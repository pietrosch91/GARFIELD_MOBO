

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cn+MKgScMmuOXqDja4nBGV7WBeIF/ysF292lfgaKjpujK0iaFYzIB0eXWu1mkHfQiveaObVLOLk8
mrHpA4NCow==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lyXUbl1fNyCoynCsgKvsnxh4xSVW7h/6+WXSvHl9VdQRm1K5kCFQ2kx6cA9GQA5tjQws4LhzjH4C
jiN86wKYjDRH3aO0ipukeid3+Cl3Hf42WJLldVcK13r9M8WvFiA8f+TpNioyqUM09aStqFjdSjjo
csyM4N1L6gYZVbIwZOI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ocYp5Q+x2567q86I1MGJbRTpHjo6XgxppbNT9mGuUHy62i1N8b9FapDfB/As1HxRsllExonP6L4i
nOrPFX5dqrfhgwJzsoiJa+kQoi2nYY4KOnCB/Pv3Scs3TRpf2vM9w+ucmXI+o3jD4h7K+rgsIuZr
FCyudD/onJvsmis4CLUUX001F3EFidOEU1Q030HzWCJJNPr3CSJCNNoHPiRhh83y8YSpsqXjqNTb
qItJOecjL9k1mrcywbi+GE7p8H60wh9osKYdQVQMrETxJObRc2pckA7TWFtDMJerirE3KnEZvIsf
rkobt3565did5AenTYngu53T6wdatItFn3vIuA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vOCsY/SF8gPSqD/ldVKm/v7jmfpM33R1VJXD0UiCtFFOs1P7Tf2U4nhuNP3HANg0qD2YjaGQ6myv
dlR6lzeuHoYmZN/DUwZJGSaiuM1h6qmcn8qFSCISMqaoZHDjixJ9JrSXtSwMaPXqwy3RINyRZxZZ
n+tFIFvhOGXInTnHa+V/8xfZhzHNthwln8CBoCm3vnx5oPwRDkJfP3YwEDF4x4X447JPTEXORFnC
I+t/Qm3ldihxuP2e3EP3csValIaPqAY2BoE1dXhtaXAVGywLawKNeUCq9IIPVqj+KxyFneku6GTO
rnMbpLS30BN7Hk0gd76CeIpd158Kv0d8sEsmpA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dhHD5W3lGGtC4CZjL3T8nBhCONi7O+vACUFgJCKoGDg4NGC33+yxWhu78fODvPCS2DpLrPJfk3bA
djnpMpnwkBjzsk3CeFcPREHpRWWK8maEH4z7l4cbfw7kGO1b7+ekrWpBI7kV7eYckr9C0k8Ompl7
lKzWRDsnDke7Jkm2xJPdMkOOACVdIUAXKGvSGFbWAwk5E8Rp1UFWwqjmBhVrZ9mRxRT8Yg3dtQPF
q0TNwwUnijSFIcDGKDKuZ7CNTFcQuy/Tc8KslLW8lYYLxncygRHOjdaP0ohBUBQua3Io4qpRdfaV
InvJO9Dh+lNQuqdcaJvi0JXgF5GixjCSKmKlqA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pz0913pmzb82uZOhWjEa23X64ev5vHsic1WjUUDytBBbAx/E1XSrB4wbUFgywP/okDl6EBGDGRvX
hoS0WBJe40mrnz7XPUgtp2OmS/NgcqGE7AhEty25v+Jxpgtk9CS4If7npTe95nuyFzYHVToQP4KB
6/HKuWIfxwjB8zuKPC4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I2mjOeLUUoNbFKbqo1sWmTLCRf6eOvt7iqKURENUw3Qh1TB1B+bnN/F2rG994bfIQZsB5fvWkgKN
FG6KCYNjKLRpH6Z5OVJR6fOANjgDmnm49QXLpsNS4efTdEf+OXCcVzbqTKCiqtvuRScAI/nsT87x
y3rpJipze8j6Nlb8T4cSSjZaNmboEH9yPf7AxUPuY/HaH+yXbGP7PNWIOYU9iBJ+xgANh+c8Rbay
KHHeEYhxcnp20ptitbVw1sh77xQpfQIoY0Bv7zFymqzyeXKX7gS+ski/Y7A9b9aGTleTt87NJDz4
ncJx8n/LI8MaThS/7y2WYyDJ5UJrv2MXzJNvJw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
D5YF7uOsXaXOZh6ypU/bp724Cm6InGp3nELa/lpDIdiaHlIrrIwjN7+XpeEVQv7mb1d/zdRZtcfu
XPcJI4IwUnsGG4O5XNXEhgWToL0TJMw4F0a1cygxW5l66WSYuWhLbUCiySPczMA1w8V9330feBFb
bF3VKgK2g2kSdcgEfezhOq5z/lblGYDYPMNQL7RGkw2OVLAYpDlZzq/De76CtbLevx5MYhxBfHVH
2Gq43uxlU8KXw4up2CsOoF9J21zigd0DRQRAW7LKFRwcFEr7abU7T16H0rVrl+bNCar8I+dMRsx6
kJlR+f8bMHnWnOMXRRED61f6JCUJzGCT5ht5qzgD/uJaeWe2uuoSyWg+/0vJu77q5fHPp4YS2Cgg
taM94DkaNxzU4uBK3MnV4rOFsSQ1DVKF1z2zone8MvKeO6FbjNlwxbsGrJWVbCRDkNjWLBOAzUOq
t/5GiovHimmSZBMnFjSLGZTHubAbafwdvEcWtIr2VVUCGPFgYb7amvQ6yXIOYb0mnd05ntNZsyg8
n4WtOjwygOnwWnSyjZyd0MV7pHktU04tQW5CrMnnaRy1xIecL0L9YrZ0H7Qk7rlTWiYeJUu9hlH7
hxhVMeXlcvErNNLDQyHZpr97uh52sl0gV6dg83CuaHV4WptNziQ0dq06mAwtU6aVRgJ0LcHIbLbY
t59hPMKMGaY95RYtAaEh5jCZvUwwuKggEVLO5dTypxZoj0tL2gCSwWkpRz28+KYNaYhDmD1ye8LH
IKrPUY2D7/1c1usgVgRRamJ0qJPFL3q5/5eOJJDi65vBr5UJ2lyAEeVOjsdf8AvfUumsflRKcD/N
+YTTF+2MALBClh2EOWWxBasZK6YzpsAXXAuDaf7N8TCoW3wcQwq0D9oh+4RCEMlLJXeJxzHywjyb
z3d9fNNsPJ/hY0LkMhoxL0P9ut8hRETBhX0bE3vYI9rHHlNxTM1w/gFoivFrWaKa8LbvjYRKKzFU
H40UnHJTDln6pT7kZ9GcnadGdl/CWmDlixggCYaOUA1U7cfE86f7PXnLUvW3n4YBU19hkpt3h7bi
0AdWqGKqigGOGFLC/rFjnYJ5KzNItvTbueUX5xzTl99EQ128wqatGPD3JLpOoywaZUqcIzN+Aype
yrB+/fkZ5qgLxUmbtrCmjeD5hXaUwb4Bx+emyFa/eYtgC7P3k0h2JTgYtkjiZ4AKBIWc4qRLKNx1
H0b+ETMgXcZ6z2HvJ3cRdd+NIhUT6oUa9zN71NPyW0RF4kxMVbNJNKaOmP6g6mzOgsDA8WQPehEJ
Xyt9uMwlAdmm4y34cF0EtQc/tGqL+ntApG5qZgi0s8/l4RQuawsycV3q4LWHoGDXD/mOsxUKOV8A
oGEwmX/Ryvd8+lNEo5oKPpTVODgmEYsk++txTlrC24aMFi3Z/7zz2c/Djq9A6MgLMylPBhefSajl
3IIR8ehM5OypeW/jybTDhy4yNifj2ZMMbgbSWFLH98fk/Vok3PwwVgv9eygyHdfGOgBII6EC1NKk
NNreuuHTxqEQH79UzQRh7cLTPb68hphC/+i71/pvo/qAk7kqova3uGXpxO1G6RFRrZ922AzdVn+h
n0BDKVMggqgQwkI4aub/Sk30rlfSo70ac/MeX2xM4SShKdxDWn9UmlRp9qa+qV/kLxRRKjmSGKEX
9jRSxN0bxzqyvIfFzhw3c3MmfO3AqJgtz2fQGHcPryRkH6/hreUzsBoh3kQ5QQE8c6EQNrVnL5BN
XOG1Vjxzss8X2S1pNjdNkMd4Pf9kZpLdXyL7csBKkqW6XbJFaODlIxDgMuLq3mbH/bmUfNaClrOl
mfCj/yOCxnsx6dUUeW1rBq7WtSHnCGrwimFcHKzX2guIlWcsG0StC2pUQIdaLnWER/EiJyS32xzh
yGDHhp8uXHckGZ7Cs+2KaeiM97q0KbnUKsFSgSsKvAte+i7R/LCdNthoEG/kkGuHOKPbFZcJiDKE
HbdrYXRP2UuVLgIr5OLBnCEZWRFqh6azIo8S8J4ACOQ1VECcKyyBcFP9nsJP21lMJ7UBCuhUd7r1
0/qvycQ91X3XAZXVYRvwGx/NG+PY0dtvYXpndWBX15jwjvAnC/RbwpfEFt9ypQqW4LaPUAvYde/X
NeJY2RBCqgMPQb2eXoz/RgLAAx4VKC59MScQ7wz3ThR6idGQBhP7YUwFpVc1iGIjoVQfkBi7LPt2
WdbURj69XiAkicX3ow2NOAAshqxZmm1YqMY+Ex9uqZe4JrgHZc0Ro14722I21P8jtqfHAd4uvLcT
J1AgPPBcQRgT4K9pMDeo7JZ7M79ygo3ETeRvu6HprzzDPoVnwR6ACbpAoNIZWgYitXPmTffDK359
svwhCV3vncZrVxD98ZjxyuiiCqDfHebfKWJs5vWvPXgg8Fhyp2QOBr/Cxmru5AZuI5I1efXntMtX
lOYtAwqSBt9LoePVfZrKpMzHQBCwHGKOnEplH76XaTmMUBF/Io0B2pMMZgwPQ/rKaMOtZo6NZvXM
ZHg8Ki5no5OrDvVYbWMkZu3fy9Wn+F9tU+WdrjRPN2HO6O0hY7hZxyGTyumLjVHfVQK54XAbJWzj
a5QQDvaJnVpDnH42ewPfUlCDN0Aq1kYrPGzoW2swIzgB5JlAYO+dAlyFQB3RzamIFXEkl9y3Jlw3
fPgykZizokDkE5pJ3m2M/Z7KGuqriP9aI4a4Y7z1VisjIGtf5Q8IoBZ6IGP7cAtkDX7j36MT0+rE
yUxoVEuekSyl1lsj/Ha+MFrRqCTJlyWOyMs1LrrPJR4CLBen1d5Ol3ELQtBVH0XiP4NbFVZTT1H8
CV6tIrL00Lkiff6cmZsplzE7yx8TxUdW/XaMkJBg4tLHv6HWctAnhuGfBWDMnIG/k+YeXHwZ9pNy
YzSTqiTchmzNiRzaEsBvqlK+DIqs0wGMYpriqYY9VwH5JglGTQyfCL/Pk2VTcZKm4XvVkypeqnuE
jGZ7tavP1kozhjH7YlbPYTEunGRoqEOnnebinH2Ct1RwS6y37mKck3R0GSNWVsuTosiVvNW9peau
CfiElLIuFPUbQRm/s5vvtMb3wiLc+yYkRvapWk0T8X1sZ71oMk+kJj6xLb+ZjJz69kHDJey+AiSJ
tDDMeCSrsUZRHOeDiKfRHZZi1DmrS2da8iOOQ3XwONjfmzGomZFgPa6MFd4B/5iEvz/ahl0rquDX
fO+DxkuwoSiX+WGRKyTxaZ3Adl2bfIrjmj7EWLsM2etEVhwfFswmUa1VVnWc02woJxxvaen5OBlp
HwQ927t47gA9PsZF2nc0copgtqYOt94PFdiQgabnwbRTS29jGcOuhpXVgOOgRHumaCYDehuzMEh4
QJPo+UBzb3azdJmjzMncU1hnkjKv4Hd6FF0yPoXh5OtftwlUpTxhQsW2grbQYxGAaKK5JvQBrNCw
BN4fON/XQJhTZNYXpIt8ljBOxoZvogmxYsDE61vtj3YNKhmwePqKdDdCT8jfqXWf8iz5dZdM84Hh
liPO0tQ0dmNoz68eX9NQX7MyXT78XB8kwQ8Vq26MJOE82GQ97XTIyS6GRPT/CaGOENRASFQF8riB
f8eDRjHGsGo4UHB1Ge92AzbJyNNCGAvNB2MZfX90COjuTkR5Lofd+TQBOD0AqrrZpABNj16WaF1b
+NpZctEr1he95U6HiB/gVWwe6VPE61048IFD58IUco28Oe/TWUjiBUi+gcZyi8jlscZp8msY/fPk
yLMZCibpsUg3YCppyincLUHPVYsYOHKTBaNwTUen0YRl+4tKDlGu723sOi0QVuohwvV64mj3Sb0d
6NyUGTNFtYqaVZpQQUN1VLpJ0WZG6TgEtx/HqsPdpMuBdfy3Yob30dd8EVBQxm9P0jISDUZvGbvo
ghXjpqcig5EDmMTnnPLAKWNoG0ncZF51t4JKmq0boSWx1sgDIXxkZHyThezbueE7KVUMfe/qRsXy
G3McOK93nIYA3BQzgJCKXXb5BBkkW0W9wFz2tbdB1V4RadEXQ4Orm+L6ZcvhMk3RBQ8VQfbl85rA
mJyXutJ/dqS2lM353bLLB7qb1BRu4oOmPPVopzShishKAP754RjEYoBHpvSIx8rZTI0VABFHpoB2
MNxS9PY6JcUQrhzf+AJiulKHt1D3DGr3uxBM/5xwZFYobBThCnam8LfQfvYF23lhP+mTUApbBFMr
wURlZuWG9eHBf+R3cciMkZWbyKC3igQpUgr13n01u9ABaL0U6GAeVWja3OAwMfmZk3jGzlXLPg3K
R4jAgUa/ykdHBGPjV1csfr2DxlsDmJ5tVk5XL98XzRSQBNjMSmt0W+6rmZOYpxwGAxKXcjY4tIQb
Ixj4yoPgn1qB54/0t8ZcCwVOxN3dMs9Ym1SpN1+T/Doy6bMVRmIagJma+SvLjoGxtlbq0cfw7eBy
S6hc7c0/wCdzMrjYvPAKwg2PeNJO++NoHvnLlLP9nOcHSphFOjeTAKXfRNolq78f7PK5twXpUemQ
+sHbAAYV1UES18vUKnCkmol1cjTqs8Awn6T8Gj5Z/ftcpRIS6dr6WFcUEAGsZhVEDuTLEVhHIEMO
CXZRDNNtXCPWRhs9D3TuiMHdvYk6CD4FeAth9IDixvJBgM80PrnzPyaFDmXk4DrXIhqTZnSdIIXp
tKq8/3njBCCtDs+Gdxc85yG63TGK0VejA5EaRAWXw7yxRWdgC1E80VCt3sujj+0IQ0mHuY3lSQ+L
PvoiLy5/Cs+xRB/9AcgF7Fkf3cXRxnw6bBWSOt4BsoU5zVAebEmY8hfQ6SxqSWrDZa3xDDdW7r91
P6alQR6szaE03iJY43l0W62hrRtnntpc46S/ZdKQxrUyiJAoTyAUENiPsEGn30NEXjLuqnTlaeB0
TnwDaDJIWZ38oYwAGDvvaGNC5lEtBKGtoVk7cOx/6I+UstmVF1Gljd+EX0IvqfQTrdwgEIuSKI9f
rfziBQDVCS2eBxIldkoBuJs++cbquMgLTPsw4wITjETRNLuEf/DLF/6enIvRxW1LEcAWooSyXoU5
PPqecMIvpgOIJ36fVHp725a3Ufz4i8mUWjooqyJ7Yu/RlzMEeFklCcW4mHnljo1jNTuEUbSgfBm9
LzJEiVp0fy0Q/K5jqc9DfeHXpq+CVLf2vb5QNK9hccU0i6vI67h0SOZAiycsagN+aUGTfG04Wt+c
A1s5Ul7BpXouzS0uSkP8x+4bIagU+8Sx5drazwJUM5V6C/5PdwRfGNb2S2/B88W66NkHyFd+6n6P
CO0SfWGmM9VfO1U2Go/PDBzYFmaUm+K3fGzREjk9CKo5s3FHIvXFz5FMZmFW14skI/xkWRvyXdZ2
vR7+rICsoIcAEsB6Lk/itZKQeCDRcDYU8n3ozbykWWsXZkRrjbQf9tiBedy11Al+jC8QgycLkoLS
kjVkhABO8BwBFvhJTWBgOV91IChvrh/zc9zS7S20yfwNx55rzWgNROehishXFeBKm32jxHV8+fOK
RXeEDS/1mo6agzvTiNOfNXfceR84dZKPZMnH2mcRn7LEjuR6AIv9NGPug7mP16FfAopH5bEhxWWn
jJwozdKLN6YwEoWYbsVDXMC8/ezoqjjHiDUAWU0PDU/gy4alkd8ausmsqmGAGQXyAwlX0G7NZ6lT
qAMPHlFCUGeVlh5k9N6l6tw2aVODeoYf65PLkj3okEuXHs4U5xOK/1ShhSjPZ418vgtVdO85ORqu
QKZWk7wjhVIwS7Eo2FutGkuizT5TXNMLscNVDRME6W8iS5b6wwTtHcCVCkV83NEU4/Oq6vsPLFaR
wRoqAyF4TCzGNwX2ZWuGnRxdnCgcNo9M40GiGBrjLMTELIpng2XOYgjLVzjhiLuRs1CC1UosPpNN
xSxc6iXc5Lrplu0EER9P0FXCYER/fvGZ3lGTnNSEnBe/mytkUk6XSsO3f12qgy77Dp3W+Wja2PAl
kKsotAN6qcPr6POW1GviuEFXYEKC3mUHJ/5RJ5/vKhu7FYWT1nXVEAjx+qr0EKmEf0JkVDELAzjj
rfmptY8llR6W+ecSCMEpa3ViWAB/72n8kUzwMOWOQ+lHyRqxJF0F9IGe1GMfXG6TTIOvWGgm8jFq
sT/zdtPlktZstnMhUxLbMMUY4BnMhQudiFFs8fDIB7lJ8dccDwMTt/OmSDOba6FeAWkCEFEKvxjJ
whRKn+BUMiW1C52ZEldsIwAY0DJRi85Z3PN2Zv1e/+WxKnI+xTSnv2zy/o4Hqo2F9nZM7GexcT9i
VMTz3a3sN3+GYKIWSuvrNTv4hrbSfzJijlMLyx5QfOzPzLXaNqv38n1+A3k/Yz4LM1ippEDZCBJP
am+yQSdjuCBt4m+KjNiVv+lJj/Deb0bCZr4k6A2sG97C+iP40oAQHF53B9XQqY2TihJgUpH5cN9+
u84qGA2HQsBwy/A28BCrccc9RKJZpWt+AWC1Dyg7KRnyVAb21Ki3vsQ9invmvNiQRNR7S2Z/DkNk
sqtT60w8t47LehaLZEp4rcocz2lTlWGoFQ0MLllsS6jScGfCBq1xhGkFqlRwZtKz1cN4lo1q4mBp
m/oKTD+BLhoo6mZS1pnH7ktOr7OgUb704PSMpYe3t9Ur2pAiNJBrB6AscgEgQaZu8wwC6xjtshkP
PRCFpR19oP7T55hO6G01UlCJAOGCjofCYPuODvpb/EycTTj1CFTDOdTK8M7zK9FOHECgxBkd+2IG
fc8+RgN+E69i86WDJ8tvkrR7pDyaGPKlKWABKerXRLWxz0Xfk7Y3YE+QpvqOMN+t6NQbwxkqJUTo
NDIdRce/aFn9D+SQDQirCGh/9QmbG9CRTreDhGZ+yVfgdYR3ReT0wfF3cc4rqXkYQeFDNaFk3spj
woDkD+4Q7ljIVxS1rDQeCMsCrfVHtH0NKRvFDNZDKb226b8sypGUF/Ht3uceppDbu/QMfP4krspC
dl3iEdTjIOVOJVxlpuPefyvKuaCZsOkGzi4a3lA3xKr8RlyF/X03ouHEGsWrsmE3QrGYT2QB7p4S
0ejOvC5mFNEWh1dwPwv6qGtbNMVNz/0RStoQ8tqzPMy8/QJ+o/FIyK+mfmDFTpByWKq5lDP3jy1g
V/XrI9NtK2wyLtIneF+Kz013s8hT/DBOzO7PNQSnzIXhi4z2KkYbLBFXMsrFdS3ZFb485JCQCuxX
9ewng9GQXY4X4X1l/8gA+q7ggiVc9Wxo86vz3R82WWsdFR/cih3+SHBVH1hc1CpSX1u1RRSaCZw5
4YZ8WPVNsvZJztfnwiWi+fyqL4JXf1uy+ELEjcHZOzcgMSDzJH5wKxebPJG4rd0wiAyjLR1rxRX8
UN9u9JB6i504BLPpSbfXxvYxlSGwvuKl13lXTgXSt+e+9XUtnhHrDHkwAx6OJh3X4D0oS9f334e9
gsGGY5pNkYNbf+J+UXdc3GH8oEgxnwhqUW6rQ4oPquinCc8thtcaDXyLDNBr6X2qVuflP1AagOXm
zgxNEhHKTJTDHOQ1gSBT+YAbNJwfnVz8Yk0COD0mJCkPY+1Mc2Jo3z0HTYK3wAiZ51AK7ClYuY5F
Xr61BpbOI2YGuoxYJs4mGjiT7z7jtEgsz5vy/aKX8myrjNDtuB7Hmi7r9uwNAC13W/GxmjIr1Tgp
iBhrwTWyhIFvKbWVsH8/waSJ7eEhpB8hVvvTqbOo9vnW1XckEw7AfOMoHvZHjGFCBC7uGEL1GzAN
BXJiINKLYKXvUa8ABi/eqZSppJlpgXtMLoM3TiAUkNzAYiwwM0Ho4o/3Y5XxlXIIxo00/q6xNxM0
JN/Xyj3t65bY1KcfeGvwhgIi7CyR7ENQu3uFLglfGCxsTdmtHsPdW4Owyw5cDN5qZBopyMu++1f2
M/fSzYUuiZWcNeWkhNxj0lFQGz4/wrUZPlc2+ZvM4mKp8xLYJVb+3KHe08JFggr005/2BUCRfYej
dFOjmx4WLS1wDBG8ktNzRREDSuoDq8dS9Q2SyVn5Spn6Vj7L9WxeqT3Fz0A5uyfa07Ufc6SnI1NT
U870YnaGFHSt44lMKOJ04nDNCoGyJBWI3C5gEOh8rgh1/iMUJsDjU+4YldZGaUblRcQNGIJXwOBg
X9FL752ic3yRHo2S4joSoL3Ybp8Rx9LQfbIO8Rf69kjs3YoOlu8k/qFDQosnzqvcHq+u7gm6PDDd
6ilfThsghP7KGxDcCPRf7aMhaM7KynqXfLs1p1wHm4rzvKMDdmBo1tg/QhC1+lwTI7s5WkQ0/nal
P46Jkofo2L8BC6cujA379LN4iw6kksVpMsFhj0S8Fdth040Kr++t4Uj3+c3W7cw62FyAS16dXHRI
B5tx+MPD6JQMFDPJ8OUPbIYVz36fC53QY6w4YQQ3i78OumkqLOvpGBP6NbKBGoH+FInsHk2SYNxG
O42ZdCQp+OpmTMQIyykuj4+gL4cRQb4BDJvoQYtQmtNy7iP2cEGpYqlll7FZSmeZOZA3jt8K1sDD
6+STMqsMKoVodC/bv2nUGNzsyGWrKckIaYzJdrKv0Q/+peqUHSX0SKHQ3iHFBvXyw3mTySPtcdKx
5MnyMmeuCqrpzcRPbPlEGnJo17Dg1q+vO9l4XvgmL17pjoyE7MSlCer9lJIjt0G2QKKm4UPRwd0v
0WM0ZAhHdjDEtW+TwlJr4gXUqFeh0kSLdp6DvpgMUhMrD5B89UupntL5BSwPJvJLWc1wqS+v3BBo
H4N07OfsfLSeird1ogLn6md3A7jZCeeg+AMbVQGbNGTmc+7rti5NJZP7Me9MJA0+JCoSLUxKDW7o
bpZvVuul56LiQDa/JToetVREDiJms/KtA8SONt5zMq6raC/s1hLQ2nfwJLGfBNJ6gMlArap/BiK9
wOBRAWQBLHLl6CA0LCG6c8iSHn0HSguF1gH9ZwSAgR4ET1gMUpniy9m2Kh+A7NKpJsQT6QOl08vP
XOJooqJ2b+i+Uw0q4Xajvk5K4OObJjQBA6rrRv64UdDcdFCfYx/n1yiaa8H3ni1VVfiOXk39YPqE
UQUxdRUvWQCx9sHCCfgdiaYKckbHik59vrvPnjKBOgdISMujZM9ijyOXWq4ApRkphOMMusXWoMh5
782qYYxufna8L94n84SUdhUGQsMwrZlWL8mMc6zH9dWYmVFcDLinO23/c2ubitlp97s11PvJu1V6
BkchW7qNkHOopmLf4eORObRNIwsZpI/qPnuzQcaPf0gQOD9su/2F8ZW9Z5t7+xXS56wHg6W/cgUP
TnhiN7FJnQhDcAdzY6tgAvMeQvwut6Zm+2ID09eXusVgJuzsZ4o/s3GnzDC/fJf262rDKoDmg1NJ
XzZq70qYX+/R3+rS5gbVRh4hctm+5IqBcx5NgJPJdVkpwoSEbf7fBPA7fOeriQ8xbCslzxkjIx70
0errFssLnyCZdrhDXPqdjF2FOst5RauyiHsPneUO8OUJRzlVUuONro2XZPs4qafqhrymEpK46/39
1KofoYjDXR0ZTUat/S1SKJlsDmHePO3FAj1QFqdmwNx0w4QWXWYAT2mCgYHqZLD6COqlFY3VEsEC
+B2rv2Rft/kb7mQWeTFXohFmm7cG8Wa4i+itVj2aprtTpzOPet86NYXtVbup4CJJ6CI2YZl07ADE
bl2DlQ7ZrAD2XiNjZj18okdmbTWu92rG7YMWDS7eKz7+9LlOVjxxbG8vgWaBhneob+4k+gJ8+c5j
QIdyf5BoUApPT2KbFj/bU4oAYYJiB+k8GSTdVQKb9VY2UOSvDsZz6mytZM1ziD/K9tn2ddD8kNmW
lj3afxD7hj21Jm5F+K7wjQjwXI1onssec0NY1FLVGJrXSnhjDK184Q3LjG3I6R3KuPEj5zwNRARc
DffdxptU6F/LYqt3SLzjYl3+zoh6/H0tIS5X+00ovieXBvhJe9UmxIMYqEZn3cYuQh/S6vZJJOsr
r6MCRCVlJ8Hm1xG9yKMJ4x1PpTH2cZreAI/W+MOwW8VM2DjwEbq/yQAosuzohHx3gD96kpycUR7c
mvH+iVI/7tRyM05cyW9viIZl7Y7ffyH8AyuMHmrM61st26+z2gzQg8c9d0y7EJlTjz5tvLgeTTcI
hyp6AVwpe+ecO3hiXhC/XSuikEbkV/PUqug+qxQhuU2ivMZ+V2Lu6rtaoczmDPKI5m8i6rdp9UdL
GIDh3xrUzc+rRiDn8aDcNLq2X9YBf1BKb2IwIUWEeUWeHcaiyCc5jqYfShzWoe+mwocO4eE2onDd
k8q+mayV0ZE7hX/zeDy0z3Pc7NNzzPWN826ojABeI2hMjy0S1AusVdoxkhqGD45bjmPBhdzf8ghr
DRvc1az1ZlRApiBm29THeDpubGZ+nem0VGQA/gC1v6VxFZDw/ZiajM5IcOMjhqfbFDGJsscWHnJ2
89KempRUHarj/r2em+kzTiTQjO91QyxTeaPeJWnXL+8o7w8s8YQ5NV86FxCq2sWrrKSF1kUzB1YA
PVKEe4okNdYk+Om5NuEJqynltNWviQdaTSczHtbiIvGqnVwypFta1x0PVgWFOwil0pgBr4lDSVZJ
ofeRQfJJCbosY3sN6kiBo22RO7bFTlPMAnu8eMJXCInsIuQuBTXEuvyBah0oeBG5tVYuqt3JS52w
WzZp8Pg4bzmsNY4E+wyjxIJlOT8LckhEUszer4dx+nWicZmbsLmoNFB+boK0/+m5Rt55FiV8VTzE
YlRNlbbu4RltDPnWan5ZULaqfnHi/l9Iuh+BLN9WwxTJGl7+j7T1uHAgTnU6YlRMbJptd0Gd6Xrz
eybqXPZhuAik/pSnHt9OYh6w0SN0fh1h2yD1tGEwWq/2HLh29e/scLMa8o6KkLGLg4/7S2siy4hj
HRYto3dGO9DRGc9KwPnE1AyegAmrrYUe1sSWGIlT3b/n/1G1TSUkR6caDBsR43cE2I+rr0bK/sHB
+Kkc5DbjO9SgT9muTVNt1Jxhj7snFmNeIY/IzXwlPZAN/9txNoj21WcYryMeC/dhSKXV+Ylq3oax
JBoA7UMx3XaVFb6Z1UJwN1OJdYqi9+Yzx7qzECJRLj+Tuq1Y1eo/YMRtZ0kelKd8hyXBsRqfJG/n
Bm15caQRgt4bWjM572ETuAgoxzX2piIFU4nB/lM2X+zEMTDdgDkM7rlIBOeJPIUp68FT5HIpx7Xh
RMdcrl2ri9XhcDGLaZr1Efnz00Jv2OD5QZeXCv4RSL+jL+ANDywGqy4jNL4ZC2O9I7WLJPMOAwmF
afGhSZdDGXK77nfbnMYMdLtKeemqYAP9zZXGzalbu/ClxFgAoRxhEp9I1ERl85jL4qkoK214VJqC
sq70jXn8ahv47XshobcPfqNO6/lxYrTZNPmi0kV79FIcXqdCwojdaqkGtHQtHJYkpR3O5slQgRvf
00qYtD/Q11Ea02RLC7M85kuKK3SW9Khp0s8enGGFMAF+Kl4H0cRGIfbTHmBCFjf/17sAVSc1FQWF
bL4LQxx2H/+PBpuEVKydEm3J756gVRbXidggRHQRFII6pJ0ouTDbpdRChl15nc8b9tw3ZQa5PWBc
K+R2MqJbYqxwDVljWs+OGdeblNg7cGga5F7xJbULZ6P4NoLKrCiCa5flRHP6u4uM9wuCUVdNHgpp
VsqpLW0EuPGkXVOC3WYQudhfbhhHyyJ3b5vue34/GK1wZs8+la/4iWTpVTVZPjaQhhNcmv//XETm
nFLoBxCqQU+Cu6T+DcB72QmJddJk3oA0JNoIMy85kVLjydBwCmy9D/HeQJ7604MdJd7s6iWHZPnK
CNFD48APGYr8DT37wkz19PCrCgVtzITv5C1o5/bw8xe2MN48SJAlG30sKBoEa9LgW4wKedcTZ2n/
3c/FA2QTNw1bUoG2JGh3K5tELjuH8mANlw7gyDK1avM2Ld7B9Io7cZM0QV4+IIAvB7EK8h98jiys
w42JqV2S2bM8pS7CGuV+fuu+nBtG9A4c8BBBYKnHjcbMxIjvTMM7/x5+eVPLhIcNJ0WaSNtTgfa4
FmGIpZbO6rP02Yrwxh+BpWAQgk+G8+7rKI6wpDwuamxyoHfu8Tyvgh/x2yzi5sxiJUsRzIH4NaM8
+mQJkpxmpjhBNTqhZFRYBLzzWmc3PrE6o2sHhpaug3h3GoRjHVRxDYUhnbmvKjVEbUGy2Yad2MWx
Mr8FzKPfR9aHVkfMtoHFf/8G9jOtpcmilYzeNlqLXeKqQbNtuOzqIamQmEAAG8Np8503AmKUcQnL
u9obRgA8awd9bbutCJSgjrDqrRDtJYoFPPrtFxtBjU5sS+ATkqUfkGnMNNZwVixbGlaIEXFUEGMR
u5aXAwejd4nOeYK2v7JXewy665lkrHDWIEMnaTgyhlsv4DQPg1Gc/mHwDajyG1ToY7qS1eeuFpCJ
13vEJcY7fy974hukbiUin50ZcgNQ4mZwQKE9DnoZMxwZBr2cmlKHeVjgpR9o/PVc/oarE3p08MEw
qIHeOkvh1tnQ4IGdOEbRKgpM3uhfguXtVsUUmwGcaAQlw29Z6oxPR0DqMixcMaWSn8TFK4iSfKBk
18ubXHv7Ue1ZuwSAaHg1pKzfQEtsE+5HvlO0NdutHzWEsuCdn/9h3QeXxHDRs/3Yke1M++Lbkffc
R4lwBuMp4afPqBsqRHurl8JR62rptsXbmLCrMNHwseiOLoHNrTDPLJPPAxd9JQmy8vWJwEJ0dwul
sh3nMDRVHIgQKRj7x5QcQIqvZND5GHYLxvXNGYjNfDoF8CPadW+FVgw3654mBUaV1YTFsFMDOZmm
M8ywKjfWKot+bUIwTuxFMYYA3oW6nN43IVO3lW7TeydugpyHzCqHiVwg/UOLEKDTFbrYDpz/OJlq
Mw89scMb7+NgPLpyMwtFHwwk4nw5sd8Ti5ej0sp1BJ88RekNJfLNBPXAyDYMQNzU+LB5A7ke2xUu
6+poRgFW8LfWS1JIikrfpieDEQFxInSeMs6oOkx0Nj277I1hsCChL069nG8izIQCgRzc+t1i1Fjo
qwOjYbySz71YhffsE1xUgatIi47ihjgbATgrCQTF1zBBpqGL/N3G4GgYqAjG9YF9MATSm25A2nqk
m1oX0suzqFQ/d27pbD0O4ssOMOtsrkEMHUvqWDD+E+MYs5jyESlp4HBGDCMLXZbV85A9AVMjDtNb
0YCRcMiQjDMVIgmoCHMRHJhvE4CYxu1G23NsNBT339IGhOKwlhhHKP6U9XwHO/Rcoi76n+s9ydSg
f/lFnYIvtDAlNynsUrOp9RaENGKRTX647rLQUmZgcwLxG6QEE3wNZKk99nu4XCVOzbkrVV58Fqw2
/G92rb2wwXcexAaaANdS5XSky7thOQWvCXVTtlIRdpe6sbSrIIitRHugaR88mNlnjovAKOQe3dhG
Lfid5JN52mHTecR79KZV6uzJe53dQ49HjiZJ/gImlC5LrWD9LSSmLgmTtemVBmCqLNxsH6kBsovr
IdANMkps+39DXdu8Y4Bdx7QHO3AL04P0XgHOsEc42U4kLaeJFUsbYLNqmWqejeVR/XT1HzBWqVxK
3Zaeq9mUCqWlcIz1M0fz1h4Thra1fVFBrhkggpvKTfGDWKGO6gwAa290XsdvyfVQQQE2ZJbD6BHz
IDmd/FHqcEtx9EHjdlqnIMJYZV+wyB4VxgaPvX/m9ek9y2T72IKlN98xA/HvXldKxQMQtiFvfVAV
480ACtloORYb7Ykznl0T3p7FDm+XejMC3YIsE4XreaDVjOjunlpAyGQoenX9z0V1ds7QeIGavB85
RdO19XLRKWnUwNeJ1wQAgA6SbfbhW9DcnykwbEV2+S3GsXNjV80fP/5VPLKDorl//yXhR+Pws4J0
4KuTeHut/wmd2uy49yjdJqyrgDGUqDJvKewQYzaPM6CmcZCRu46Uesc4oCyqPT2J2/eCJm37ivdD
GeeGnHWd1goALx9/tx4yyBI+EwDqchh1rIqrWXeLDKdY7Pru3IZV4yiUomI5pIod05DnLD13AwJ9
Wia4LcBymV45lpKJkMOAP5C2Z6GfcFn3+8evvFKpg9epCPJ6xLnFqYmdhCa6TZ51IrFfkubT8s/b
ln+V+I1BJ8L8/Hx5/YHDfv4JNKKUnRjLSgoYrkWBeg9ZvFO8Id1eCr7Q65N04jQv+2AZMstPb6WU
sybIkYcdqckQ7UKIIPDikCVLgqSmcDwipFn2qwmldbOg7J8+1B2Umb6mUNR+uJJcwKp97cq6cr50
ldo0pdovFVBrp9cHxRe8B62VhTbSPOmBgYkyYrhq3nAYx9/XPKo/qp4RyDJ/Jma21alzZ5mG9Tb1
4C/8O/27d2dVr4nJAKnvoFNuzeDfmrHN4XqH+IaiY+m7/9qgr5/zIzydxuJ30/zRM35xtbl21q36
RL8KD2nq7YJ6jGZ537Fs7EPn37uhr6kJPX8Z58DkUuFVl0jPkzt8F/Fvul1ab+Us+upj5Slv/3PZ
depTuEXVgCcqCOtg7WKHcjuZvE8K1lBFgzYY1tGuQsaIeu7vpaYdn/seRt7iMloh35xx82XfcVhZ
3i6Ws2XHJCV4nqpS/AfasXBeB5pgkV7nB7RnV+huhhnJYpZ1jA05NVWr0SjqklQm5XZ4td89xXwu
6vuRyEkUVWww6CWEORPj6zpjIVRjVC8eYVNbmvJvrRAzWZfBQdd+Mry7DexrhSoeagqgUsD1ufEB
/2CZ9j5FK9EUmEnXkfxi75th6YQkVi3RYrjbJNtmTHEueqgH7sMWuupbTvOmyfDAdhG8CupHuGwI
sW9v5BZ1kvGAs6rmqPYKol3EXqilGG3dO7Pgikj99g1b6vWgbNofqGBdeJzAEmH1H1+J7LgyNig0
eF7fBfILSXYhQADwStqIOcdswgjp6OF7XyxmROapA05676APwR0EmlrWWOCe2k2M9H21sIwl3jUx
DgXzglT/rWsfNO462vdId0I+7hgkDonEhPKF9ITtCm5kKj1qkw0SFieERS7WPaQ7T+Mj7C04DGv6
eJczwiHwVB5bu3ZFL0Id4A49uu4/cwz1r77/RdpqLlM0p+bcROShbhNrUzJCSPUkyBAwce4jPf8l
M+aEOkNU6kyIQdk9Yl/S6cOWoaa2C21LYMh5OqX+d3+/sHthzrf9MPxP0PPetCWmhTppu7qBYg9b
k63iJuY1/h58oFxADz0hVGejIW5njWyw83dWJMMAd1xkenjq9a4tCd6aFSQtCLVWaMF4bFGGzH/Q
BYbN5zpZczBoz3h3+DnWX1nmlWBlJdiWzIZu1agNVl7CGRomH6NTQy4rVq85YCMdGsUTjLxn1tFU
j9/qt4N4SoAnzwOOD/1z0fi6Ba9ZZyok1aYJDrZOCKLeNTttQ2YQu2Yjx0eliE4yXsTCl/Z6orLf
ncdoxB2VMAbRkIKQWIlT6LjVSTY2ZKacf+IRIppji8PjL3apfMhaurqSbnNZ6gCKcd3fBn2lS5QU
YMQmnm1rKBbxPJo5oHjlwQoMLm8+Bf5ujVUv0fJEp4ok3xI5CbRYjJRbb9ORY+Pl5CwMdKVfepHF
i8S34NYN+ZVd09vK5zOz3K9FvctSY3ZfqluJD4juEKGMI6CAVg4hxPyGYOjEJCmTIsJB8f8xUjcr
l93090SyxYh7Z1BIyTUhfUcCV9ZOAYIdiRljqtRGeo30Mnb/MkIvcFvIAVH4/PO3t0fcccs42JNh
mRiP98Nxz4COGw/L/siBv3sqnJvyPT4D7MtkwaaJO/pRApnLfC4zWGXjHmVpplofcmYWBy3R/cmj
E40L4uotnSJwe51hucxtjbxCXqFv2IP2HrgwPGQmZ1uVNQOtThlAJeb7l/EJY0ahE0OlK1HP3A4T
iQUO6D4haxXHxwz4hcfspi9q2Av94pVkP7KqzxO38K+RiboSug+YbVw08J+/t72mBHk+Sx34C8Vt
6ClpB8SO7UkL3TA2WHquQcNZG0NcwjvtqOT2ka/edx72eShMsRoxxFmCPM35I0XnRjr+QVRo5nQP
f/GAfCglZ9AP5T3sikexWfabHE30LP/Hdl4wltWkAmV3AC7xnEKbyXoqjkjO97nY5l7fjlWbDQ4J
BOXvKj/sGnhGh+C1AskV7f7Jq1FgMamX8PxSKiw3jv/N8TyF9l0i26OYtyz/eTFRNTRdLXgDL2RJ
Q/aOpIuilMvQTh7eRFTswHBShO7gGaLmxuyWNNrkMNNYbfzUbQ78OQYIRV9dPiFc+aurGw0+7Id5
Fxx52nggB9Yo5ibz7kduSMJIyKzkOcpGvlkRVP7uzp4uoUhAp6Zf/LAvaFHeZgktLNSmDP/bR1hl
GDvOEGsVVb/UTu91lneUMeRgfJi8gGXJ72qclcGTua68oJlU0VULrlwT2YT+a2ijPpw0DjDliRWb
7XKeL+CnTBZVAs2kJE1VQX0ffq4yF2MnF1glShBU6hFb4GZk3dPEpeP2imLmcaABzHwi6NnWAn4w
+GDChf8xfYbyzsLZZk5LJgsMoAUW0XncwaCj6Dmct5e5okiw+2SN9MukLsdLDozpmqvdkGx7a3+D
Q0jQ6Mlc1rwen/96EoZyXmYZcrMQ1IPks53B7gXIhBXWxhKpkzbDIntDw5ye4PIBXScco81ucQT0
PuUsXNn+h6v9BJQrbhkEBshYN4RbWFoqhqqo6FbMQ9vt+IYodaVUUjiAkljQ7wlbIGl+o4FaMeow
sdbuwWcv9pZY3VOfSBUNSL46PDzahJZEzgbRe2GiYS/ROqAtEWe3W/JvUf64naZn6NWIMONXin3p
JEhM7ziUhLsTPuPdWvNmyC+ZsuDD/BNsNxZcPGpw94UM7PJOhNo0Ndb/VRNQzXojkMXjKrV531yg
3IMJdhJvh/WzsyX2nPz/h6OJ7iuetsBUMmhY+Kvl93L4qU95h4uDZnqON0leoAD9p4e3fzZ9JSLC
E20JZgIi7kdVpJGBXKv8gQhL8uXH9iII1zf/pn6OwIdDUTbAjfF9w2/TxVziW60Q5iD5fpUhyWJ9
JC5GlYtxdUoPfOkFlI1509McxZ6rNj1YAGyFmciQdpEOXSAILCEV/BNW2/EIMs1hEwmYi26NSsnX
A7n3Wmtxs28LAirSW0coij8X2VHKtQobjpID2YF60lmfIQqs502ad6uBA1AOrQARt779wzBsTfva
whunVQkF+Du9TeNSBFAXeG9+t/252fhHjGdsWdz/g36qpdK+mrXpR1xPgGQPx9Ggxvr59chPJKqC
GX0LFk3g25AEkjYWyBL92W4mfIDg9fjljIbFiDF5qI6LuuBA9mlaGv3GKHeVkgYdX3t+CwnzbP47
IOOfmJgpR5IbkDxd8IEe1tY2O9TvKYmvJL4PG+ui6j25f7oHu83PhMUWHp0/WCHWVcbL/8/k2Goa
ZXQcdpA61EZidbneisETQkHKDzyLSOPlaW810i6R5oo5smb4M86t8z8GEaTcU2jTYV4qbMnqkoj0
TyaNia3shz4M3yh7GrudoXaFurlvlnfLNOCBM3wfm5t6XU4ofnvmY0rD8Xg1kCui5uGop4FXGQiT
MLcQoAN+cXLrGOyX4x+CXXjOrHzstATcEA2Mw8RCZDXTy0XHfTK0jkxgX9gqoWVCPRtg021vlcux
Iux8PYzDqx/mTELf52VmRkNnCXGcnUJ82adFEh+7TAmmdEDCdAadaU4NK+kzhgNk9Cy4ajZitzpP
jFuh5gRPfclbToLr4jwL+ux7qni6kZRvQVELJbnmDayYqOv3DH9nhnOje+HgpHAOmOlQMQEcFr2b
rEZmZCm/gF+Yk+Hk5Arx3UjCJWNlE1g3pzj1q9TMEUgMHkGICnB9C84tt/IijzuednOoec0nIwCx
IgrGGkIiADdZWvZcd+9F9bJLgIVopZn1b/pOsrXVtrRRNY5C6cICOofDrS+ms+efN2XWm59ciycO
bEO5Y3WGxOui1G5I2OU3UDP3G4Cji5ZuFHDHmt8cdptPRns5SVVbgvZsXVIWj7hY2d7kDy89NKsb
fh7gbmcybj4ghOdj6iC9kZ07IqjBKzAwa8S39fK0J0t++Kiu5ldcktQ8fl3lDfTcqbehi7TqbUor
OyVtuFmgul3OOgFAelNilJdFp6/RV1fWW67SUtgNOz+w62S76v1ySFEHe6+6+ifnB+fVx64rAm69
Gh4w+Z9baPpY89UZSU+5tXTmDXU1FzF7YLY+sRuCfm5f7Kgt1CtXshR2Svf5LsKYJlWRu/Wp5vTS
5tPDtVnQQjnEpO8ypJ6nXMRU5hDQQPvwk6nWFkrMFMMwcLNl6IvvdPOjLKOdbq5h4MWDo0EfD1Je
VLhHW5f1xX4kt0gM0fZreqrJsDj3nKXoAq9LfIc5Mr9pQl5IiSHbRkrjCsKyRr85uzXK5oyutcPK
sZJ+fq+O6+MxkqKvVVIpB37WOk9/BVEfT7QjT55H3Qew5uuDWJUqZWneXTbhVlLsnNcwA9CxRIcT
UCHXAFqx3vzTSn2ERM/TeJKLwA0mFf9lpFqnUFnP0NzKzQebXKP0yKjwa7uo60RFTH/eDSSZNjiD
jPqIFkZ3kdynDsiVRqjp6pMrxFMeI4hWZHWdp3ZtOAarKRvMiAxrSlmrs4d1HZBQFKkcII3heVCv
Dwhgfi6TeEDhhppSm3VDEI1rSpnr+xxqhAYC4+MQoJAPG4EconoLzyE+tEBdkLQxmICMayTH9nJh
ej2zl4Kp8SiTVLR0JnanYzFXGMyWDY/IhdL1YPJoJdDQyLdAuCE4Re7oZYuBPFLR2hHgYF/Zdb+X
CN50zOIJTZkWnI0jPmnGQW/5cKLBrN2Fl1gUXE4exr/2GX04FE3oqeqbDWePRzSCm0T4BA8s1FGO
HfJCtVXgOTi8QTWhNLoIGuBt9MPrStup98JYum0dvb2ieRnxTm5dzuLwnCmagB8jndN4mIZ4OyaK
ZjQsVEPAFcqUc0+KqBA/1HIJtzm8LyakF33n7yEvq/0nUgUv6vkxYvumIgDuxN3abg1DivN34ddX
wgyWKqywq2nO9poTmzJNx/a7TNmYdi7GemSrC3CuQ9HHjKso4tdI6mh91bYAd+Gz4XcDDh89PnhZ
fJDhpfx7TtWipd6KywB5DnVqJ0pmLZULaz6opl005pL5KFmtAWbWcA8XBsET22IQ0PA1ZUOEyLCQ
hBKeQUSHT+wHShkiuHGI4uOcFtXyulaCxnSXbqTenh9OJMHp4RxA2EAXJejViFhKGihkgtsZW8Zs
MMtpCV1ETz2ny/laLUQd0AcUSDKbyoZCy9y76CSja8SDjTocRHAFwxigM/b6NyPlh2rhSt+EHTyg
m8sP+cH10lYJzfHuu/dSXruW59XYBnukxTF2Efat5oKMOIFB0+k6YskoQBJb9Gr99SjgZYVeT2Av
NErGGUw4OVu0OixFg8LBt7IaZkIO8qO5t6hQmFp9VTdZk/JPlU4DvnRy1QGJ8clINXpX8Ng3X6pH
vD5wRxYoiuu3rJeiIlTIi4WfIeytiEIvjVdQVOMc2/kDtRpW8ALsS8sI5elJ8e3veH2vUXWJJc1d
Rxf2Vau22vztXn58eEdorJnsBIuRZZcj4YdqYvCQm5mrmwj7q3fJJmvOV73PDxD6UpHvHEDh/BZX
9munyD3TaqGQFvT93+WpBgZN1UQUBqS/D7pXc3f3gFO969gqOiyMl/GsEhI5vretw2fciKiqXD7g
H19e/RkOowEUxlwWPI2sZfTI75O1OJ8Xoc9PlMwFzYkJ94tjp/WlMSsKFlJYnnrHKri+X2Oiw3gn
zWya8A4kPifr1k/Ve56nOhI3x1rGSUgaC6Lu03rlI93G/XwDfSoqOAvwdMdUM3EMK/YFBpUwr9RJ
VNbudqy1knpSdcDEdv8EqRbs9GwJZmtgWpQkWHLJrOLCvEJmuwIk38i0vjwU7ZDmchQjZqMTPobz
dUoB3CD5ilDjy6w2UNnJKzzdus/1olhiNxq9NXd1TwK1lSZ/+6Kb9yffjtq+7yktwanx0WmbZik+
RhjmdnzeXn1F1EUXerx/FOzVxzQxL/NL744W7A74gKQs3NvZqUShUzx6CNJYav6+EVW5kw4J4Jh4
n7FjjaTeI+tKE1BdPuY1HHTSak9x34kDc9TIdAkK4SOHeNLUdtcUYBbCNDK5DGdqg4cHrZzqBoMs
bfdj8fxGcu/9pmsZk7IVZTQKWUsso5lBS5/uHnxH6J0CnOZy9qqJeRwim5sh/9lZJvFbyam64zAa
2fxo1Eh3ihcFdk2oE3J81rU6AiBeBhzHF9wfdct6vFl2MZ/CqPiGUEmq3Q96Dp6hb3x+ch8OKJ99
EtG1+xBh+d8fCRmC6OBUTWZ6zfz8ajagMcV/2zP0jOtlM3rVNj7n2SgR44Hl0cB9QqmrM/h8hsnT
Znlvn86io8FMB3RIfxYpxVyYgaJzgtwZq5FlMlW4PDHcjRVWlLCOmDGTEvNfX+O9ULW3W6JjqmAQ
d5tZmDD1BHVCWRCBSq7u+OJV14ua6BYvW0nP4GyQ4k/4cAUJGjBx4XFA2rAZeBZBXo2V/45YSkjI
EepV0qYJPq4dz4tJ9LH2oCp+uJT22oBXkjLh8Xgf6+K5VDr5fN2SXAypXzn/sZ2WgkFIOlaN1L6q
ctmU+lNxV/G15/V0GwFcZqvI+jsYOwKQZv6BbdDHHSoEi8EfsUjCzKtokwgr0P3CU6Tf3rQNuVX2
yXv5+4jCxLW8PurL8GNrZOAQm1zl3FOOv1SAhTmcSLvB/t5T+abYl3SDHOlKfdFrDL8xdSSzRvn5
T/xDnt88PKWqZYZshh21gn4tu46faoPmbsEKDmveYZyOosUmD1YsiJ7U5Wh3p71qeNwQnBA1JAoP
KDIMed/kiZnO5IXiSooI7kwvEp3tsMRImQM/QsH/c8G34+iB2TsAy5yy0oyGCvvYBHVd9MO+5QlY
O2fJSiw4MRu/ekA46rzbbSchB4dZJKT7kzID2lQIu8uiLusy1CuO3tmBX67uZvzp6AiojVxS8bAZ
/AK8TgpD/ZkC09fmmEyTp+jjBm8z1wHa+K+BddveztG+pGKGrJ8HKSuhrzl5GQv2wwb+3EH55wV3
Q0AVQYEjf+8LAn5RwAjiJG9M4fJHGWlxJZjwsY4lMUJ98jzGMjnBLbvgUoAO5PgI3LOSw7fZHgqY
HEpU5/lEFfe4H6bxdVuzte358K/4IAgqpY8s/zeuKJSiTCamB7w3ysuF1r5Tlqhn2h0fBCQyrKtj
Q5rVqly3bXC+IBUidhm3QNAIO01fDuioF1YK3B3mYuGC8oxF/YGhVMm8lOJDp5+5zbQbVK8KU7kh
xhsKRNZVgI0PSu6F1nwFFl/oJvjJRDgMU5qDcPpZg3quw4ZGXttU/m2H6JtpPzLnfI7GQOhULN6H
PSoISjwcRKrz14rOO0ket2XV4WrPOXodl/MmCwG+TEOuQkPfPp1Wxzbo2F5OuzwHN7yCYTagvBZt
R7OfvTPhWh/RYQ25DatWxYs3nTkXYz3kqeoC5N8NR8YtKbCzYfErNZV5GjST/iyTA9B/DgxSp4dD
7for/VU2YYn6JP2rLE+5uIevqhYJZhQ9Xek3qX6Vx8VpCgxQn3T0K6avxSfHVqN+0PAHx8j6CUXZ
j3jo/CNV0lojfz7veBakbZxcEbfRvxGFzcD6/N5Rzb9hBCoQO2Xnq4wXVZXlQDt58njXIwSqx9Ox
GfXteFVMP5YirdKwQYtXtV2Kgmmrhu9C68D6TidQG+R/Di5bo28RRc2IaYwc7Rnsc5rlkU0bAELp
e7UM7t4/kuhnfV+3w0EfrXCGes9beoiWiE1jcHKC+VYkjfQkhoU6DHDCj+7Dxp+iIALn08IYJ+lp
Ym4e6NCwJd/YANYA4xqFrlnnxcluLGtfXYfLm2xYsIyjUf8VuimZWov9Yo/4FluZSjgQAqeU8Lae
1uFma+6FboqS8i+uOZhDF9bcDA2/a5SmV80YYSqptW7DbqDjvQ5f1WTYeugtha/dsbemUTiYiQmd
Vr020RVGJcIUvwHpEJDp6/D+P1vOKjtAkfZixN6JVUD8QGn4XiCgVItmxnEx2ppTgkayT6hcptIN
QhYaN+c77q2r41Uv6UWwu6BUqF2lT3YEJJgOOVBuEPZICIp5gtMeVL/auJdM7YLJDarKvT4NDoAS
qQ84rqeYxRgpbTQGmoGALXwnKqmhQn+mR+OWQca28RMENfdI1K8oZ3NwfjMPzVRl9XDype5pNJm7
gzKudfJUHisojmKU7PyZW/e30GFv1obeUPZ71ySshCYDdJI9g9k1MV611i8414VMgme1k4ewbl3/
DVCegRQo35T4cEm9WNQc/PomVJ6w5ljfpMU93j/keL4P70NppvyG6ZMK8A3Vmr+GaMFtL1HOcepL
UXCs7zeXi7jqizT00OAAiTG4ZIZWfEV3fCuY+ETyU/0Gj4NPsAhI8bP7qH3AFfRC4JUhqBxrjBh6
EGhsRY7+H985Su8pbxiDECy6nD01RC0dxWUZS0+tJrUGXsV5l0/cBguxzYxg/jo1kGILguwcf+NU
TayWODWXCIDS/Jpenb4zfzZUo7YX6/HQGndGKNz9q9Y64eSag9xtgL1UWjy7aiCNvlRCcLQ4+cmU
4XFpMRS7guD7To7GuBP02u7zqClBf9D+aYVkVHC9eiNJz+rLZIwINFRNVZ0g5qNxeT5wn2rF3uUh
TXx6ZsvHXLAIqGk9VRShUZjvbQbYZK1/+W6L+RwDPhKeOfoEw6vQgrFaQfgovcOfIOiPZuBCwFTf
vg6IWf8JudYIaKusdb0gtkGUohApWZhVH5vk7XgPfBaKX31a7skXW77um2B30tkdJtJMOeNrZ1Nm
TrH0v1UMpRyD5w65udZxPVPCJSK3QqZj9QZa9jSJ6vBnlUHl8/0y7gi4aqAFOhF+oUEUyxT6QKkL
ecFEXaIR5Hj+9doS2IVIFG8NntKTB66ZnfhudA5cKinyAKt4cSSEhE8mdhYUI2VDb3u6Qe505Kp+
uF7V2vuNztsyN3qfLGazrg/OKYPw/RqeYX6ZSgelvyiYa123X4kI5NyZSd1l9gfK8UjEHRhd2tVx
kVGbR6/A5s/526tCuRyr+H46ApqVMtHdaU1Tnor7cGlV6NJZ12LEkh2Bsyvabr/RuHNr4IOgqBzY
pWhV5Yj/AouU6H4UAIA9Yt4kBn3SNvxC+4HkYGYHjqfyo0Xcg9OzLEQhK0LbS2PAIsbgCSFsNnXw
djI4yhAYoe806niYyHZwuAJl1iXK1d8eMuV7MeaEdSNyVSzivjNdT+AZVjtZEtO7a5uL+gGD4xrz
WslmGRaBW0g/QXCQmbBiPkW4PQefFxB6psA4HEOjMz2zH3fSUhLqS/W8QtlR/UZlyZ3OeotdCRdT
AaOW8en/u2KffhEGCZByCOMhEo7VGDz5AOxZoWTXNh0HrSJulz9oLqSQDm953gXNFzByza/DSwd0
rL0gNyIMOP9zXfrZkzZzTZ3VLs14Cef9npLIuzBwquLfF8Zzn2g7kyCZHqa50zzn/+1J4W859fR2
PI8H6vbluY43UaD9BldmO87qeKrvhJz8i25nYmMB4THe9HgoJv4gHnE5EUii8p5NVs3oCACKScSB
X+nF0z52WJrn8BZ3leALgQPIrzdKBaezBV1REFSamW/TQFvoCzdn2CZ2WIzFEHJoGEPWGAAn3JS0
7TXpUP5eWaIe1Ivihx/GuEjeRb+NcGszi9iHbPyJb7tXDrONgP5uhfl1xROPcRSFENeL65drkMvv
oQ6BGWqwLRzSdObdo7teAdMnMuCKcjQV+uDA2wnd5OoByaTsk99M0vx1W7HMROc7ix9M2JOhBRkl
RS6oMioQE9HaNA5EqnObgX/9/6HfMExNh1Q9L2z09B1ALCdy3tRBZU8k6A9njr41luEqqPcBhaA/
olTOWvFARwtSNV3+2jD7j9ghNc9TgT+w3FD1HBoptWsIc1Xk8on0Bvfo5ifQ6tiseQQr/n35kHaF
Wm4F167KJqUXUmmUlHIwAgZg/BNq5XaDByMQxDzkldFqbtlxXJ4peFbWVU/zPpMC4NPSPju2VAJX
mfmUE1Ti6HJl5sWBLg+BMhr32X14jrFHqvDrGqmCi4V9FMFizTAv+8+5XSPNYaNRer66Edo61oDN
e5cdhgLBq5dHmgVPM5R8fjjS8sHRnps42XF1zgXed+/I6o1mqHpTySOTuavWcS+3EtIFm7Nwb398
uVd/kChw/8Tms2GWr3uubuB0hBKVooqwOxkwRn38eruLEpgY4683rXTgPOoT+y2GynHZlc14FRdn
vvcHzZdKE+RDr0LlHbMkpCRGW1+4yMSp7qyxMgXY9fLYTHBVxOPb4WYYUn3yUnK+AoJHvwoIbjIc
yjgr+A9KvbIy0bICCfmhHzGvgce7tyVhIWT7qkXVm/98VqNn3sFsUH4NaCw1H2iLXKPIOUn9J92o
chPDe2aasIlWSaQHy2YDqsuu2o/xDvehd0sQOrkndn+Q8nLWUKwpxV8HRnIDFdVSjTzkzA8JLTzb
hS/XEr5R3QOOj/Uunpu5K8vRT+4mV2sVAzAv4fep7TZIv+p1jhOlBt9fvzDdiWuXqWNPZfsMqfMb
UjKt1nxzTAXVAwrPYSkML5FpNDBp5brMit1IQ2PvqciSL2rNAD5kxEIHMbUzYoZIjAWXj+heBZzx
Lsk3jZEbbLy1sOWiRO/6zQjgbC6Jt6xKEO3CTYtWGjj2EtuwBXwT8aOK2c3pYDZT5G3YteyC5LC+
0sIuYG8hqqGW/ZankGg/fJuypHy5m6p2iMp0LmQaQBxs/j3X4NqjdrNAA4GqCcRAyuGjr946ONKC
h3czSDolGyTX5Yn7555frqhnizEWhlWmQT+6HGjgZX/40AAiI8M7TiMosNtbjhjr3WCl3n0U8dP6
8kLbTZ+UFss7vZnQs4a/uckWvUs2KIgYf9BdUuPJdHl0CUjoKNAxxs/ztWBq2Chq9IOP+ASj0nFo
72gw/yIzrlFNvRlbQ9Bz8kW3HzS1kG0gZuigPFMV1KNj7ilUuR9+XxJuFlAoqsjIAq3/h190PIWA
f1uyDsT2+J0C9C31HE24hzRHkTTCHVCz2A9WBMNihOCgEcKUg2x3sNYT4ZMxBd6/OSYMWWaModx/
S9ZShIf51/400Qs3xuQHEPrBnAHihEXLMoGgT7C8vqQiUG4eZTz1ciB+fXrrxMRXF1vC20gTIxaP
Lwuw5R+HpxHz8580DJN9gyvU8u2Ia+O/2gLbJZk/BVVqOiwxToI/6PP25c9BU3K+crEfK4Jl+bR9
jjZcSrLG0/7ZT+6rMyhddNRpDOjgmNZZV23cLKnCytgS/TRMwGZxe1KVdM6UkSs9kKy/VEuS1G4C
ecKsSGWKcnganBSEQxd0DEPNltYw/m67vY9+KyHDgNsOcoyXLP95YgJ6zkLl3ngRdwQBsFN4F2xJ
UflcxzGEgMw8Yy4OcS7BJSNlRISA8R8nT6BaMa0ElvDGQTHjBNHD87Qn0XBRQYWtv0Bp8XQAfji4
yIwPzZJwRm+GGBsfN5W3Eg5iR6S2uG57m1IONO1MRwubfHTBf8evwipEsnmHS4aoETvH5Gq6jIvj
vTWbCU4PsttR+iUZ9bCD9lAJreH9GeiO/BvdC0jsuoKCvzq4W+GmXEXvOzHF/U+hsaN6ysDhtbKN
RmGbBG1HvGZy1MZ/G1JPH8FoDR6Pg2xIfPYZCLm/r+lD+BxJ+EuHVzRZEh7DK5UB+Xe9CiLUY4BG
09vHmy77thaCZfNqwsrVq9NuMNT/QB/7OcPFe/APeurvkGcJfLkaCVdgWEqs6TacXKIxm8daB+oO
lB8261Imu7HW0pBfGZX1Xgn2YaIpmEudM5Y+mCMTD2BFe+xjSzquL+ToY5Gb7kZgPdPIY9e+K/jd
YMfhyODziREe0WKXwY5LoPfDQ3dTp1fBDMrCYUnl+oGCF3ptDSJzKBXJ6fxqykZ6IP6GnmXw2GF5
BYI+23tA1z/vwrmtX+A2483TgTomRBBOe+2Et4YT4nGSzvZ1JzpKSPnuvX9N0NbzH08EE8yQMLb4
lHdDBRkKFDhxSFW39siEyO5Gc44RdYUdP+wQ6NDSZ9sV6kctAJmSkALUFWsr3aW86kqC+iVBNCuJ
hzhlM/PNCeC6o/DXKVLwQxez/XY3NxlN2IPKdfLLGuD9EYT5IACFvc5Pyw39swzCK+5XbApVnZt3
+g3LYZT28cwNY2cPFmjdkfiP4iHgORo/8QhyyFFfu5Rk1m2i0/KzAVEuVzrfSzNXjnOv6ZsOgXVe
nPPEVJSgY/72obAc4VZXA+VzEWkQK7p3I4wjvX0D3y0v16KyYQBRA1UtZUJdWx7mYLwFNLoVESVP
on+r3gGodk/hu8VwTaUsWcYP52KZf33rQNYBlan8DTDbvHEHtqZ38QWLE1qdAWt8VmcBACYn3zaw
OvrlbNrbr92QTzudCSwjRUFbpQExiN4BAjBP+OfoFcPjb49SWc6qbw9A2P9hvln2ZbV0L5GK4fEQ
4Yk9yWGPttWNL8iXD00Y0oYIynf4zax1vfhPkyCW3g7Ow2Zep+jE9EgzG63Chm5Vpzt+9Cal76VV
A9/AF0FryA4h6SZVncLfSGEFhouIiSonasWV8mv7CiZdbQM+JEli2bNagwmNWmZBvrD+9hN52/o1
UkCZllaKlJLslDsqTtWp1xg5MGF0Yv6PkAns9OIqORk8WXorafgprZBseQtK/qSB1/WdpsISiQ+h
pnp9JhIRaDE0ufOCeoK2ajOa5Lx1MY+CuVbDrXem+8Beh5d/RCApbmOvHHOXE8qOfR7FWWkYFBN2
O6ucfaZe7LEL1ryHRgO0jsBDqBWwIA4FUqQkP5rXCFhqMOA/HWPWpTrFDtIoZw52JflZhXuex2l/
H9Dy45a1Dezr4YtTTS4Qk8KFQ5SzPUUVZ+YzdLc+hSGMVsioHw+q/x7Jso/iQVUDVT/CnLCm53QL
uMgjzPCxWuQKhh13o05SwLmHMzWymnkVjiVSWcjPpqDG6vMVQG7BUEsQCkPcaHL8FyVhwv66S2VW
sZ1VaTIbkg==
`protect end_protected

