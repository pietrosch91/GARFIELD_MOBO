

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QHA3Ex+CmcwhHYj/Cu3wGvj9D2Oh5X/PuqFEaH2NXNQZh8T+UDvbmRy04SPk/2ZNtGxTEFpvVC+A
OCZnLDmVBA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EpCFyIVFCjVsV8JAoVIvFxgMicPOE+gA797pZe0ptQ+JWzBRfe+ko7I0AJCcVXyK67/23E/Rmn28
26K0nfbqlZMWRo08GQzdo2Pvg+0zdb5xynhVYesyBJF810yAmWPUXibisA0Uz4hy5us4urGRvXui
1VlpuDGRFz8HEMlbkMQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H91qDFpDLhLKyu2zO0jS/sr50G0AneZOioO9iB+qoJcFLnwgo0vpwwtqzJX6wbDVN15cu+R/IWxt
dEt2vBf8d1vLuMo7BshJZtbUM8fTrhTZcFoSdUQSe1qC2oLTy/DpceJuEMWuDApMg7w81zUOWyVZ
l0ZQx93l6uEMApiR26abzikEl3AMNYgld7204pP+LGkuQpEm5BNdhJ2R1igYEH2SLr9PoNXl6Ybr
Jw60dHycu/SF1aZZvyjj/k0RqWzkWo9OF2bMBdwweatK0hL4Za0tR1dkbQIVANMFXr81aRAsb+LC
ySA4CauSi00Vi5Uc9EthY+ZLgX5Ay9HkzjDp/A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UQgJtyN6NYDXy0tjNwGtkb8soUmLxZJVzWlNkhMS/C4JfTEXUPg+A6vy121UgFOz3JMSNyezviZf
Mfex2hTID+DH3Y/f+mS9lvkRe2ugr1UrbCWMuo61hHhoeO3FlSVy5OojiRVr0pFZAlcHpyRyAMDC
2ubNAtCqnKhJ4O0W2nXkasQr4eFt+GOK6JSg9BIu0PcXYnr8Z96U14IqU8qoaCFnjmOffa4iFoKt
fCItpLPWXVs7vpK32UsZ6CdWATv1DRVa7rvpoKAYhB3pTdLEGiZwBFovoFut6DljSNKFNe31ZoBh
ZvEnbvlCLpTfwwRuxQIxsF7NsbghGxInSwNF7w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLlPz8clXjBHUAybAGhYboHKfTw7ps5cfHItKbfGW0Maog/3BI94ghpter+alXbAkH+8KTGFy2Ck
42pN270kZeA0uP8+FP5FX9Hdxx1rjSJSYnLaETC59zrF0zNRHR2eUpWdzjk3Q0IyjEcI0hzDMWpB
BTUA2W+6VKIt7CwOChCNccifqqqM2/lE7U6SRri20DGmnKYCeA4SLYKMVgbYiwIQ1WpXXJqIDpo1
bsC7dc9a1YP5bjwk8u1LIhPncODSxREUNUwGR1Xb9he8Nu6GvsazhQaKR+ckU3zv9ioeFohkv8YC
6S+WxXXst2ppErBUJHaQ9VRsWjop1VaIGfPf6Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NOuQSwyLor/NCRAPbb+hLF/fWkzD7blUj5CmRCbO6PxyE6eUcw2hCJ3syd0WNFx3AwuOr2lG8SgF
2djEMbP+862p4gxkXmmNOf7tGqVDHgC/fgmOIsxfkZ95hvRAcEvi1RVx++fS0h6KGuC39yN9BrTt
nmZ8JjVs3v/ky9THrn4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BP26diD8XpcagtcJpVVq+RbpugiTQYYy381rJIl+lewz0g2oe3rZrSn4SemKHDAtULgIN2oNIFYj
pWqaeK5KLTW0n4xvkxIsB7rciQ726nTjcRddBUmvF25tkhA3Y3UhvL2S3bElyqF4lCnStpJABIFq
XT3R+Lyq40nBC3EXTPszZosjTkHBl3uO8EFhwXxLaoSimXXGgappLzUn6dp03J+zr78NjVyMcx18
lwiud2D8+5QyO+QXigVTSDyD/Zd1vaDmZ5CVwxsypJWCKZ2A3qx4HCL5RoXw/1eLwI03EXKqEgVE
P4uFzHRwLGNImIZpDLhj8SnU8I0lOUFiGGuDRg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132672)
`protect data_block
uKaqaRXQqd4cspUcT2rcerrIup6sCeNG9Gb9ovyNUKiUbb9aKezIynlvaIkPfPA6SPIp5TEG/RoT
C0ZGOLmsVQMgk3d6TO8cRbGOCjzaRTPyJbIFwPjlGIAKJORPEKMQ22Nl4chGnaRLcxtPQtYEMqYn
s6DDNYXA0KyQDX46Cy9bkX3O3DLLBsnkCH/N+nv9taFnMCBqxe9dozzj/WI0ETK73+DBxSiqzpSz
k6m24DS6ty6Jke38Px5mmqEp2ALWHGpYqKlgDQqKLGQTlKau/ReSj261RUceIw95PQCypb/TDpHG
d0DvLrJerNF3fcMddYpS0A5cjemSI1eijcmiOInJS6ECiJJWFuo+CiRPeYN+gWiK2tmSli39Azj1
sLv+sLfZFm16DnqCu0b0tPHCreM0tIBq399tMG53C7WNNimDr99pftPXHPni6l9gaU5ahj+gcDio
QwXgGdLozZ/DVR3aqFpWATVesGIrvQpV9ehtHM+57Fx03IzCFBbHmPjMBkhEtzLPVU6P1+5EQFpz
WOat8fixhkzztgvpZ8oJq3+ZwxLqjGHZNP7GBH0TAt+L1xi9kpjyQDSnitkGHY/PlWbJwMkWVjLu
hB3m+Qyq/OJcPt5y0WwxM2AGqCf9Ch5pj4yI808q/R+bkrisTduwuE3ey2PfVeFKthyp+S7y6xNv
nVh1JQjjUQSsgl+yzOHI1lYWDVO0CTMo+k+N0RTyigq1HVPHnD5xqjbJc/o7QwYT6zqqo53+FKMx
g9k59pQB6jQ8SUhD1DrQRSELSgUFeA+gYCeTKKeU/6A8z5bzApNYbYDuR4dm36ZjB1jOJ5aawbei
MQNNaK8Xsgq0d0Ldq65/aH8OGJ6bgCTjojyDvdwMVwPAvtwfhYxIPsaf0wRxHYgwFcTZ7tuvbzP9
D458eEPdS6NGj8ekW6URnoojJM+D4eD06WROhN1oJl1dEoKUcsQ5LC5LD2Gfwcgquu8wANMAqhfS
j+4jCApjtpZ3qWIIDn47Nn9thd8pxQOs/PWyfGVdnw39Y+wxukeeACgnNGbOhXQ70HKLcSkwwt55
9t3CcKI7GttGGeBH0nS5WejY1wYTr2gsPdyogiNZh3AkIi8FdoMXJS+HHULkFDljpo40RpEmwaWq
EdrKpFQiWijxi5t8dH6nvWEXC0emUSB8zQKOP3EHscYrKw6AqrnXIzCf3Qb9FRjrOWCbDBjQV9kt
BChr8panFjJYHeTYHkuYVTetPd2lr+khtKRhBoUio0lb2K/e2Wq/88DiDv6B3f+cc3OWAiOINEt3
QpZ2hTgjhQ23+2+6Vlz7In2SO8ynCwxbETP9aBD6V6y6ieawHNm8eVeBa0eGSr/0yBwOdIGXSIXM
Vjx9WOwSgWVWbmKw82EA6eWP1E8GTOWzWwynaCBBKT8bZw1VXeq9RBryQ9AZ5VgGXWCHJqNyUdJQ
USRypsT/70xKKgXIXQjW3Fi/7YZz3E6dNH85LcfcJotXLrmBuXEHtuyGgmTKjN8NL92mRJyuecIq
wEwYI3zg3YoulMR+pCp7SCvJyQvi+0GObRT6uAgcM3EQqIaD0BmgPiTwnlVbNhWMJM28Cdh1Cr6a
HavLG2iIXHN9FJpzQNky2LQ1CFI+XKWNbreHkuK/D+7ttBoXxWk2QALGL30UPQHFuAdnVFQngwIK
ecY+a3jDUGQ0Bb0B6cDNOgDbrhAhqCDW87m1qBIYsSMkF4uwn1tg4Lzkfh9gz7+N5rXp6rh+P3ro
S89fFp1XDHd3idN+fvhStf8939FcGrG9s0Z0ClaHB46KHbESHr0/k7F3Ybmocv6Sp+MeaacdFy+p
S63Av810gKN2S4O8LrOe4/2m+uSFyC/IJk+xhhQs5VNmTV3l+XsM8+uP5LnEuohuPTeAwM6wCCIe
L2Ls06PEvXJtINUkbk/olRL+vvUhTRBtqMGnoMd8EI70Lx2XX25ZDeGzwdnfPbrVGoHsTTiluZxb
KUXc7+AMJY7eAcy8UosFoLMePMhf1TcsSjCTOakmhTlcxAOluV78HKJ1y62DZgSDQQE/WXX67slx
48zx1xEG9qKTa8qNoNpcBL2y4eTA0Ndh9uqEo+sLzAIE971KN8LnffIGdbvvc8AXxSxDYpQUB+Tf
KMjG/El9pT0wM7B3/aehiVtekLPzdK4JrsF8E6LFoRRtgfX7Wu6j6hdS/HFQFi8wx8YtZ1t9ES3T
mD0rqGYlRYYvEyszA2sFfk55FGGRepldEIytWl7ITNYVf1CxFaob+5wNFApNDt8Er4HzywV2p+91
4w4B9gMT+nZZqsWD/l3r1CujiYaObwXw/Xmzr5gpkqFcr9vst5xOmnhruJaOvub6OjqQuy8xl+I/
2RQnajipeyZhGsmdA4v11R9gljBuRytP1Vqly9/vvWiiXb53XIckkGgO+ENGVt/nzDUswTBconTU
yIXoi0cFBGSfHziTqsmMaHhM6zNX2NqCOUe1Z5/rORl5kbIomH7cx5w8sRSOt7WXVwF6ziKQslAC
r+VYi5JlfZyshNp74tV/33p3rl/ewru0NPNSRtKNe0BmeTZPmSeu6n9AughR9MEOaLp63v4y/IRY
5HKQrL98NiI596B/LJsIptSKEzkJOEyPKV9JboqwgNyDaPljG1X60R8yyh/le9nwQaoYRjaRG/Ug
JzNfXF2b8TzJXLymXJ0otpc8mEuK5fo4boluduvaU7WPAxPohvDfHAaWKhTzfTHT9faxhzt/Fc6L
XtjhJI/DeG2MzFd9kxyls47CSl2ncSmwRZbEl5BDEcu22KTRWZsZmuleKLAvDH/w59LOYLZxf3IW
6VIlpDz/f9Bml27e8yy362gdnRxFbnRBesvLirdegHS1g/TWG2/Q/KB1bc/u6pHfcPxFXK819Gg0
IKj2NzcQLRPOtLmTVeWzi9J122BPhM7togFZlDVPy0koHdjbGFhnGD7+ByVYigW/Y8o/wvWrUgjg
4NEdEoiph/aYEoSuK5lEiCo6kSs9goZ6bAwrETLbQSWavY68n35sYqRLm6pKdOFR+bbT1s+tSZHz
KYGGdvEFwRRwcF3iFj6MI+JB4+WHx5zEkSs174+2fdZ6m4bcH+JkEKXmIUAk0ajMJBuSwxAocRs9
NkdUENf28ghs08QaSqJ6wpOFoMO75PnKSgUP+b0wFlCQt9G10mkmTSZhldzU6MCox07IvYNByfWw
UrxjNfVzUh1rVwSevlo65lYc6J4x1uCitSCyAjhgTx2XW6Hr6mNcDO1QY0PVGp/g7YqzauhJKe5d
N4HZoU1qhrpledNXDyqVWTRs1lF6My5xhhDxZMtqbrcYQqsGdlvY6YQdx5cKpx9Qyc+/WNAA+G4y
IKKa03biYt4DO/4Jq+5ApaIgGtMZqhBNF3VtxE8A4Hw5yCsPz0CpayylQZQRO4vJnGGH85sXqBy8
4fKsEPP+ykrFvOVBrBVIYyFON3j4Tllci6xVR9ZjyUr9AUk6s8Oznrg0KGELZmoy2oNGKPXjgfby
te9epq+ViXYubjGTFSSCrAKTa5pL1weSbRX5pz5KmBP4N/hAnBBAB2AvQFaEPRpnu65Pwt00jzqA
ffByAIxB8CnGkCqTRCAQKoyfu3ZNaFEZmwVvxeHPtMjNOCrGp6Ihxrn28HGuHYT5P5nL0JsEhf9I
w5LMnOMYU6nZyJxFI8FwA4WjepVb19gFEdOc6RR0+Pz45V82v7t3A2snbTUMxVnp4pT3nZJzy9Jc
2N6kPuZfnTJ3A1HfzVtCLC0pxmiQWRUIGSexca/DKD6hi/b4xXm/HMpCArjizNrDv49Eb1+ffd5M
LhPvZ71yNBRnwlEy2zVlto96p1UvydhDQ16IvBEFk3grbxNmyDX2xVLgq4YGJNxO0wmci/ol7qSi
T80knOIfhK9GPa68GEqg2eDHZQu/IEaN84IhQTYKO1Re04sl1c515vkgbkkOr9TBOtoiV8EBdoXL
9JYawBlfdaMPWpvBmp1BydQ0DVUrbD2hz8EN2W9uI7lXL35ZpL/QjplxC5FciRfe/g6PsNswK2xS
tuni7a/JluAkbX16kKW59xSf+62myLqMWEGZZLlZ+uhyAyhnkXLTpq1gJAHgDhhO+sa5veIz8y0T
X7iE2LTb7QlHT/+GUhrCej62fctCT86aR8c0r28KSbT9O4KKVpuwRN+rlrMa8fp6VUiHZpo+ctyG
e1CHgq9GGPKXyqjxh4gY+L9TIXT6N9+eR5yE3ZGo08s70HJ6mcLFB1w5A/TPrxGwsOk7dfnGRWnf
TTQrISTh7VidOS7wWFubYFcb1s3urRkgOK+qnhk6HAf4zzUPBg/oZtibE5IoUQRnKQwbMkAHgDNU
4LxVpgPNIE8EzqAAPuQGuTqhDIF2Rzz2v1uuRaAO/ojNk6fMA01SYJIR5fXfdwpNNz0CHkFhwGDf
5Q8qb6zvX0ZbsrJINF0myOAcMWweIHMG0AkhZeJspb8sPP/2XXy75wjNl+mjFzNlpBr8uCzZX9GT
Bnbursa8WE5qtEJj8Odp8VHwt99vZ6e2H7pulK3jskDWDOom6GquY6IQq7XPP+uKSJE+9OsOBNo0
+l20K+J7dtQtIQMi1goV0HN46EZ+qd0FsKdlRzBTfHekZw33AwIFVqI2qv6rgVzV6QDiPZ+zabmY
d8tgG76VT7UwKMfTAephfgYcsUS2Puq7OAKcyUpl7bHokhJ2HlBDqmFHPVN7SRaVe+2/k+mp+qgW
BVR+iW7eeuLN5ynj6SA+cQjWVbwueTXD4takQNHkfzVggb6aF6Jes2Y+gdgv+krOqh6khM8utDK/
YwsjacD9J1nszfcRaVagwdYJJONFYopLSZYjaxJb8bIVw9myI44Je6IYPV/Uj8WbEf++Qg6D8acw
c5PbEJiwpQGvIQSnGOdLJx4/CbS3r24xx7LxjNFmogV7eWiCSJM0hvaEv3JbkcoBvJF1oaayETwd
NyWDPHqMAeJJmwemtyCA5KUewvuE0+OF/gbphDwIJC+e+N8FUmdM4jVHsxZv56lvrG2n0VMOg0un
NG3f7rTHb1Bf/fZWMWntodoqplQ3pmmgJ6zpTTh+8ns+O3zgJXTl3OZFENp0bu1nEDPbugcUFJ3e
nmVYkwxJpa+GOddWYEBJjl2gqqnsueB1LOrZQ1zM6pSDGflXCVtIp4uO/OM3j+JZ7cAoEa76Gkjz
wZvPrBQWBqDHmXf9N/j9kLpAURsDC/W0vO4du2mZMv2ZAXvQz48/Bc+uQEM9q1KyltpODZE9Tdgh
LsJ8DescahOkFZZRWMfNA9qpr4LM7R7owRfdtkoLWSWxmHFKtA309g+MmipBCLOgSgFGlePivZmP
ubxvFrg7FywubJc6wQoJ+/TjReqvrL08c3Bp1XoFNM0BbuVKLi1Cul9zAEyy4C+wX0o9mNnvQqmy
yedy5sBnvdPutQO3+YKiHsNJTcoiqIG2jdpQtqPvX5zzqlWuQJJzoAk5MlO5lupmB3Wdl8PGmBc1
dbdK7WbeAMCfF8A1HkyrRMZ+6Dguw6OcYTUW5bR+O1eFIAXUg7VjV5ZdFfmlz/uTqqtzrzstWbtU
P9GveM5sz4CJXu5MlAHc6OrFuR3LHM5B50ceU+X0Y5NsyamhoJcOjLid1yRtSqOupcRAeLQukq44
oych7FIwevMD/KdYASVS/KcJ2hWElk6oS7J5LTx45J/EAA/m+9f7nD0pTbI6QfY9HJV2FwzEGNw4
zODejhBSG0fzt7hSturLGUWwZiiN7s47p3BFG7UnKVWglh6HpzcKGGFvCndRXIrf9BfSYp7IGg+X
uOsFPHeLqh0fAd0d1KnjnuXBvDjJFCnX5ZTQ/3s81M/WlCwbyUsgOIPlX8Dag1hY7Z3Sd8+8yr/x
VlrpquJy4DRW9y54vUR+UehiW5jLSSncCtpkeiP6OanPfeWzuS2vZY+6BcVO1b5SE1K5sdc5P3Of
N1hQSn30DluGP1K+vo+msC2W4coFhurBaulVJN2GzbANSYmu9fC+ZQJXyjjxuhj+OyqmgrM4qTK5
1OGvlMUqSCc6DcW14CvAJDNUjv9bYXXPNMmrIVOJ8bookmJsdRfMvCHvA16VVYWl4PGZnRPi0Sx4
Dvu6RUw6iIjT7rpz0hJiAL8FKx0/TxA7TzFxSlN5ynxl1FLf5d60sOJQbEFmY6O/x48NoD5revne
z6By8WgZ7Km4bkNKAEfRmXSzPOCF/cvc+I+QBY/h57F/b1tKWyGJmvnzHGgswTYAzubl9Hcwdb7q
P0/IlEtA8DkRdappwBIHyN9u1ah77Qeyzr5vSO3dO0GU+XQb6cGYBvs5qBkzysUpmiFIe7I4iwNr
mGHHD05sbzyGTiHbUTUfqg1t7B+H7jVUUuLvoB8rFaMz32CTpU4cus3TK/U1gV4xhmz7sGihg7vi
zpwgjpp3STWt8YUzQasYb/9Doy1da7tlx30pLtHriBf9P2UExwhBxma+5qSv/vDVei6GlblTUeLx
PRSZTD6vouvpS74ijbu5N2rOdrAg13/MRPC2Ai3FpKRskzRUu2ECTfjX5OzPxRMIE77JbX5LGqCp
+EixqQ9CQ4VHheQLN8dxUwZWpNKfSdtgt2JkQGLTyM4ExhnEBUjVMdGB8BqjlkH/yfFBGHGYf1O7
31lN08cZ+6mO5zHCs4EWR8Wrjk7AP21DeOo1gBdn8UKQHD7fBXnbtUduT6JgmDo2cNmB9kQYyBL9
4Fnt7kbYWhJexKI+d3Ix00xm8b524Z+37NBXERwHOnqi8Bum2a8UB21EYK38NwbysynqgldhlbgV
3vwj3zZEf36Qvn6mP/EXqgFHMaqXqarECijpB9mc6PxQXwBGUBFPJW28soBE/mqk29tQ0SxWmkPd
btImXlm46oU9+zQVX5kvFOdXj95yK2ZNnTPt9aeo9wSBxl3FYT15wMd1d3RNIU1nWs78dRmc8bGV
Wskbr+NTjZeyWRDHJXH1M9ZDm3qTsbbJdzpMNqQMp966NSFUQuEPNRT3q0vc/npbUAw1m8KisZbe
xeZeK1wBDRMnickIumsbACvBRw0MS3aSkyFz2ETUYPCHDgs4a3FRSjvEBL5wfnIE1o2PodYaw2w9
4WBz6dNmlsbEtMgzYAoKS8nFkV/dMWA+9zM8mli5pTjUykvpIJCUp/qVjB4PU2jPj71y1RhB79cw
R/2PMlf3MbRIO2XeIOVK9rFe70EOuLiYnveebPhGmK7lk6uibXG117uc/M0nxoj1f5HQNHB+JA1x
2VhhnAMm6mxRkLi5JITApw1QZRAzFl0r3kYJEgmbc4GeiP5Xy6HUtwnE8eGT++OQGTFSxMve8Frl
fKOELXHs8hBpvP6zDslAcQk6rGMMq2LkuSUiVi5VurHmvyg3IPGoZ5v2gs5DhELU6dLKZS7wQrWv
JKwPbHsFhhV7xh7IN/QRMYhHfWDtQA0SNjP4a6OhIu0jmxwqH6aNnSrUZnaDT8AZ0RbLn/9nF3j4
alWmjbpn9Aj7w1sYLC6Nz7GAsuCrbB9OjlOXqGus6S0BKwDuKBYMhO5tggS5/TQo69tAZ6QIvsSD
QYZdH9cKVjx/fgnS5SfYNDS+7Nf126xOaXnAolHnscQTweNNVNjFxiNKk/YQ9L7RV8S45VHRMVww
blAT3QJG7qaRm+NRaSI6dJQ/RxzoQc93Awgo2YYNCctLVgdbewbV4igzsfY40ef/Anky91Xkq5D6
oGHY2P0cesyFVXqXx2hvk81pUT7ZDQ5tj2eVySi4LivGoD0SLqIxs6wuJIsE9roqol3BC6Q016yc
JG85qqTT2m8VJianmfxqNOT+dYDSvE/QWdeJTR7h3ihHUqqOlYo5voLjfy3S9qJnSwl5ECgthbeR
kPaQSeRfj4dHLT4z8E1RWf6Y3WAaUX6wKK7/XzNV1Doxc9MSdUJUQ2X1iqiM84Qq8dFCjSKMDBmZ
0jL9HGi7yofHB43IholSGxhl/t4p6QAcRDMHCZTbLV+0S/57XzxUq+gqwu5DJAhHaJ8xVhBXlrVU
XvxoUPALp4BPIW1NQF31iAKGP918IiVTQFjDlHTjD33seqEE+Drjnt7Szm8MvVjYrh9XVu7O/hmb
x6xLXy5SMWOEmNsjx674uo5xN0WaFkucn9z6Yf1JilyqZQyK90TXzBgKyAVnobnZs/7hkER84GiQ
X72aHRp0rtJtQUA3gKOcyy+VtR+2Zl0tzw9BcM6YTzUQR3/PjSDonNCLabnMVBRnDCHldOM7udPf
xqBwnBjwvG/fKmaI2ZvRqOzJUo3Ep3mT6dik2l+/hOAjekSW/OaLkyUVlkxo2CZvWvekmRVret1T
yziwGP6RdZU9YJfWRx/ckDgIKVd+c5aR2hzcnhBXzRvcT2FWeJGE6k75KWOrLcSwNZslh4JLRLhv
38aYx0iyzPaRKMekpLeWd2/AWaNMNIMFN7iTRW17H3L0QAF6d8UsOSSDiWnZnBOAHiU599QKTgJX
YeQeNJw98jTQbLzQPwbl9vsUkfy1/FgTSpF2mmOtCZTtTmNkH42OYGIoM8X41jVsbVPTgxWZVWpj
ZkIL1PDh0KjpusCzZUa/I3xOuxEMDCTAUp18xiZ8JJvOkOwbrKvkptQWwONhfJVtYhP/REE1hJDl
6nh5MqPUjTNEBA3yNYc0BfZoShC/3pGy0TgthoVIMWNkZcojbca+FvfdFO/Ecy1rk4TUML2PRfVd
E7TwC19hi34UOwOa3Wa6KIGLKsPwDOsx/w7Y+0+NPoIDz/k7tKhur88ieNYsojjR1l8GPv0osFDl
w5lHFijdRoOE65O4s9mG7Tdm6f0BdSKIRLkcH7SuRCZl9UW91C2dusnUjx+w4EvsAv1SsLrRkm7L
5m+jFYLr+bXEViWl6x5Dj/XQc5jYOpgUnlCXlBaglQYi61HpMx0Txjx5dCredYWN5CaEDzyorgyk
uzEo8DDtn0bAqqew9a0qIlrhgh5QO38cmLHBhuy5XvWvQHr6wHStIQ8HNpPCArpuWpptBxenNLJV
ZXU5VAlde7waCvO5yDYztME8p722ludkS0OFXFO3siAeKKFNXg01xcSjL0KzqP5n2pH1C8zqwHTE
24Hfi8lF813o+ekBUQ3BAgA+Aoygcham38oirCwwj7xdS9f4ONEjIuTEFgBeR6G2wdnSeODmnF36
OLT7wBN3cQTCBVw/Q4V/N4yETcK1UtJpmBwalF9ZZ8EZ9DIpB7ug1BOVJ3/ldKG1j0RImwc+xJns
6WEktx6ZA//3wWEpHHStyZ/O1KxDDoFHOfb8/KyK3Nb39nGFKhUgerNS82VaM9h0FUBhIfd0E7fI
tL78CEMdbVOA1gyhXyO1aUShaOYLMwoJzMXQrmKCKaTDXTHtu0Y8v9cn6IfhXNtqKNDLN9lxWhKM
HAnIcUpNTJ/BVtSstig1tqT+l7BUAps9QSTZ6TxceT8kqNGiN1ojlU6K/RWgJ1P25SckVTYCbLRK
uheCS7bs3J3GkruAlrrS1eHNCr9nob6DClABODnkpwmLc0qW+nKdwuWgBVB3h+rKJ1lR9/Hf4/yq
4768I7PqEPRv1wD4m0cLXyomjeIX3GPut/rUtd79Yr0XSzTblxFWoj2+/O356IqorY4L3+mbJhvn
Bjqh3r4gBD7BUByjHBa5rNYSdGpUZIaFpVwz10kx1eLjy28BLUN8viX5PBkoRNQw1GbNuW6llP0o
0Xp0/9rWPLtjPh4O6Zv52kc0UWWNiz7ZPJ/0FbNlTF7xhR4Z/FHk1l9LuuRcv/PIxmp8snCFbJig
nszZbc5tRVw1/4P6jmzOwBSEe2WzJB5HeRL6IJHanYc5W8shaIuRWHTpxin8rkNxL+Z5x8enbZ2O
JfV2N3bECahOds/vwkVt6xMrNHJiaIl7mexssIjgth21kJqJD8GQYZjmi5SL62zgIuSXjpCsiB1f
CqtJ6pt4KBb/m1ssLYpliSd8Lrd/hkjlYAWW3BjOrOHDAe2phiDL2biA9rhwO9F5cyeHoqeQ6ufY
HFd8yCD2ckl6FOAQvXi65s+qWoBPS9eZWcbHQK4tnO4nNC4kGwO3UWI9NYqANGkVW+KFn4gjyZkU
ph1Hi6jq/zITrO7I/RvqACNLVRzxYV/kVE+SBKI7bCQLDlVOSJRMWvi6a1tEer4OSOuFDlDkojnr
ll01RCBiDWhRopy+fYvaTV3AmUQHcL1/Hs48lJ0Vs8vRsnUG4P54dG4q/ywk0sTNXVqLjCitxWQ3
+P/Kf96xwVh1Kk/3HQTTn3BQULEnuXY69+MXjdV3v5hYYdj2O/UIfAmNCTgdeP9kdzegMNAxIyzf
9BtdBMAo01XnciW2L86tPeWImBHrMdqNoS5z2LXy17XhzSawN7EbAK96SVlA5yvS6ihl7CsXA6fH
hpSGI0IQF+2lt0yGtSrDztMXZvDJwQ9JNaLyTtjRWqX83OIwqoQPRIX+LiyKJL8GMU0jc56CzIvF
hyTGN6IcAI712nYqs2ceWuR/fH4Z0I9IYUrl9tpTd6SvEGkPk3q8Z9WlvBFMzyZ/5NAjL1Eb4jwL
yMmurLS7x18+G+jd9eMNowYIMsUqzYdU14lxLKBwvLCGJ1yO50bouvWCvHTBcNa92zFoxpY08QC+
KZ4+a7ITGD7pJoJGmouoC0AddCPt9qnQasp4Y/e57A9qWL0Egl2szi2Zuoh1QMqOM74EfNFd44yS
B898Ctf5GbTgxjHA7sJc2JtfcMTUpdZwCk+lecMhmLrtFkmNFHDzObgUEDloHfU3Rm7Lqt7nXKrV
Rj/1fqpb03B0jaTfoPbrbMC4ZS68BXjnMc+xUVrGBDLN2+QQIe96IQ8/9u/IDeRSy/4q3vhuxWFu
n9axPc5N8OstaizCev7G2eoB3vyInFmbptF/sMbwkK6Ef/eQp52EUQ4xeoejpIlPBYBQzRIWVzzD
MfwKOCg5qaWR+4SDF5WLEZ/lMzfEkx67EFcO/plBW4PLkl4K1SJ3jRCM+OfxMsqd7HvNmBE+p7Xt
jJmXGKyoZCSD7HUGwR9Ptz8fSnLa3V/dyWP+PikDIR98BYnC+KUktH3OZPubska4GRZWDUAHn7On
d/y6ETNQiuTaFkMzET5K9WVNKz6L1N7aWkZOHnnCmU80o11J3ZOUvamr9WkJRvJXHNWmrnxyL2v5
UtqvsaXjnTVk4zoAAkB7aXxGwwYpXfSz7WEWiQoE9+3d+cksAI/+6YhQ+ORuHCpDcZ49y97Ig1Ka
Ld00le7v539ctWkitUevxGgP3hUk4BaSz42TUVVeV7odTYf5NWt83i9nuNzo97rrY9OOtBqvCEsR
1ykp0wtDqCtwS9UdQUjCRKkzBqh0gmXg/442/GbGVRROMSObaZD+lPnAobOOTXpM8h1ipAky3uZl
JJe/xN0wJzsVNbTFG+gJzWLj+l3yOuKXpYi6tunhmAHExL18fDTg1Y4myCT/lKhf55hhsc/Jb55u
FUUwHzLf8C//kFrMf539T00bBN89UAgrZTB1rGpo/bYgqCWilxH6x0ACPskz8LhbBUu982I2ds+B
w+9BDopOp4IZJ1Bclfem8/3ovdnVMeVMeiH+9K6BmU0SRjn7B9ui/dkctg8+3MbV+eFq+Xg4daDW
SVRFSUOXuovVt+NpNSTEUQxqBKUUSrFen9HyZAJQpYXZ7CuRWH6m7nSFdptpcv38QB9dMSGfHUMC
DjfjkGMRSrvDlJY6NRRTHUWjw9X/S9a9GW36oYtakuQh44eiB5GBVkUAgel0GpX7fAMrheffH2xq
u0pTtLsGzDJJW1NX6UOYL5YzPG3xTNyUZjRKfPrChBVCVFT9FnHYMjMI+xdky0fkfAyvkriY2un5
e9VAkVYy5pYkEAzxGZLkhKQo8UEmCay7tOSS8+3urxU5ueFUyt53RRa6xrBn0xCIjqC+YlvJMcO0
EdRkEcCXLn4PZSJIZv6j6RU/HdYjVNPn2n0Zl6ogYevyd225ccJXkhjt13m++qgfd77JulgoY+wb
2XGmXjSq3BlyFqT6r8tqXRwfeTLEezInoqOhDXHV8iobbjECHpZ/rkaxj1eyrY95O+Jo/I20K6H9
EC320GrhcRWBRqU4y8GHE8SQ+VBIlAoCEuSb7yb0/63vScQHtHA7WUFDE0b8omaOLdtQqd3b0wjW
Lk9F1WR1DvAAujOBMduoAWAyYxnj9/SacREwPhk78qHqNbzvxTEVT5SxIWzrri8Nwo9qBgiPhFYm
Opy5TjTHqGPym5U0HhmDk38hp6iWltfHZ9VkgR3/gNozp/L3tbtEHApnh71yPmccrEri08Exc8oE
95edXmMWAtkSmqfDRkVPmVoc3Muf82k5BNpzE1ThXzkI4qpS10RhgdXITRiKNIAnb79IKLgtVm7h
3ibbtA4E0TmowXJpCnU/K5EoBe3NTz1MswdZiYtL+uUP5mP5ipvSBlgef+ky5NeXAJ07Eb6IPfLg
Lgnbl42+lSaGahny9cNRHLtYSTjh3ve/y9T0ilMGCZWLN3Em+QUcrWcW78k7VcL5/u0/GZRRG8Kk
4XM/V7ioXccDqDzw60ODDguDHHwKbHGQQl5cyNtOSzCvc5vLoF6iUsGbROy+Y4K4lcNHf4O/GJDq
Fh86qMRgOQIrr4U7d6fgm3mtXQQlxKoUdK5yx5zBHWo6ZTqHZXwykEO5mIvYqNNm0Sz44s0S11KN
dMxsXcW6MICZcmtQiswq2KIPdXSC/ocgIhUy6qRLyfHZvzUjluLRZvxqhplQVaqbnOci1qm08pZr
BY0xEmFsC7lvXmqDpZyxo+hosC7VU6f1ruBb79IR+VMbj6qBgpE9UIc8vzZ06X7HrmkyKgMqns3G
u/6bS9+WQqE45+5Aqo2as1TpSbI3YZvybLGkYym3GwgNKs/kkUMixfnMYLJcGfh2bxRj5sOrSCpg
YZyveAhc9XS8Rp31Xn9Q//WBugc3KsIJHgIMKEKWobkgOweNWJdoKyE/z8H2ChrJasOl2xedY893
lIOvTJF+DCJrptkMhXJ9JqSe760GyILwThwATn1v5aL0MSIX9I7C/K1mJirbLvlyHXCcerii0cZN
amkAbcJ6cScvM92ePFL8adrryEJ7TGhRhBsmbMv5es0act6MmiWBmnfwnzXFu3Qmcs9xJOre5WWy
Hj6Ym2qSHmTt+9VuRSFEDaRrZXtt6SL9URHTJtXQaACLvhVzWm+fMRTjteoeG0sFpvzBhKraZDQF
0aKGPT1f4NfcQ82DQd3EnhvtiUebSLQKyQZenzhsAKjkq2crbpHWZN21SIsoWi9EWFV2JxMGJrDC
WB6ULUR40vYNJjXb+L6qp4EpCZeRm24t+lVHEvi8uE2CJRqF8P7mV9375hrGZZY+Hd9qZwQZQoyH
WJEd6KVhYAr6IJgtGP9cQ7q1EVEVv8+iVdDMAyLcx4UgoJqnfDlhdySgZdfpYj54iN4KnWDDGS5X
VN1qK/dCu2wNlzU+75Ztec42h9gvSD9GEdVGv+GAGz4pJ8D5wP4tSrqoOpZj9uZ1PikUF6HsExYJ
UC6vaj8AQ1/0NxA54jEga39IMY6y2dliTCyyJkf4/xEphiXCblb9BkzV0HeyskxQu2scg8gwtdLL
ASP/0fVzPSUi5SqvWL9wamh8zj3QVIv/UTvPAIg+2WUk6Ry0wjWf0/milFQuYREo1NwNQjA/JIhW
mClJKh1f96hXYC9pWAgPdUrdxxkc/WHH9CcD5mWYUsghI9MKNaYJMpl+u6VewamAnhUsioBcCvtP
wrH02uEi6RBGJnkniBnVEI+3S3ovUlESIvwpdRm7dERCP8qMhCCjVHzBLFQ6HW2FSg8YtF0FV7Om
URpc9CzRtdTBoVudQ9GsyVrv2YeWElrtxm9XxkC/xnL9g6vU4PO3telXGOY17TdjlDwXO+WshSBa
esmUYO8DYYF8ykbyqDyNEj3FI3NFgUeBRU7H66HM+7HZYXDPus4g8BUuAtU164paiXnpYDkPeboI
Gldsw+gxhikakCvmzwMJTmiNdy4xLukN8BAJzQBKYA1piXoOIVQEzC42OEDLIRO3I+rb0PceQ1j5
xgOQHQSHZ6443Efk+0Hj9deP4vRMJ+D1EJRBNBYKxLe5Lt9YuLf23e1jDBvh8UUlgKzNF9eXU1XD
T8vJE+mOXI2PK58tH2NspgIABAYnrL0RRc7+xyAE2WlucNrXu1Tu95I7ufIhR0LtdJhnJfQZO0Dh
TE6cwxDAiZwhRDO1o9/FGV7qV7w3ZzU+vW9z4Njp+i94GahMT10N4t77oOnPZUANJvpgyrK5kd2w
kBQ4cL9+ZIWyhID0h6RUYdDbupn6qJ6b1TWrRoyxwibsyM9+WdE+W43hhsf4NCfYjFzYsSfSyB+s
H+VAKrmoa+M1K2n6QvGFgwDX1L7kGiCfiTeM10yHcQW4zCZ/8gOTkAi7enWkBTxHf9iG0e/8ACgy
2NLbZjSXue+mgEp6L0OHJvuraQGPIg6Nb+jUvGkJh3kl0JNtIKsWIYrymJZV3AOLDkqq2s/X0Ntm
L53LPPv/Q3zM1XyDcaWtWT6lvFmPFP6YWhTG2vLVBNuGE4Z1QAJRjOC99NKJ3bWoIO9tvmnppXEv
kEx4qt37z2DB7KyRkLl63k3y/pV5FzJH02GUrbzCw//uKS4WqAOUZpOpd8D9lY9i/xiRxvpSCvxh
+958WoITxU7Zh1DpE3/vTysUkY5OC7kMjW3h+TK9AZkh/THIYqGRonhlH93+iSbMJxjyayDJ40oL
eEROoVFCKeHSVsVW1OPka0tRJFca0KYi3N5LVZ+sziQaT7FKDEe33HFoUyH9OXW6bpx8rxJy54X6
f85f963tSA2dzc1P2g2BD1SZn2GlP6ka0no9RNaFSTA4vuiyR8meSdcVJ0bSM43Enq9tH/GaS0Br
qdPbx4gFieXcKIviS+59cSarGqRanj3cPyoJKBQWi1Hs2jfUWxJVL9oWKbIgdZ8Tu/JoCDF/gFtp
/83gZ3hqQaXf4bHE1/sYDTfd6z4FFgSyWsH37L+qiaWXRg1GkGFdOafcWocwF9Cso22m6bBGk+xX
EMPH2fvVK/pfMUWgWcwtOIfweuqS99lMe6N64zsHVYHbJO0TIb8ziAtsQdpJ2VwBI/qsh22MvaQc
Oo2UWiRgtPjHhI5pr8blSGe2tFe9ucL3feJ90QO+2v6b2Dat+zSMeqwKfXJo50AoYJiO1wyo7X19
II5emjBrnyCbveqapvU/Rv7N8w9Q0t4LqTa4qs93BmntSmSK7qNdXUF4na4XbDYrZfMsr9QfvXJV
gZEyGvNlggj9NwYGL62x+OyiTaE+k5hkN6AhFptgEXdsd3yJifIGW1VFwEoNi/3nTK3KVAtpfRxc
Xx6K0LxWAnGws4CSutbX7IsLTlaPE7wYQMoO3s3kB+NjGO7D+83wry0a5f5vwQPQEs7kSop7HqzD
FxrY18diRm1T7Uh/s1o0ZyK0Ppu7GUgLBADKyQ+DlpgiU8q3++PKFhOdYoh8V7KOi3t47TuHhdWK
ZsNQ5IBJIhevC27Nj8vsit92/p/YC6z5Dxks/ZAYGXk86jwBU5MJagEPZ7Ob4mnfIedhGQIbBYkJ
Ivu8WoaYtA9zYPObX0bhXBb8qhqsG2Uwz71jiWFZecFFp4KTD6AW7N1ulOAtEmEPV4/9S8z/ykcH
i4VUQFvJj/0QrJGgOZen7/FmyzUEndyNfcyoGUp7LNWJGm2OgJ23mlUK15cuXwwMDqrtFmFCZflv
XFmeS3+M+blPDp/6kjL4a828kUd+UAgZZK76vLqygjwrtNbCmjBilnkCXlk3b4e0FarPOKcwoOcz
2LGukDyt+IbTjC5cXvkhtY7/wvbWvdyZrlq4bh3lK1e2llLUZTZAEpVKpeINDfCPOXz6P8i+U21p
XoSDgZqzCb7mnGFObBTS/1JKAZ4WPiILiRlZTDVM++fwEOSQUgeVDJ/z6x1+OVRkk9wqq5wBQVRT
GlMMHLN3OOseyT/b2znYJn5dx4hLSD/WhPgWnN9mst4SP+qWQt8bPnvsIKqkJtyL3AWX1NqBVca5
zBbUuNjDrTBSqlXmZcY563XhVyHFSzyjoS8xOX/7lS1V9UEsH7DXx7ggWXR6DuX9Wte/3Ncl8mIm
1oNBZ3wXiHkJWoZmud90rXa72FZ4KnVh+tPtPe8L40P0qjpoPMtGh3h8OEg4iZGG5lReNHUeKKir
gAlnoXwB/rpf0S7KoJF/eWQZfZTXJs9ggErgMrgFdBUqiSIEajqgV7NMTEHqZhcSCHGysmmbnqfs
nfWc6hEACmIVBjbImF2W27Qirqzwj+vIWCOist17oLt9Kf2MkbJ4uV7JgU2RUcOQHWp3BWHHPrj6
HO8PE7fXSY/CIa+jya0lv66P0EcqLcwoJzSHoxzUcQq/fo7KPxhDufLyzHQxaXw0boibggez4hIR
e/LeGnZkRFyeP7NO/UrA1WeTbu0khqDD3Q+wUUaIZixZPLl/SRum1W6K/aRuUn9c+cViQb1SdzoX
LJjxXCrU+IM0Gl1fXH6Ftzvn+eCsYyexFsxD3C55oysywppIjPq/jnY99Dn8ekDPvCZ9JmirtQJB
62029jdWNKxFPDaV9G6u4YD6FUcTVPbx2+VC+asqBkkolZeU/IHisWHzsVryq5JgDgE4KLYXdnYo
SSsCu4Y/BNmJFseXITx5AEm/vak10KxCGN1kmwHUqmTw7bWF+aNIP6ZxS46lFlY+3AXzoKjRQ4gu
+pE+w8xwAoDC3Ma1HlzSlc2WqdrOm1z3eBlNTXbTrpjPSgSQUJvSqgaCSQ/CavmLa8zGglzna9tg
Tvn0OcOzGMQcpaxr/5gPoGxEqLthng8ccmmv6mVCuH0cPgfYRpTLnpdLNYLm8fKchWoPnopqZfRG
fsBjaK8J3hyyiKWEyWYzobRqXvO7JcEe5oaXDZCWoEBwbzXhXeBnei6O60o7su6yDGgbxwa75EXS
wLrvka3gH+lBlDOU8xXlzqKDpVAnTFbX5sOWiS96HdXrn/6KpKsQNQqlqM5Wbq7DNKQKZnCnWmQR
VHzO/FqN8g5SxHvBKz3OzNrd5uv8BKSRMW5jJMMikM/BEOCN+BF/yuHvVjLxfkg9y40zG3X5BlLn
7YEhIBDpV4RKxv+orVT8pZx9wUdenSKOyFUPJ4o6j1epGeQbi6gIwjuG79nFKCfXmSlx0vEk5ybR
JGiCecZPsZtApnQfunj66ClJOc99PE+e9vBrHKh6EeGJOT1jCpqfJ2Adw2n1/5jtqPGkk3JdbQcL
y4B90PNeBt1WO5sBORZXbjMagpyY5ztwV2p2sUwlTCSzbf0ZAHVzxCKpbY+7MtsCeZ5qTFxtUJ+U
Z6/9jXyYLiroGNgMIIV4wjeRDo426aVtTzRGnZfi3xT4WMrFUAyWtCX3bOS6PbKtAaLp82oM8lZq
RtbgkYSkH+QXjUBbSrbVm52EI7iAk2nzMqUBGjzA7gvFORqX2qZ9gVBL07d/uc9dlz6aFfie4sq+
InRgK1tRZvNmvhYz2dVRyLweC6OTnEqRdQNtfPCd/BwQTrNHRu1vndIdS3uKXlm1F03/O21XRzxL
0kJtitpnzLXhHBWejigaM74yNzf4ALyuuR7oMvkM1d6gvbGKL6MWPKaeROXR9w4smYG/LVM/+xNr
TTRLDbCHBYh4S3PGNSA4cIQ16RBWay1ShjjETVBmVGUqIiq6Sv+dnU9C44JWdOzTkQ1W14W6Flro
Bqc8XbagOCOAorGvLFxQWMnNs27oMnhZX55sZTL3WPat0lHCo6BMxA6X2BS6A/kS8KHxyesmfhN+
3UPkHByF9CjLq7/ov49t76qcvZDmsy/YydfvBDJKXYKO0Z9r7artcs58gNsAX/hXRN4iDizMxU6i
kPAmMLhMJeWnhqYhFq3YVd0/hXbJ7qx15V6tMO7Ft87+8IXYcdcSxcFfeWVG7Zbu+ynuHVv97M3C
Q+QXCIvZ4GMSpKC+zdibPRdHr7zwcWmB56AvXu0OTlvmzQHprzCa3d/+5vD1EFv23FYEKVKaMHwR
FetoxqGY6CeoY4ImJY4c+0BtzugNjrsj8cp44wGvjXSYEHC99MbK691NrZS3Oph3SOpmpg3kgeDi
V/g8+UJ9s2BdG5nlPOiDsRa2gZqMbCn6SMAsgzlYznYCO85IxP3CHDLMPL/1sdsm+GdNg3oRsLP0
GnZemJhg5llZCHdmE/5jtmlW89RejTU7UUWRpNW/zC7TguKOM5UpOuiNhj7fyC+60W4nWBxWmmCE
mBRA/hz6ejvOmHSjcdbZuo+y1MDfyTym5v7LfxTGkEFCkVfI/2TN4+ihUFRlfhmra1GFvgi8mmcp
HLkdWEqJGh5attXWdUzyl2J6GE2l95Dp4ZgYO2POqfoh7NKjjVON/c//5Dk3PBALx+tL7e1ydHNU
xpKRVzHUmFzxPvx9Z49d+RL0Nmz0st1S3iICfbUX/SEPt8/xB40SPEs5sJOZzZkWiLj2fWgT9F9a
Mp/qP4ihhk/2PLmGbUkYgV13UQkE447AqupNQe2ocZXBGq7aSOKf12xWW1HYWDyxm3IKapEHlhOg
gX4BiLoXnH/Pow0QxECqE7YCyFuFkWNY/msE8MwHCQttCMIvkPLX79zu6PUrXZWdSYsHrC/hYLKy
qMg0cNPMLx+OrBApP8CBKSK0lO4yoSCKdXfEtL7jGARikBwQWJnIp2a2eHel7GxwtPL2UBPTjbNg
Uq6WdJ7nVin1Shgd84BYzj1tRbipKEqJ2xHoPmulAAcTZn5SqlVRVt6OZ0D9orWVFk6/3EGJwWT1
LG0TMz1I9HXyNoeJKH9ypG64fL2rlk8YYsrxuUB8GyDBXU3Lp/2gMv65jFdhK9r8HSLNRH9ZDyq0
tukAsxPDLLQJ4Wclg+tSgAFt+eUd+ITKO3j7aHG/25dmdecKqwGap+EbClL+FbWQ8lxPsV3uzP23
vqGLWqtu6E5XcMCR2r9UcZncIpvZX/Z5/IqK3V4ND6IdzJP6tia26VCcDgSv+UiUqFPgHPp/sePM
xTZzJcuXwCHn4PFQssQlV6oFOs/s10pZpfwYeL1IJBTJxqxrEoB/CGUgAwHX+OS0C6Tw2bLg1on1
lr6yRQQ+B8GXUvyT2+Egcx+1C4kXseH+7VkbR5NHc21lPHHNNtcP5kxFokkhyJOndCwEdd6q52eG
fNviIYDsxb1/RN4+RH37IOA4gC6xqEH3Lh8dnEWaP3N+2ZoYJ+4FNviA/bN75ltBOiNsA4XBvmrF
8M1id/j1ECtlcgb1mGee7p8nBg7793jk13vINWO3q5wx+WLdpm7C8xJm5Yz3cZGPzl7m0QYtEa3I
BnNyfrHysQsEkKafhUQ8ogWK4+1PE657iyfLZh/plvefXehxZMtAZb+yhJPBJrVhRND7vNCVtbWp
/lKyuG+WF0XaR3PJ/GQj3zMaLlq67XaziLl6v8Kn3sREZwuYA2fDADeM4ONxG7myHNyL5FsWF+8V
n8VG4H/6kLoC35z7S/LExacytrlAL4c3UD30UA4wbMd0VdGYoEE5QLj+03iJ1dDkcYIvXEiJPejY
aiIxLODUjRLvrqYVLG/3w8dGmZI9cPgDMWEfw6U/9c5Zz3FHfeqV18n9O3WFSuu7BzSxKXszdPIs
W2J9RYORwhuCMQY4eVXIQD8d/8L+zLB5d2jZkzMKJ/J2nK5gGPLdH2cGSpWd9ACSd6bxS7lJCXKO
kXzu/b0p7To5iKqmX0UDMFVRI6CpcKpZKYhRfk3vli5c2Ipu11yuCwAOujlVpuQ3DkQptj3/2l9O
TUMZoE/N4yWqjZnBPuIyFM2kfhNy1SKbBPNNjG7WAk7d7igRA/M8WN5jFH/8YTs669WQObJI41b7
H6P0+rD4KobPovD487UZk3s051EYZ7TO+nmbKGHd4rRlrKhLJlC3KqahbfhFYLtSHMOAFqvSxUXj
11Q/OzjdmxLdfBlDmh9lUkardbMDn+x2lcZ/PN4rlMQ2fan06FOD24CkQEgEkfJq/zviRJy8ieR0
vlspyXtqMt4RoAEHGg5eVMBGoW17M/ico/iQd4m9DFzXJahwfjp6cmXKBbipTFG7fmj+XJbrIv7T
G57dfu5CYlhItqNnPJ6E21lsYyO3xa1KFEaMh56+yjkP6vLmfm3jHiD8lhiz7uwgUdpYWtG0XB9P
7a7Z6SgP2cBAFQm42O59NcX386omuMI2wylWF2SHbxzchyX3GcN4iVm3rORHbHpBG7KFQylWUe0K
aHyJrexQ2IjKVj5rOXul0qbw7QZ4YvvD/b6a5gt+VNCdhrrMbVorSbZjQXP9Hjv85+tSnQHfv3NH
0IO+qli+yMAIiLjlT65vFPL2qLIjCEMOScWbcUGcMwTEJCi/Xk+fSYAVRjC7f1s+/bjbdK0faQxS
LY5Ga6LR8uZ6UukjqZBiN6cg2aQYuYo9fGISQ2ePQU6Wzcs6QN+D4hzDjOqWIAhphk15XMIMuxTb
EVD6+qd929g85TFgWr+RRvWrDpHHrm1AC+W+UDhlVNgQqmkjakAqfjkV8gRGtYSOlxf4j/6acFjs
HDZAswIj9TP0wNFpa+VMX1vJB2EaDiV8JQqaJagQ3SsbPc5qrfHmdK2f6Fyrbps88FvKB89XTHUr
vdQEogxBN/AEotUsFt7Df2oDDHIwQ2TdLNN7yH9ag7zsZYvO1I/RhEVNIueHd3jTylxdNwxohLg4
/kmokW4BL7jhFgQy2x9YAt7H5/4nppPZB0CCubSO7PWf3BBjMAga9dzt2+RkO/oAAMzBROr0T8Fg
pZaa3aIioyl1WfXGZ/DoIW7SxRczAZ5BFkqTngtu76ZM5Qs+i1IxB8oWwx8z05g4nBCVCWcfdQh6
B28wtgszPiF22Wb147nAHVOzQevoZ4YzerdfNWDhCX0oN0ZzwuL2V4dJdcXm9Dvzi8x0Foi5hUwb
lVBOEc45V5PDN99hNYNX/ZcX4CL/s0bEcOScPDyZvP3X7IpRIxWw3TynBh8gIEWtjRsNBFm/k+zd
4Vm9ElTT4kvyrkgC6F/NkPaJNmVBKNzYexur/fauxPnqVIu7KpstKtM3nkr1ztjJ6gd3BbJ7HLkt
cR0fFp1LEdAVYYm03JZANhVLxk3R+tTnFc7zwl+eiIS2M8jH7jKja2orGh14D1oBVUn1r4ja66/C
rQ3j7PdP82zU2O9f2CSli+03+MePkAJ9BO8M2S6c0zADPqJy06kYsD1HywcZ6Dq49mp363pb6OBu
DA4/LAmvz3nvQRkNPjlwi5JM013UHDdLuao6UVhC6puxFqorG0XGH03hw9XphbiybeVowdoTRD2Y
Yooj9BbhoHWhtbLinwNm/73ODu3+pROiSUg6FTyclJyfCIjarHH8jchgeUdgqNh1hZT+Aum9Euyi
+BDhJQq44/ujfoH0Pb/X7PiS/vVdlhHKTdFLeaukmUSJbGTmQhNjI8wkyvZKLcLwRY4aB1h17eJK
M0v9UsHzvyUUT6nCu8ksEiRWWF14v7Xa4GekGaA96cdGjBTMcpX7eokNdEHkiSGzBRzxyJOQzhpn
9wMDo9gTUZDM6+HoJQMUceA4SxqwZd0fD55CfcoKIk530Ix6zOmuBfdFii0SUR5YtpZ8v7ekzZYv
OyBE3p0JSbhSjN7hzmtZhAMh6Dkwl4B/FyPBZRK2deBSsnFcIE9VHodnVq88inIepPKVi8QfLu7u
6O1FCq0lzZHwQCpKXTzrTXgUIsCRnOvuc2HmlNYEGmhqwnJqHnKXCpooAAJfjf4NnK79TAXJdhdp
OjLZ7rxbFWypoZ5021AMlMwLyzxf9lE/gzcp4/SIy3lHwyAhDcIUhWFEVNHh/wc+9iSGlwXFIX6X
+kAnXurd4zmqp5GVn6C8B3XiPDTc7BWPXXCjXZkfHfq6wDWMm9B4WwRwpAo+FDWNVehqHhldWCcn
9mNnKbvZ41Nsr8RweizZxD5sIkNPZb3qqORwOFp4RPwmvroc7PmZsh7yJEtQ2iMxWbRPn7PkjUq4
IOaBW/D28/pJQrI8VWPJQrp+TnQWIWU5jrycx5zyy+ocynvRER+XUv7puMbYFy3EKWBmDZL0Q0yV
f2h2regHeVvuEWtL+9v5qbKjjeenVnDlk0+JTNqEdnqpDQuRBI0PTJzUUyXTeRELOYUi24EpqiF4
9bOzGJHs0stCm9Bo1Y6oGcP/C75AhZ8gZL2Esll8oBQ6rvTUIjlS3S0S8yfGwHmw78cY1WyNRp0H
c2nRVxqZsVlXMmvatiXfMy1LDcgj8FBRseC8ieq7WuRpzmgVDPLXpUJBvj1M3H7j8LkAAK/IVgW/
RQgU6zJaRVnBVJ/fp9CU3NdNxAgv7EN4pyAwOxZIy8P1z3CkKKnlqxBdtREzN3l/R5zW/ZrIIU6Y
2RiNxy2kAURHkgFG5kcAJhG0DB4qw14xRyaZfiAsrQV9tkjY6ueiLekqJi5stmh5BDOA/IPlGh5g
GTlU1yUzObDdO644ShvKxdHVgJfQ23WlZkwg3cJioo538DHqtuX6/CzlUkIOB+EtEaoXaMXeyP95
KGaYEjpjBTuoBSgBNy9sIJlwtuT1//0dgQhGtHnDCISH4XlO8HUm02fYatJOdblxrqJOVgB3oUgc
BNNazNXckFGdZfMm+6jUWPeCYJkBr1VcfFsQlNAwkikdvJwThN+mQezLPQpUJzfMxO46eFHLz6Gi
gWDsOZj1Qfy6VmxEP7aEa9j70Yguj8GmNkebIiWM7kEXPTrNG8dKh2QwWR0ewh/twNVuHgtF9Mnh
gQmsvcTufbKf5JYeDKPGz/GzCGXXIPN1BGO4VftQfjh5PwG662ZXYiAoGfYZ17wPp1cYbeRdFiBG
7nJzRNuxZYnyzoe3PKNwD1XraKejtuYd9/1CTKFhZxu4qjy1FNzkYMpjFH5gzi0zdLYNyEODTKeJ
aEyIfd8rmuUATiUBICSGU6USVZinZqF4PKzRahDArxRpfzUHbMAJrwJIO+DFdtjfn3UWC8e/sjKs
StrRG3ax2pNBq0Wz260ZUH2TjC6oKNaozQtwhSB8ucga7JopncKfWa03jv6ug18xf48HpKnJTk6L
7X+btKyy0d6u+5OCUWsNdUDAet7VTLIaZlJimaR3VVcgFRKCVF5zDQmqV43iCPhITUc3HAlM8d8X
6Qxq+oOSUIaAvHqHsw/QoP7sM1J/DjQP7DXWz7BAaedh2JZQttKCIYPVqGy2Gkje9LmqhMpEZnJM
kVO7FRZnejkPLJyTQuzfgndqeQ68TT1wxSpmUSgsLXIRvu/VNPkG204o9iLvcvMMG5wb7L4Awlqz
LupTu4sEzXKZ0oCGfGzV3bWHkyQWszJhS7lvpQ4bSifdx2sSDopfZAAz6O5r0HJpyMqLiEYryzGi
CQfvAJDRnRUkPQlKe8ssglp5w8YV25AwdF88QzRXZj0mjNsx6/74mk9JCoKRGQlx1Vux7Mc+vVKb
HioAR1f1JOngklRlxye5mElMTW8UaUdEpwD2jk9Dwa4lekFJB2YYEMuCDEoxHYOVAeGSzE0HBfA8
ZPISJM3MjVtHPZhWj/aKDTrNttWoPEM1nLCWQ4gsS/HG85uz5sb/PewhWmfsu7KJab2qjwhUa9V7
vMtUUngCOXk/ol3dGlE8AJPoJNMZsBc2hrTyDyu9Pk/7ed/zHLfqojug+zD0nn1i6oWIsOFEmkKV
IVtx9HaB/ogx4bs0hK8T+alUywD1vrGXmmAxNQSSpM3UNEWMWofZ+lmoVB2e426nU0CubK58pvn2
RgMYmyIdxr/ZFDKzIq9lOPSbtDD8XlNi21Cmz+bxBPgLKJoF4biz0jNU37ca67eXRWRPl6FPYJ8b
XrJ6is1wY8QoGTumDWQf6InGo284iovF2fZfuBTrU8CjDorJhpRtNui/BJZoVoh2hEA+oISvVv8+
FXjbcDKQgQtrIdT3j8PM9NyR2taZ1ZgJdPwsX6HDifVRG+JfP8W2et7DTPYZVetvDAZVXLZCZth/
oTuwoStCYnmaboZ3KfVfN1LEoMKhnEu1H6fZkrmWEpdHbC9oXd++0YhEMB8LH1pKcKAIpzngH3R6
ZFY3cfU9dhKG7JQwPwolcGC0Em9u28R+VpA5rN0t7c+Sfv9ciLRV5mBEdDYg8t7Y7eVg5Mvqn+LQ
kO+5a9k0syAJ0Tz4lEpD+WE6IjRW/8/mpuIOBrAYmpj+3htrmapdhpHm9t9QMsEgxIXlCo3wxNio
ucMq5YFNCI3qyN+nhP1jddrYRSwYYo6v2+biYfLKzRp0T9t8pD1lMT0jFdYlM6e4kDZqF/asaBdW
cY4pRMbstaoWjpxcBbWtzaxV5aSVFY85NSaSteHy+G9zGG/RajEKwyJfxkcay8QS5DPlVFQra5Zt
erEru/NwV0rW6e2APTEb4kokLmKkhgDDFmG2ZOF66t5gwKoG9Q535UiGFKVXYrO9/zH06VAoPRrt
gxtlMfljzQErQa5VZDK4N3dWKvV53TvBR2XZKqXFQEqSVqXOguT8fAYwjSxfZFfeOiV2cAZdE+x/
SCbXep1eb9Rz4hfhP5fyA9u3m/tuDT6SV3pbFqyb19a5xQdDpT5GfOos3wwCG48H9pCcdwKXY1Oa
nw2ZnghLO7EhkKvo00NwfW9Gpui9FjZ0UTLIdhLNpXAanoON+X7bGW/WDd617IJypz0GYL6HV+E2
McFtL1tX/ZEv5wiNgURzh20O96myu0tNedVUlCBwyTmKkWZC9yKvI4Z61QAwHeamxh6R51c8pTmv
QYA145whaJtvChx0OQW5CrB0ldQLvoPC473XNMrwa3rC/kq+nlRq3fE8nXE36dah1h2oFaCdIN2l
FpFczaYiaY0blMuzlEiARZaigsGAOh4+R+qTVfb2SXIBFeNSjtOzSWR3RC4Z0oNzr/UH2bobl9pq
yyWryl5o36X2g5oTI0gyXRIKpQYTX46eXG8N7QxmFYorIQ2AsgvkgXu2cVtbvUyKw0RZxmC4iVJH
OE3pjRf8JP7jgJ7dQ/tk77TZ6GCAbhaP3vbiB4aH5UCRS9ZTHsQqnehv0n6fjOYLAf3IUkn6QtXI
AS+s9PvAphJikqedrbVmLBAQzCNeIaUKryNVzOMd3x8rPP8GSNhQEgQqkoGBg7lry94J9JUZSxmp
ySt0LmeBe9tx7nEQJHlgklWCgnfiZXn4AEH1IaWNm3ou10Z9IZkL6X82cXsRpK9zNvNrd1+0MX2t
f1+dRBo1/rWLCVZ0lnjs11NQ1wo7ef1vPgyM2jTTYgNv3zVqBZQuQYqsMvGh0cFOK/gkbQDcdCZb
Q0az5haarMtTuBAPvb+PT5neMKgImjvXs3Lm4W4zp4jeqgkGYNiZ2nD6G7zP1OX+YEXgykS2vLqh
JEGWfJahK75YaqXoct1z1q/B25EB+xhp9CdxRRt3TUpdyq1RYIv3Y9fU6zHYG3LLq3uerHm6Xv8y
D7j4/1lnndjY2pCnHaumEXrUAU73+pqdITSXxLPbWEARpOciQiMZSm1Awab9Ox3hLCMqJHYUyfYQ
FWLx8NL+AA5XguhAG8saRGPsszgT987/rjykna/MktplyphMudOUnfNTcx7lXy5+3E4ubOwhd504
FnSWSDdoMzm7BXuCxLvb+5iA7kwnVoOWVuOYiBXZGitUJRj2MiNPed94KQXGzVBhUdk42r03jgC4
8o7+jVpERBwVOHdlkoMrL9dN5o0aVkRnFbMMy6C00H0nmC8YCw8Oa4/bl7WxGe4Cwz/r0/NATd9m
wpKb4NrL0lUWyNHqS6z/iXXP8iT4ZvkYh7ckpfYRWndAbymtIna1disetTFBov3wIQhtoXmwtDKl
/fhgLRb4aUtfcSGfUIpbiQCRQrUR0ZSz5iNkVHclF55/1/YNkFPzpMQep9vgbzRHkFJ4ePMbkOXe
5vX3rOen/c4RaatubjbAOFVqk7Qx9wIWqEU3lUus/p3zoBWN68UmsEMrnJF/rbBQEsETl0hcNoBC
bf0Hjfmb+GSGa869GdcI9kOEZEgqzAvlcI76a88xetyOkq9Vg9J0JVN3y836zv/4K6+xgp6z9sx9
/1jhLIS0FYUIH2yPu+MWNu72wDvd0rFOKoNEpQ/WJOeSb8M+IZ0Bg0nRnsWiy0dVYUUD81U2XvGU
WJ1zjnKgMzbJW12XdVa+TMIXmcPy+dh1CB5O1WTUvoBgAcki6uePSwc9foVcxrUDjXHGRO8GVkfz
xqAlEvt4UOcRZtay70DOWttixo6ZmPX4ZX6vMmye4LLbnhsSkZDIzNXQ+Gd3D2rRPT88dV6cJdBr
Bvn8R/65AmbbbEvrySS/j5IPnku6IyR/8RVdWY64q0xSvPiC5oPTxTfry8F917kkcot1Oh6zaizx
zFvMz7eGcoBxoRjRYcgxCOrpYUeJdCLzcg2McaOfNS/LpE5H+4PvO5REg3CUeA0ObulApDAatzdO
cfGdX7oye3D6Rdee008N3PHgF4I2nmOYpe/30ZslJeGj03kGs/0olXaKKsk3jA40NcHtdpT0aUeq
at9HVf3s1E1sV76jeVUcSh8vhdQL4G5e+TOmIhiVOedX2+qif9XUNR4tVNLsiqPkinaoSUe7Frk0
CMuAfO3095sPSyOoLeNRfpgeTJNFMDApMzZRI53naVOwJLv/dOdxeRkB39V9UpCQCPXVV6JvrVMr
xkw2vxzFydR+1iROEMGFPeAM1eK0HmA8Hne1mfgUvqQi06/QAMZhvqwfT37sykG+civ/FhBwImWY
zuT68QDo0S8YUl6VsEXBvOXPkqLqOJhJshiRZ1zaIci5D0kazzaVwSCxuhZr1rE81sq1UnvihNxe
sC/BPX446elaGcoAT4KQlWoZf2+ZnSzeLz27UKbcWxov+HfPbmJZA6jmVtHVznGGXb4qy81lBiOn
ncYAQJxhQ7r3OrJLBKEGBzAVXjosid4Eq9LlHubBY5yrbAJKFZakUdmHiJc44aemtL/lFvug0bTj
JCV88F5swO8VXzHApA3pmnKq8VYR/XnKyMZJpn7aaAEnJbaNSL5DOZEW4eLlat//G3bNeKJKv5Ap
r/LRBAlox/HY58rKiABcrF6Yyp9OCj4zHNg3mdkDMgNUCNs32J8/tEkBqFI965+cRgCpvXGl1+Op
gt7rpFX4MMDWjdzJtAlEDyHVkPmroJmytXgWyeEhhl9pN0X6ZENY4hLtmcVwfQI4WElpeTI/dZWM
OqJ12Jtq2Kq5TTjTei8BbIxY1tEyHveT/+eixFAzSJUr73JvUT9trnxX4HuTqIqWkRXcqU8aPGoT
3RDESgGumpURzZMNV8ojHpbhGxrDahCtueHVPp8Yl2zpQWLKOAHub0eNQk/QUAUs4x6eCDRjvmVQ
0sMMfxopcgAfDSf1Qx41t8b1MbBlTEAwzGOuLgQrQu/NnAz6jC7tFAAjVlSHVNb8ZKkB0BkvmHyv
3QUOrsyo0ROng9e/Wd3jNai+CpYqGxHILpvwZ+r5hG+CGLchEBsXM8k71MlqsgB6R+tvHrrT7T1a
kGAV1r5kN2AcK55q0273ImxcDCXj10j6n7rJd+oGuvr/Qr/BRPT50uOzlSW9FMhRfhdH2h4VkoFM
Bsjup0++4gNP0pV+ZMoUT84bAwev9Uun1eSd9C/CMVtDeviWPLsMZl/ZcZl5eHpV9UzApjo4sQFy
pqaUEcwhWzkxqYvtug7aIohy6IyNEpYMI4TLUuUkoRk+f/QR7C9APzdD1LN1R4pTJJR9Rj9wM4nI
dHmMObKu4zmas2OSs3WilbXjwqSjI3lDOzy6DdU04jz9NTkfnbWamgi3gp1LRHDNaP4nvotrRcDV
gSDtddU9AUoNyXbxTkmdfkSiCpGwT7HDxOveqAO3b7CJAe6R2+3MqN4jj5TtPpfiRH6qs0GWLFGE
IvO1BGfiQnBFGOHFQF6KZaa3jQa7T7q2LdbsfkMjBouIU5bzfSElOQA7mI6L1DFPcMmuePuiSqS6
FrvTElIk1QqXy8IQ6WZyLivDh7q6Co4kac5jGt8A/qxdZLor9vw1/w/PukAJPeDLBcElhoUlUkVX
p7Glvqi+hMkf7B5NopUNnk3wuUHxYOc6g+36mUJdK1a1R1bKtYEL4Z/GS+mgZnsYW56FlZ5Bp4se
C6+iOfGoh131DeZ5hLrsDtXrkBzAYshVyO9FLbND1U3LYrFadab8pLiM/Swt5vFWwg/Zj/6Q4GXN
WgPtdWbN+P96/TDXauA6jTV6j9vDHc2rCiqyBeW+KOZzZ8hC+XcIhV6GElHTkzAzETtVuJ388BxE
pLFVbb3mqTRcU48OPVZodpA0m2IIVsta0QtowGDu6dRGiRvUOWwlJl28DxHSbzLrB2+sVjpb9/o0
dxEViQ3b0ISrk0IqVobHfaVb/9VrVjk9kp6Ug7zFMJcqv+13m+TgjHl43aSXgKP6oXG0WaUvq5qn
yVt5UUrxAGePSUT0VOqjVHZ8K7AKjPateuOJ9z1HnoTX+pZgPzSWWUhArJjLm+rYSVCGR569Sfqw
CkEJJVKnIqoXJj2MeVSZP84bhT2kLAsXONlETlaSvBZmC9VwKZ3k2R9vKK2n9/rMpp8HaOnYdfEp
2xuvD4cj5KqlZtM6p30WMsXu4/+qA8Q7B75ezRe2JfYaBmBre4rYSHaKuO9BWCRSSlKgcpdqhTl5
356FtWQFGhIKdf18VXYp7O8TaCg+x+GtQcCE9BMT4yC4ESXg1o9A+PU2aEjtnPFIqcx56IFkpAbX
oJbtAg9sEU3bZpb0sSLBmkCIqIpglh1JYy0p6UXw/G4hxfc1fIuinwetxQfQfwga6J85xO7KNlHw
w66vxsSnPuVgcKNbysL8QYYP7zl0+qavEBSUsQDrS7q0z1BsPxmwFhIg0B7aGNL/ySh79zBV6ctM
oBu9etVgiWE9AbndTpa3/hcesoCvhK1Jr9Hqu5GlCLY+pMPCnViecDR4/MoCnDS7KDwNQrd43LUr
QSdnRV357Yofp1i/rmpPOjV/4LiBKXWjUcF1eg6BVdb+roTB3z1/YPlk0YHjqMKH06jvriH4L4vI
tQQj7vpWQITNAhn8JH/gG6FIK+JhiSwAKKlAVmZ2Ul5TuJyTtJ4NU34IEQhag08YAPNkA3amBdtj
PY4NTQppN7Yt9H/2X3iEwwa6qQmbFZv/xeWI6rICpQKDHDUw70CGQJwvmrSl7J50d8D8T5KoPZJY
PfwQ2HelNQGRaXXK33qPwj8P/fEIXz8eH7OUFsidHIRbDXgPVkXhbJwBGffhAGN+Gn72GWn1/z0c
PhgUxFrfdrT1apmOqgPNXBz4qG8PMmXDAzcbKblqMsaDwet8l3vw+8eNf+/mjZxj9YHCdSyww05z
1b/Y7Q2iOcRGYLOkWAy5jke5sYmvq2UihYKhezEHzsHqeCX+ZpnSJr1s1Be0q3H9ZVHuAvvs086j
nbGLMkDit5ijF3BXTaokep8UrXMSHzXBA11+5mHYIbMtxhQ15weLVFLwfXyPeg8bnUjw6YssD91e
n/Z7RPdMXb1NnoHFiuWifEUiplnpMNTyuNpq+wRFGXBcjBE8uDNlqAvfCD3TOFkeMwDJ5rjjrMx/
UvGKZLklXA6CXk8GakOGZmP5Ez5LOGxG0upasbrT305TNzqzK7UQl1yc29pTHslB12si1+b92x2V
Ehsxohf1x4HOQ9TdVUS5rf54Hd+uES7r+hOLjPRcdffsjU/ejJE2G6619DlQ7jG2LlIh20IHqgB3
2p2XOhuGpObL2GYEMpmVRezl/cHkXgFRl7OclsDvwhy/WW/tYt8KE45jPcy2Z5nk9RdditYe2dHP
dIF88xG8slLD+gSF2+CQmnmN4Fi3XHPAZtp/BUgL60bklRin7kq59tiaC8Gnm/71pwGi0cTruzkW
Da47fpztaOoLo6bpx7f6hrqUM1pEyO+WtS8DaHCiFb2oomah40lZV2SBR3RtFy+S2M2P6xOMw4VD
tNF4X0Ftyaz3/kllMMGVyEKl0N4tcINauMUDCZlPM/6IKYn+E23hstw6l33LIz2ETO0Aia9pZKEz
IK7kdwvqqerY5UqMgBWqn9lB47Mox1CNPwQJAtgig2RZVfjczvhp4g4FfJanfEvEw5YpjQTwYfDx
mng23WSmCqtvKqe6Jt63tOqbgwkMJbM5SdDeDNCW5MNPocPviQaLRiP0/Y8J2MnTAtjRXSvN1L4D
zkkkODYlpnDueL7uL7b8/FrvWmJgEwZONMci0vOgRhRT3zPjIL4JhYdfMv4eYrDpOKPtxgRZK2pK
osiIPWndPWCloqO9AP9aIyzcl1oh354bTrSEAMn8pTL9uJWDO76OtASSo5ITHUsDvbfQbFwa+kCd
n8aBUnWPk9FTudjwObTQ+hC2WdmQY0xVQWr0G+ffilUCkCTpJnY7mD8JEJO51kELX358um6K/7ZB
twc1wFyrwdeuEHXaGQXuGavUWZeq7cLBMO3ygsei6+KNRDSgtTZxWi21cEBZZzDjX25D6lbTRxIm
Zpba7hCbQgyvueU+YxLanxsUWhdK7IXcdEoc1vM9rqnCuKIpJ7i9CaBAs0wd67mOT2vngmOwbNDa
U+YDwMxtolSuoGwXcGvR9r79qdmV9W+dH59G+8wTutKGqgwxnRx90vJn8sim9kh9kg+1yNLZCsDA
Yju1BoZsxJEgxBXhnL3kAu/tp0NwgV/H3EqLgVVZe/qmuBxjkRqKNFIsgD2dJZnEbg86H/iJ6o7R
eYK6zAOfDmRe373BhmuSY3UbFifAFat7/qKHxur2VHgRXx10dQcJuY3RfeNKDwR7ypSa40Y32Cqj
/WYcS0JcRcpK2s8s5L6havNE244uOpIX1KbEtj5ocDSw7d+LpDudmzVvk2vxCfbWypTeSrIrGEp6
sxMDRE58IspuKoqPwy9hBEkXPCejWkU9xBeMaURrMM8TiFoXePOyhmBL+PU8JTvbTLuH66UiEMkk
/0Uj8Jpa0xfTrFJuEWCZzRTvSO2CCtqJvaXRN6Vgh2kJQ+hKTzDKLKZff1YLe9bOYD7jci/Eumkq
YxoPcQ7pKtrNDkJWSnFk5Haa1Zu+3SDQdW1IfXrwuRsgsjFelTgLrHL5JIeFELGRmREZwEixytDU
NUGGkNQnE15+lYJxpnAwkmrocqbRS5mUCC6Xf1dgGS6GGACUQUP3ss9QgP6H5hbig3TmC0BVeLgw
Vv33XzKC1dIZiz7TWbNZT6FNpe65vp+tAk3tT+DBIsvdd51t4euKW+3sH/g1EUjkcAf5VI/aihD1
1KVtaolpCxPktXet7Cx9UmMGaEW6s2KLVCXbqInoObTb8XxvHbhN4e4KTIj1iiGdaT5VtH9HR1t+
OzS0tSbl9vB/i4iKdEd4FisVYPVwoOlKekPD1OD2/6SOCGYZUiCfGT3yixFy+Een1q+I6m90dfX8
c4HEpEwRcxA6VfWqzjOOeHpUIuP5hH3VnlaKk78BRAxfIcGOlW4vPhZ83TWllBM0BANm4eXSivaM
D40YB+wwHiN5EqIE/FORRgDWb97zSQIawjguV86cOwv/CdR6I6tveB9hkvMMNz16U6wdfi+iF7/M
a5BO5p3qdRIL4IMwj/n3ixpK5WWjN4Tbk5gNq2WNe0q1Y0FbbbdsPzuZhdH7AL/lLL7FKnb/vCXg
FR2ReEsUjZnPAr6CO7LmiGA+8ToRaqtT3o6SzxO0ecHjX9sMOlZyj6kFuIoxghPwnZnRRVXGjY3C
VytbzCIcLuyvBNv7tv6/2pfrP7cfpnLonH/WWHU6V0Tjzu5hLg11RYKDneGtz16V6Pis4107lXIG
fmxMT4F+WubeCTckdZlkb11zl3zzbXUYNAof05KeSd07gXc2sNsbfNNzHLti9+TmK8Tt2SufnJub
ALg9aDXhEcvr3MYD9f4kaTR+kasTCdXsohMFFMc7TqJd5QKpKgJz3KVSPV5rT78ospYg5xlG3gNM
Dkz5d68uY60vS5XGSLUgikLOYDntuw4jhqEPd7kHs4oJxvS7d/3ta5lHsXkryE1ZVVCNmwLsvqXy
bFP7Sd/wUZJfhwOFyV6gIUL9jYbYS/ECLq1OGfjJujruwx/MA1r0XrAb+40ilIj3EIBNp4D7zBRa
IPwHAUP5gtUZDFjrX7TBzjkBwhgG2ySFsVwukbG5p3pBEgqx7+t8M2BqsA+z7ffSO7ug/TS1RYmy
a02AJ10MU7JGKQgWlvoqGgBjgRYq1dDyjLyREAb1ebcjb+4Fxh7/L2e+alV/a3TbyECO24+Sq9qu
JgchHGEMlc6+QJj0WHopyEoYD1qbs8CWgB0l5iFFe23PMdBb3YFk4zybVPwUWiyfCEJEdmjjpdOZ
2Ye5hp3BGf8c3qrTUGHwUG9B3/UahwBxbVareq/7F5z9EFT2febtvkdZUKngpoeAiCtcH13niTyn
yJcAydyxwbNhafibHfKIJiyEaLb5lTaRrHTeValLXYQ9H9b6YcggoAv+vVkaOn0aEDalvV/tTZe9
Lym0fLuz6XxMxPFu02I6cKPj5a3CNFK3vXV8IOnHLx2D0TZEXR3PbS8faBKx8yrRLekLjtmq3mOL
E2UQzELaCiCzaa68tqkTOCtooynnvrvlWYdFogwjcrQqtUwdciKHXV4QK9vbILaJgBH0SNYpbvjI
iCUKs6srJSHDIPVrysnoRI/8OQ34EsVqWODnPrfIrzx70gQXydeHqaaHZhcWUnX04qguCcmwD6F1
n1h7fT1mMdaBdWOic/6BV9Bs3UeXS/eT5bZhKvQc39LiLL89HxC/LMhKZUW22X3Wjd6OjJ9akGIt
cY2mTSmXLSw5UQC0iA9ochgtvocwdwRkEDgXI54kGJrBhrju5qFprdNNosaZNv+WlpVXHt+d/Ir5
SUyLglMhTZLQ5G6/3dMGJcNkeA8j8PxvCh2EyvtF/0GOCIsjtxTQbUwcemdZzdXdK/g+WKX3E/BT
3NypJLyYTJdbN+eHFX/4dEWTBZ41PyaExQHPx6SwQzxIt0yWPpDJsyXEwptHnf+tVpdNv2W0On8J
xLjEYAEuTH0L8IaLb5YNH0K37oPDE46GNRIQKd/TWNiUtDii0NNcBuyjS0qsGbKmiASzNjjSeg3s
qXGqbm7vdru2mtTKjC7SdY5mEkZS8gOrnpXKhGdxaAqtnUASO4b4Co6lJfcTSwgbbHBLhdbxJ0iD
OjovUHAZZNGJPC9Adf2dWOF8CvVsQg/0ub6rC51TyjkIEP0J/NikwOsr8zbh5vVoroILqkBS65bX
9GCZiuLOh/rkZL4E9KIrCuHPHwWUIhSFC7SXyZJAYNT97T18ladosTQJ6d8rp9dbwIwVU8fNEXJu
2IjuAEWb4imP+p/D/ItnahxA6KWCH4bkUux571sEyiV5P7ny4ttY987nWu/RuwawGYivtzdFSyy1
ZZPpFCbqTVGyDtaVR+oLq3qUM0xyr0bhkyzIaQ2SAO1RpH6z6fWt2MAdkX4K1DOAl0gZHjKZwlac
T+mBILWrHGP1la2O48ygVAqA/2H3UjCiT9Sfz7oYoS+3nGlg/Em+sdpKbikbdDbs+eHziT0F6Mfv
20SnSdepiC0Bdaz107mPmHQ1n14SWGImGL3hAxIRnDBZtc7J2bhz0sEkWVuxFbKf85QcnWtyAeA7
9JDVdrPTMGGHrdW8aP6asqQCDne8csw3Et31uk9a1wOWwoc4Wjg1uc9mT4ha5pbGuNTw9KNocGmG
7wW83ytDojkje7+y07D9l+6dXkuPsUR3Qx9BGbes9MOXuWUvI+bUGtPEi6Pdpq2IvD/1KZBQAUsd
U+doEcGbmbykOrKQTp9qvTfI4A0fLmQcZymaMezQdqVt2Olp2tpUE5omdW6ntR6KXZh/oeRW4yEM
9sB5+WpIuW25C5LqYRt8SPUu7iFoosiXmBtEba6SPsZu59LZH+1dSfgRN/1UrxHCeQFe9IkiD4Vz
bLqg/WoB/8wYDVsAkPuQdOg6pXAib26/I186Y6vzbRJkeD6+XnLmUo/qCMIUPi76eFvwpItl2RAW
I1OuXdv/sNQMyRnDL9Zy4kMByos5dcZBLfb8cxnjK45QR6NxX83XVRD1qc6uVSBlc/+zT6eJ8dFa
5z01Zh+e2ErIW1u+WV3R2IMoAIVOqODcoevVIkMIIt8aUmEQkIEUwDPS3ibX6ZeO2Y4FuTVsGryy
oh/JXKZ1O09tbfF/7rI677mqBBIN8+XjK+GMTKcpduhu6fImfQKwJUot7OQjqt2AKJy1G6N6IFct
VKz1N8WsywVt+dcNeyksQ+KGTBU3kINo6/wdEgiiancjJOZOepYUwBYD5QPEVOkRVxedSFRgCTi1
kd7FAbCL/6dxFSAujYINt/TXvVo0glb8KQm3ETAB2QB0Aq6kLa4efuBM0SRa/HK3sMLttt5swO7B
Kqmj93CLC1jki1gMwuT0DfYZCFAnLgf+kOjTeund6sR6AMZj1p64GaqkBxj95AMJZYFT+Fp90xpw
S2bEegnCSnO4eGS6To36Rlg1qIsHkVgEr/lVdW3I43eH5Ig69fnr9sjbPUn1OkmVo6QUU0PEVG/r
P0pVl8LR2EK/yTuPcUxDKEpPpZHrquSHvzLuriopjc+LuMOsaKTeAdjpg9pdoSFD4SXqyT/niEFI
vwjSTOQwUW93SQcMC4spWvpMBuBgFTEciNdWBGBDT8U70+pCWTl6wElV/rnnI49zBKNzjR3irgPo
2J6SkenPhLxC+nPHonu4DR35fmsDqcag9B+hDrUmKkcNq1aHuEzXoMVnWKd4257e86hI4TZHMaQl
iaM+r1G5ttoj5tGss+0Us6ljOVNP5CvyMIkEoRlWQtnJB/BZ0x3ti/Ot7EU2WDFiijURfHeA9wGn
4Ay/81Ox7FXGuwLkGW7OL06FxxH3qrQViftaxgoE3oopwnGvMCKtL+K9tAgY/W8x50TeEmYPN/Cd
FlOBENX3MP29+nS15ASFaRfctkhmG+KeBTaARzKsDaCRrSFhUoBmPc9vX1hM2a1EVi69udan6ctL
+Lcw/ft8SYBEta5j5f55/gYdXMsDAj73+CuItllNdEGb/MmZhDu2ZrUzPxvJrJleMx8u3c76ujvf
AEnHxVxsVzw83athD/dg54WayvP1Qb0+T7jh7bgyirHC1hTvmYxfDgVz50f54vB+ioC8e/52m9gd
fnJ21or6pNxr0ZwkMvDClP4Twvo4itTWiNjtFASwwd1O+d/+bUkm+N+eg+eIHROdvvTOYGRfWc7w
OctkJQWGcBcwi69D2Hfc8g1YIbyJOGFqEqOpzGac7hdOe6jdHCnnZ9mJE6/InZnMe9PKTzHWUrPX
fEjS17ztSFPWsPqwbnadH5m3UPUntpDUsixCP/YXW02a8ZtE/Dg3+J0DIeDRscOou8/NK05NnrKL
2I/ub7UUbfSVnHfNSllUzA14pTx4oxhux259Ol1yXei1//VHHD6PSJQEhDxblFfjjICkRktw1r/d
FjF81GTmM+CrGY35Sdydl7prfv7p+jdAp2LKxcQXdsC8BCtCH5gEY/czEWTcRbiO2ySCnFEqrt1G
6kTD10iTkTJjmfBcNwFYd89r5iNHSEZXon3PgSRG3kA8bOI7XZPPm4mprD5Tnj8+9qJGyLEpTFkk
Qu3MMv0N3Lwjsc8DpZYnndPwEn798jvHguCzkeMOgLFVHo0IqcLG0BWFmr9PzHiORiehJJSIorDs
KL6JWnmGxs141pWhm6H7NyGqYrpj62BTjXBrWRnd+cSNMEU8B9iTHm3Vvj8MMcFWKrhHCFWlt8aj
QzOyZ6DW0ShN0KrU5jaGivbFQ1Dn5mdsGUjbEBw5qrs3T7gfZ+hHX9IymSWj+QHEKQ9rs85cBH6z
x46HM0rnpeAgkURXZls7ly4jBbaZWeJHBFiuAk5/vSCQNyZBUaRRjt8WDLBTCAsYnPei0VQCwsic
b6OciE+2N+WpX5njN4e5Rl8g2W+6kCKMOmWHf7z/Sj3ycmnLqs3DRQAKXd25q4NhVn44B8kFw8Ag
tRuj6hTyYnyRcvI5dfT+GD05sHCdwmWKalSJ6p6W2F0YNI7jyYXS3/ZKBEb1kMqT4t3HF95X1l8z
6gmszifM2CM16mRkR7CnH1CH8AM5y8owC6p7d4cXiZcCh3uIWsQ0VtkilYIPxaRdlDmNHAqEz6RS
hfUSeDzxPBV4SD6IqBrpgSX2TcKHrQ7D3Cbfe8maijIWaXq1Ah45IsJ5emc3jqzspBc29CiV7o9b
ZZAUL81MEhQFnwhbTzDHXlOvZ1k+KHHf9alTQFwk7NDz1PVjEr5uX6JnxieaWJdZc4CDD27w0LPT
yLc/MsjdiPIY5EJ1q4yBtSsWf9BRBAD1gTfk72rwDAw8jJlwenyv9N8uIEpDp7cQtx5aVceoRsfU
eeZYQg+da9bD2F9Q2KbEniYiz+I22V+GX9C6+xShg5/uOF2Pi7S6Z6LHSLXVvF9p90oOzeJ1fjv7
33np0LiO4Y6qvhLjb/ONuOHx1XkKlueRl5zIJuGqFA9piy6BNGu7WL/d0JhuFltW+0pITssFMRbh
xYzdYjtpSXTlWoYw4tZs42hqcZ8lRe3x/n2+CyGOw3LDxY350kBdxHKqWHLG/ZIW/BIVQqYxx4MV
T9yPI0uGFcEDmkSlOqIt7VlUAXeIYDL+s3y2g8TXsh7Y15PiN7IZJzZgFT3i/q9uSCUZLqx8kCYK
fSzn7sYdoccU5HJE6+Yejm10/pmjgowCCU+CmQk/fH2X/2WhXrwJ2zabi0yoNn8yS7tLPN0CgD9r
fJgY2d5H+D2P4/ih5FtFPR2W1aajsBhiB2byMRiSRexrvrqaiZkmBxoqZfDIyDd0de4cA9zvBOpc
HuIkFEQjOLHuMtKQ4UOcbFzm4gosbdYBt/JXskcclgsokJ1v/+HQdSXHcGtSQCwOlBsiy67au3qP
8jX7LnFeXx3p1pgUJeyp7Etayqo6Wpyj0axSrLp/euNsy6Db+r22jKb3MvjGoA8anfiKXHVjKyaz
s4pg9DtjEP8bbDgHMdbI9jSpEAIoKVQvf94rQU6RzRFvrLHdi/EbYRekxFBNlmPxFRtyoygZmHLN
PYs7pIgI9sijXlk7E30+DlZVS43XEORkKhEuqi4aNRugBCGRSSgYicKe8ipxkFD8Zlyliv9MrZzq
HDbICzxC2ueySBC9YN3aRQKk7z+uT01rj8Twj6r4o1K6iJ6cY/Mj8JW5JOEgbZT5mOhGU9KMaoft
oBvkhdkuv+QSQT1xQ2FdYyxd73xqCvsFYRKCfvQ8DhEooM7RhSNV+p3apIiShNOTHbhvY7cA2h83
Q6mZuEBcekpZvjExdjzAqM4gA1mlUGrBcwPbkd+ACjH4krNMOsUpmmR8LGxIYmTM0e+XNoPq/nYS
bW7D4/QXo36F1vqOYMvdnEuRNiMC/4HzPR7EiCMtf+1PQ2kSLLcSha72t+ESSckWH8eR0uGuvwO7
eITepW+w7ThWooZmbKRDYyBDRDWwJ7RKWXynmSnEgTvaceTd1WXJhA/DGNj9f1v3V3AmxCbwuJwy
llbZtv3Jc4qGX39lxFVomfThKNnROiyD8IjhyFDEZpF+iLU5VXQzOyTPpbeaIJ2wE5JVndPzVFlP
KOwj6J1wQPjfxBXvzH7tuNpVUsype+umxEqd7m86vpt4FONjvxduhIi4cKZ0f1er2BCgnw/Ta05t
HgCeHMdkbrmYJTLnT573kj1Pq9Zzia1+WDY1aMoy5aDlFDhmkFOfjJCLMetBKDiZ8cH0iasBa4TD
MP/ztR82CnghdDwezOY0Az8nCewDNHOcvJyZstrX/tXnXK5hx+FCu1zGdgFP7ylpdLRxwL0XYXJa
tGkwRaLymPgCKZlpUDyuQnFMG/1dQ31VT70g/wKtpyjHhXMiRo2x/kyyYl2QIGDzLKyOJb9KQT8k
zlUkjxQlwHSk52GqN2eV+/Lu6pKSXeG95ixh6SEU6cDrll8+cOwE5lCmV+kZil9fYbvb87YTyFK0
2GGNKsfKLqwV4RJt2Jcu4/B4h1K96HpjlIrWNfrwkm6gi6z+9eh46pevctSvQbDeJLBer1SDtdzn
uWi1DAyvRkHIOfPv1aZUG4Q//PK0v8BeGsIFfrNOCJ3GR+NB0hITRlEA9341H6+aAqi0IlATOcSj
Y471+H+v2XzXj+axIKtn97kTBdvPctybDJmo/bzX8n3phL+U9vgj7Vhr2frrpTHhU9xgslZtoRaU
tYTl0kwRc5gXHkPtSJfvr5pP1umk737fLEicqgEDBpK6OUee3FHc+8gjFf9y+iKHiwF1yYYJLu0x
CuH/gYW6jWYsSvn269skFCFaW36uwd9mRkRgO+Fkz8skV3q8+A4AbtpJlDGLVZsYtKlNO0tw+ISi
0KwX0xRTgtl4nqKJvkdiSZsoL/Xxi8c6gOJOZhljNXuFdne+heRvqIeMyEZSs2hef6LthK4lNvlr
+HMgordvJ2hUbeylAKvLWZYBXCOpO3JuoNMfL17IC6tybIpv+S69ewITNmhN41n1k2IYQkrHzB5Q
DzKRsjW48s4aBTw0oMW/c8FUd/MFELhBUY3AJHUFih6vqG3bzI921IkBPWCqss8pomh9Bc7bvukN
gndTdHLqkgqK2cgQpAgrebT3Ui7wKdXmMLDoMxHnkS/D3FU6fWA3tWuxdurk10tEf9O0w1iU8oLF
TcDmWJtkI5V4qQoME9zY3c5kqAXHz6PVbBKG9Arz+x2yExPDdok/jS3q2ZEOuEqDXSHh0kF2X6F9
0NnsJ/bTvvaLs34yMDzVf6lHxHgtLdOtDnj/4I3t7Hq+7d0XAvXrbG61drp47wONmesX9TNpVqMH
bMjMlk62Xu+j+1tvaRUvQot+QziTHvR9te3AdWQqOCU6MoQkqXg8qucbrgBsKQR8gzPzY/huIYN5
dsimRzq+E42QtVfn04gMXJ9jaIKYl10tQmPMfE9Bi6aU2wQxwp7QMwmDNkpIpVBBnFH/LwFPOS1V
KgJhSsC/0pZtrSspI2UxJLpS170dbDLNFKO46m6njBtPB4+ZjCR0gTUO0bsotS+SAEanCqLflVcX
fGlf/z1ngQIsryHpSLEVpeku5LpBvWlNrZxLj4SvsJ1fLXh5wXFx7re0sQsngBoclynf4I2VLbNG
C7Jq27mlXtt4pzDz9K5uYtLWsKK0+3p5Hb2NVSKmJbqO2Sg8bwd58nqsiBf3eafJcsW8yptaW7TT
t+mVdIbmcoBpr+QY1ISDv5MGxXzEXOyeh0PCFRQrZPLbczrrygdgdn5UNUs+ntbWct/+JaXx0jv/
zX6GRImP83WIX+TXHY9WjWZJcjWE2TtZHstE/uZtctPMkB4b275D1McIzlB/FcmFTIACk4dSPUS1
vHGvj7pKDuOJ0j/oP4DWG9S/OkfH1EAbB7UgtWkEkeye48sBkhAURetLbmEBIBRDwSi4Y5eLsdeS
IKB5tZ8NEPDJeYw4P0H7YGvtP8j+pXS8lNxmwM0sxvXm6FpF5EAx+8Kd7QQiR5bgaD5/Rne3kT2W
1cNEYkLjHpIn9ATV37fA4L9cAlP+Ilg4UUVs0zsrX7PsKeChdZKAdfl9WLA4wcXpGFLYoZapnFYQ
fTkuPvD3ApcvIM7xr2JvpZkch2d8Sd4zr3hlOr2onnaUK1ptCR6+hJSEIOuZwpUxsbix4u4GuUKx
0TqaPednEsi2x51uPeOkZkSvTnpR8lupLL/WA2xN+7Gzs28MQKLLRlPi9OprP1AoKoYjflmdTzYI
ptuLb6xdaUL3AXLe/rd7vj5mq1cbFt34fleMXKyVaOTvBUlpCSsMJ+Qqf9UulmrjRyk5jMLq3IAj
Xx4VPnQMDC/H6EpdJneth3Nm5J1GtHtcFA07F5n8M7Nen/USu/4hl89hnGt7u5zdxTZr8PS+ZRQ+
fVNoPh1zpwLTcSJsc8KCiJBkamcTwC9VrM4TT5Ei8k8vI1Myo1EVGED796yamgK3Dgm6w3cUkJVU
nzZYSd2UGYM+MzbKBs1aRYGy9+WU7Mwey+fm29BCoeqfSuoNi54CoAeEZQnCIKYc/LbjVMOB96EM
5M0H5W8EA+5S/UGnVFPkeermkULpeJQf+2p7qzmfL50AIea6oxQ9wXykpwvJY62h+cZvWjUKyjQr
Wgl+7U/DoRXVRDfMC48My5Oz5HBkIhLMMHiv5hMeatOzVfMLTttVN7HNYZTKsorzytPcs70kaRXa
F9X+DU0tklVPoSpUFMNUsFmPnHdKtS2qYEWxJf2RRu7qkyvoAI1c/QjIWh9pUkwbcbvb5jCxMdzb
A71EhT7GVaFcZ2ebLDxFE4f+Qr1ZGikQw6o5lYC3eMyZ7QnOMAIlqQpvwzcdjarUyCU38MqHsqrn
vymnsVMI4VW/t5yWmIkWnM04cuKZL6BDo3YNdDcSjv6hQVoNxdZ0OHiJ7W2gwvYxuDjveWeXpTg9
R6KMtDbjRZhlYc4dSK8WP9ML6hF0mKXn5rjPGAbZl2JFS3K0uamUQRdcB1cFFeSFJSY0ZTrpTgPx
PUZjrfHno6L1e8CQL/XM/Jm8L7yCzLjhkrL+8mXvTnqwJQes1z0RvFFbaP3uVQZmTpb9pwG8f5i9
0PYGXRdsaU7wjcy0Zts3cKi8gxwNIBvDHE1hY08Sni6yQzdbiqkWvuyUYfwQ9akmEjElVN2pTG/B
S3OxKKLNv1qco/z9cQEYG2B6uTWEp33bwFXKvaiZ5wVOUYodSLox48ljFMFSNB9LPAkZAepynpn9
F+lqFmhZy2RB+Ln78MZe7qcwnVLBbzIeF5x+agN9K8yuICk/ArDcvB5piZlVmU7vXj/iytPN61pE
gDjr24WgS3gVdGoMQDqJyXz8tbgZDWhP5bfnG1tff+iYb53F4Zyp0kuXoCCExdlmNF3RyZG+154M
lk28tGzGCOkGfT3Wa7oKa9vTyXeQyu+CLL1xjDyJXBiS6wgWcy7QTc1fVxjyElPJk6QNRgkJXaG5
A4jRC2iQ87ha0IqBN9h7ds2tGP4cpFln0c5nSkh2tH4wipzGJ+cvb4j5uhKrGHCRirpLkLjldnqK
qtlTEjMrXfHxSSzej5ufj2sp4gTeB+mf0xxlr0MUlUJvY/WF7Xwxfuoq2qithzErm2XmSptXpMuD
Dm9hQDzZPvarjIiaZbCpnpUazrUImUjitNN1aU9BgvmULLdnwl3D12hESO9YaFz2xChs5zaxeTbF
gpDOoFOhysxmxHv/MMB5X8seAjWx8wz2qf4LSPf30MYnxfxMTrFYpEA3hz952owObizIiAN0JnsQ
YbyWJJ7oOTgsS9/ECNs5y0fF0kmoNkEwyAsQZehV1h8lpLiaxLlz67twqGMTFERWtHcAoIR03U3D
Khycdf5ADSMU4FfQ+BHIkvwB6pf6xzCki1JrV4KF4y0tOuqFXhhVR6HIvOJPIhRmeyaSWSWbpdDi
IoUHczF/X3hDa3MbQQWf9NkNIocRrnVyyI/R1n3XehQnb+p5kAVwku5dx2A5hCq0QxoSjAXSmcoa
Tb19jQrYapPn9D8k8pDNaCRv3tIBryZ4NkSJTJ2O70J7etce7rRO1XbXhPbrsDz8tFKSuQFtYTab
xl/lY9K6o769eZeY0OIOfkYOgbUyJW8sSJ+ChaTm2O4R8hm6Kgw2zqU3AyMpPKkOsBksfiYMxOha
5BXG7QNBKrGfXAyjCId9m2g+LNt2wtvD/Izl+rc4BfqOmXoboY2Zi8qgsKaEzdzQ0IDvZd8SDxKV
rsZI7uwzKz8oAzHWkPr2FWTCQxs7ofvzP+CqzyS1eDYNm3unbt6zXQmcwSWQg1rk/QePJdfeGbtg
eu+6glNXKKWMUJKaeEGIqHZ8+YOJM2PycjteS3CKHg8WbTtETZ8Cj1QKNhWG6K8UNqyKCGCkP6/d
xvpHXJp+FJzeYwT80UvIAu+g/GWGta5/e680EjVGPlRqKC/DOO16FW/Mz3sQDjLFLDCNCOX4s08j
Y5UNGfhJfZlsmoAgPzlps8M6XAOMNud9MoWMO5Y1rRD7v/1cGoaIUPo82ONgrOnTTbdpFv5VWQzs
fsA3tQ4CJuz5N39iA6nBvPmEcgo/SYY5P2DPMNNDnfKxrT6lCtGhmKrGLzDxwDui4vvaZjHw6F12
Asx8VDUVAkZ+Xww7sOUqe9ibeZ8B6BThAN5L1nRHTDii2GSkwJM+AjrKBk5HwWcaVOeRJ1ZJr4RI
HO+dOLBNx7YwOArnzgLdeHaEB5aMP8E0JZ1c3msTegvLV8eUgowE3aUL/WnnmAOJyv7FwmR72Nm+
9Rc1FNMVwXbzp2zgCui/R9PmWlxbl7cmchjwY8K4exjSN28bHLZolb5f1gsPfZvoPUcuzdpfDseS
PZmx5XmEmYSSeKjvxw9RKgysE6jnR69TPAMBDuaentVUN96W6Mm54uXSzQKyY5zzKvreTuo/OSZB
FnNVLd/01iF/MUY+C29dRr6bqptghIwg1LNsAQyuPc3yeWMYzLAmQxm3NSDGVw9QQ8/A1sqhkWrH
ylNadDM8fZOyzM3V3rDIGQZTvaKCvNsBIVIMCNW6TH7uKSwLNdQJK9eLujaEBQzj/pvlg1QCpXx7
DSlEgYFKugT10xf17uJPJ3zG03vyVIImN1jOpdzCSYdeYjqe0nh7jHtnGgaUGrQQgf4cbW3GD+dU
1MUtvq5vPh5V3Fh2nAuSu0HXj+n4/8N78xa+ioMfmsvkgoVC9a5rtPylmVKxBs62QaZDE15tR5AH
EWcdgZQU5hArlAVeBqEU1yyXzKjnpmwn2QOjTgTfA9Hbc1CMNeHrxjq54lcgrbii9bhiJIOnZNLp
gnxfUDOaCABDZctUsa4cIoa3D9m7FuQ8Kwstd9gWbkZze/YRoQKRISMtrSE3rzmPRsLBcFME2Fud
0kgBrRuWlpKAWem/eiNW5TUAO9g1CqQoPjXUnOjlMASx05FYKjHhEAe86UuM49xAcic3LkdikszA
i841S/SE5f+Pg6Bj33JdAwe8dnuebhxALFUhKk5Nw8c4T1qUFJVrXN0iZXdsXFmKLgT0fgxrA3+C
Qfa+SEqnCGynegHjYdZpXc1fC3KF0ut0TAJ+GO1tjSdpmldyj4OSdUIWvK+uxcddP/aP9ckGLOl4
D09Xr5q0E0Is2EMQPoas8u4X9snedKUH3SEMQ16s0YaCPdGeeWFCir+doSo8WUn+wqGPolkSH2ZM
0P/eCqSzYm9GBxOcYf0MkoRZo2ifuUQvBeaHtAiFOPUJLhXxGVotb6f+ZZVlKSZ2kgL9mDTtd62R
IBH69CHu2klvhRLd8rGEsTEq2K3lWbsgh9pAHGYvcf7NzCm0ao/0E1xH0dIP9Rcv9f7xqhCXIdlj
DzMUyQtq/thak3WowVdNzVgTeronTyi7HCt5w1FBn2OcHu4/sy7p6dInzgbrg+L9Lqke32FF5CJA
rYIA9wz6bNFIOseXa2zwZvjIcNHSfdJk0T9DKLfpxDTynWUmBUAMYw/CQdQw2QOP24WD6BkHJX7N
8Lwo7NwUu62k2w8r8uori4S2O20BJ+psSHbVbgCrnFefPddP5MWApZjNFnNJJw8UwkWeaPpa61HQ
kiD/hbnf4wVYWUNBDiLYKpYw5kT9Jsbu7XIh7u1sbRqUfiCctxALNTx+Hw8qRpyd+oRH9ruzr2gt
Q+C8hA4PghRsSLB3GLWOTVuz1Ux3L+z+ZFst6KJ470QvRdjq3YyIQ6K+bhM67EIwRBHK+h01Xwlj
kEouSjp9yyWOwpDfQtiTh49u7H3Bb0AmFV2v3eEuQvSszo1LnDVghhkki6u5rbIeAc7m1JA+4xhe
gQpfiPBRAvLi/sKOJVDB+bxdn4sJNzLM6S0v1U1WNottl/VukcP5nBghnxtEjsDCm3k5lWoKgyLK
2hL9JtjSALkCDa88qRwvBEfIIYIoBpjNqt6jianVOFLDxiQmZDqH33P6+rQYjnXe/r1vJPvQaDqg
j+uEvazpDSEiFYNugOsAp+zug2TWi/IRHu3UMBySCCGyv6kE87/288jDJDP+66P6HtWxNWUM2aAZ
1slN0ifvnC/8jKczaUyRrWy9go6TfB0Ne4zFZ3rXievqF2kC5S1Bp5PmFeapq5DoO1t7CNqKCxal
miaCOuPjE7WDOf+kthSC8Z2nPzR9UCJo4dVTo8sc2bs13r+lnCMdcOEAaCLa8XczNfiJzXn3NzGc
m9shj4JcScDFce3Tj9NCkKhnoxIe2pSrutgEkwEjtfdXQ+8xHadYKHrp1AqzD/YoOflG+Wdeg7nx
eRxoe0Fy1f0oahnisY+DVuZOxNONFh9Vs131Lv03ALTEa8pzYtXIbO4eOs+ebarR6233kQwN2+n0
/0wI7A+r/JTjP13x17ii/4514ma5uySJswMgE0tltpeE87AvM75B+WWtHS7TKa++/yXhXww9lNr1
gTFTtybp6P8Jw7IYpJN9maHxPuSXQfiFr6uBj9fiM5owfO7dFLrJlAlUva/OfCP9inrjKIq/FghB
1s+bm9EUxGpwmKh39guu5vnrY9cWwtHQUhjOi1b61nQ+9JhA8w/XqjpFJ/ddRnpoAUA9wmd/xUSi
fUsLERiopa+g2OM5gkhSaS3eKCLXI3ckslLFGrYTqvrxfDQG8r/LE/eJxZF2bPrU1V/U0Z25giu6
3giX7oSVLtKn1HZQ9XqUTd4f3a0qI4ZPAhuqyQwceOUshYkNRGQ42HkjmmewoLGEns08v2YjYqCu
ois+pZQ0gh/ZOyUFKobQpK61QfyOjRqhbmViEB6fmMxLexX03/GoK4h6qkASLngyWDuXK/tro9yU
42f+wQZYbolqOMrqNHKjO4tSB/3h7ZlB1XUlFr/v9FX39v4/oE4x2F6/ToXgv9ziSPKGpUDc/x2g
fhWoJrpgs/zPEIQzTsJ1I90dCAuJH1iiA0jYNiE6LHWB3AvuJ7Lx5/J/nT0roAo6SLAJV7JhTaHj
ixZZGm4K/2MHlFJUModmCUJyu3AQX+iDBGCR+LSHy79B2eyfOHQnIfOloxdDjqopS2UGpExKK5CU
n9x3fvotrN0uvkOFKy2hNQU5xWGawTsJ8MRxTd5I4CJVUxk3JHwycKNFmIIUw4EqiOvpiZJijzfP
ocrGaaWb6z/vs82GqN6V6YKP2syqLNP0L193vtgRH6QEE/TfLN8HB+LlB4sEShtQKeaMEB/6cdLr
r44ZH4IPEgwV0+5i0X0Jxomy8tn8C41fROufQOCw/FtEkwtGz4vq5+XUkpOKjD5iZ1N5iJDK0Tmt
bC3tl0Bbwq/oUz4ZclDIzWIhasktPtRNA8B9Rk/hasDImjwBX3W97Qu8TSzr7Yyk3mSbZ7B8X/FB
DNZKS2a0rxg7v4R77eZ2SFYk9tXzQ0yu5HusfkHthyPsb+yPGcM4ZDfpdlubFqd7FD9VewUKFATS
M1umUycny+PREiCY5d97XcONlquYPDCsJOWZ4JPw9xcCTdmFhlWcQuhSSDFU5Lw1xJdaoZNKuvWz
vSd9gC0TSsLv/16w6esZ0+iGk92am4SOnsHFMyv9wM1zH2BfPsCHUzWLbmF00VcYX2yrZYESDEVE
KwXt9eaaGJH40XnVsq8C9M4vgGYu+7rG9qH7XMJCgAbgu44WqgkQKBeATAKGa1vSuFpKiy3ydSQj
1M+Dkzh9KhgtmwJ4TPMz4LJfAedTzkTwUBKYhFiwC15+DqG9MPcHQO58ZacFFbk0yIJbWbwtWeKW
hnjF53fmjUj0Hnst+pByVRX4Ebeki1MO0jNGxPuFTG8Mf/3OvJAgyJpPVOpQOOxPmVaAQ6l7Lad9
D0ez9myM7RbxpvGGhT3zgV+BGc+y5j5yUIft+dSOS138qCasWfVhPEEdzzZXbYY+IVoHcBAtbFem
fo/jc36whC3bQlDA8YbB7G829rTvN4Ol6pm4oeOIEGw0KnEbjH5E7hnbbnSXIY5PFofJxaLUXlow
49gU3Odt4TfCxddBb7itssIFViuJ24uzCbdrEZ/kn3oCr/acnzxJ+sQGE6m9Rh6eso6aUKHw79ON
RozzJ3nL842YyuYRe0RNh9DzllqO24vPwuiZ/jXWovx2AaxETvGj76SHbIfi9DxxWLEr9jNirU0a
DOkjn7f8DsaiFbwpC8f9x9cOTvQu6eEFwbONpRT9vlKo7VnUTaH1yuv1AXNR5XpPrmtu8KNacCLN
TigrzTOXOtDUc8Jit5LpYykfDkfG/+Apzfk8ZC2bueZE9aDIR36mp+KU3rnhUofWZP2vokpw+1XT
j5XM9SO5m0eeF5WNN3SN6AvDk60lyvxOpLrwIlOvNhOdNipq+m0syDlOFQgVuwI/cfrQsL+dvcRL
PjVW44szvAKnhbpX8/bOfNmv+Otp+twVv7yJJA1oJiWoFaMqgLryQKQ9CysI5js+yZsoZiqZmN//
og5FycL5DD2HKI/L9dCLthxZ4yniwy3vOm+LfuNs/9bTZKCS4CaF0rhGj1N/aftCTsUa+7rAzgeG
Y30XjFJpZBZJ4P3508XBY8/KKUs1xJNlJoyeEetDOdo8Mt+F22YwXbRhcUlNGe7l/KpwUGzOd2G2
4glXnpsLgLkfQSeivIe3+Aa7k94ArKOhI+L0ga5gRoo1WI1hPGBqm+EX4RE89W/lcGqvYvWvzgJC
9sUR7JpcVteDs91+01oUtORfo2RAd7jzow95hiw6Yl1K1mHlVTPZEWNleO0q0VZLVbBpxvFpILI/
JavNCGpKo59ZZ1qzbYXGXliwa5V4+UGh1IwODAb97gtfNo/vzrK1wLikMMV9ZEvVcO3QfK42aADf
amClUqZE3qxxpVuTxUStI7pkhki7bMKj2qCUj0nNJ41Yd5YkMNUGmhRXB53i3WM3eRpQoyDzXpc3
av6nvlTB/G/wcdv9bLrF9CMYk0O94F+dz33U+y1riQZIvbhBalR2xD38JXXwBi2zlNsm6795ANJb
PhrDb4ZLZl9PaUxm2rHRv8rU/ASiC22hRz94a47oqQz9lvrKw+0WK83aWXC4tZyEmRnMpC6MHg/j
3DCpjODZc32HRDOajMaM021XNY1sFcyVw8XSaVNzHAxVWv7cLFjSoZWICU3pZo2AqGXbdVfQVixN
O1vLBiwSvJ0Houbfi3Vbw9cwauvAOF/rR9AZ+IK7xTWlwzbUvEgOQHO1aiYQq8SjsufObUUd3g20
vZoClemJ3SLUeIZvIaxJtNOYWjpMN6vchlW6+n3hXlOUtx+6IGxpbA9BuxG4p9TiB4rFxqZQr4Fh
+7ahkIpAdhge/xpQ+KuuEypO+Ts2xqT002mMUXx3nkYPL1rTnhZlc+/vCh2jOm/T0Ku0aioj7Dek
Ec6oebSoPaASup+lWZAleYrHSmOPdeG/aTuDAUpz9fTwGMAdPsfI+CZSRBnALAQnPQTpRAaBePNI
cMPvviDG3rJ9nkMrPPPe926C4CBhW4FYMmr9iplwMArFHbQk8OGEyeM221myGsIX04N9vk6zX1sp
5urQhQfRpfUsA649/NmKA7U9DszzbWD/fYKxAQgQEZloR6pe8veNyVYhCzsJtgt8WWHBK1+81+Qb
L0hg7iTjKxZvoqprbZ9YUYTS/daTx4yKUl+CuqObmI/C4Q1O2JsFRxFEqNysEcMLnOdhyRTc4c2v
JvrU8qNOkzoWx1YNIBLU3TXAcceUoX2/onOfVbJdY+JD+zdL7I1y4pkb33O/+HMJPbNYZ9I0jMxG
PNVz+dBRe3Oa5qnSru7plcvCCkkpBcBB9sS1cqD8fi4NzXHIrwH7Og2YceOfGmFX/HuzajBbAfr4
jNOGU9D+TgXoDZG9XFy01C4Ijtuvn3QcFiCVL074AFiDmCq13smD99cQ0sW+DGO8H2z1wi7MCRQo
0Pp6feReuJN3+m0bsO8Itl+3VmrqcbmibHV+KDJhv+G9XoZGM8GVr/92tJT0J/T0D1iwl1lWvO13
GKejQ+x5CqCqT8MQ94DcTtbzglSsPEZ31z9k3PCdpsJkRWlSmDnBzXzAzXZrAx3cBV/ONA2ote9A
zFwgrOWtgpZNs+JkaR3MgVqy7jGKUWW+ovd8u3+6JsksCEoItjU0BFqG7Jo21cMolAYVZ8SsiWbI
ujeuw6wdyb4zrRqMN+xF9CpIzwmiAy7P03bQUy8r8z988bO6T8Qa90NSHRqs5pwn2tbT8JNrvG6h
M4Kc9g8NOY0mQDEaZtHn1GtW0lgPL0XLmy74aUb64NFCjNNy1dty+nHG01YlfJ9UQYPdV8oo0UIn
a67lRi720VeHv5Hq1GDhOoPsoBAgAlWXU5LxBrb7p6RjwQWcidmnehucopclA3WU7+IrRyaYr+Kf
z7vbfKqMdhoTzo4H7PNyeRNDkvy43cH+mxBv90V13clwMsEf8ilbD6AjWH+AKA7wp6NoBxkPjRin
8T/ZIcvKFJzawzeh+JNv1s4nfUlZOgmCIalDs2dh+uSAUs8+HcvlBV0UHoHrYVWg322HzjWGw0/D
dchZONuiVsF4fd0nDCReRQFifcmh8iJeDfRdwXQiU3nooBTZIakQE5LbniLT2HR0MIaPGmfPmjtJ
0I8navdNCtoHEY39M9sRowpHLJolhIQktMeFlTu2clg+lczlq5UqNPTGXbmGnKSzQoCrEUl+9VBD
K7kMFefYfnml5ewMWXAcqUrqtKCVySIcCIdumw0l5rwCrSqslIJa8woR5BhwIhVXEU35KmtcZHFE
CZEmgFNYUHKX/l7v3JOHcWOV7HX0MPzIPkVJOspVIOln1HIGa3xtv+I+7BZfmu/OXO1FXjvlNGNz
UYWF02b8zqSDBNaYc+I2CtALZTB2lyAKdzY0oalG2C0L5yqopmPazmKCeoqVsUL5FWWHNfKLVu6H
GrkMnWlji8+iO/HsctUjBAIIEn8z/ro6y3cYzC/FEvio/cSRTn5sQ7gO2yFjAe2EKFZ1lI0zWrWc
uUay9icex8B5WsKQbDyuPtjF9B/4rxsI0gsyccYO88BUtl3BTw1MNoSub6dti6NCrRpdYYdKJuIu
kG24My0FHiLXO+Yv7aVnwHpcJDujONr0dJokCh997T7rUYTNQzEN8QrDsataH64g2zU6wbSkYSbV
5Dbg1dmeD60HFMKREzNNP3JRDqHejg4MNF4vK3S0iAV1YmpcxXKFdsGqc36UtM/5LFhYeWnRZ0dq
a3MaETryHICFq1y5tSE+bX1BdiBk3lwEDttx+svr8K9/m5nrpVg4SnYhOmQMTlg3bSdDPF02wW1O
gnQEWI7BoWet04csym6e1xwTVW8ecvEZtb6KKdNhIk1QvPYzjBUpkq1hm+0juRFmeApTNI4oYTsr
ckL6LIK1o4GflWFTsgPWYEYuJgPUdIzfNFpPj1R77SQxoC9K2tlKZrDSv6mU6JupxrJ0IQmPhvmI
Pkl01dk+O/J8/95KDumt12mSke8EfWG9FmS1+Qu+kmrG8E8gR9K319xM9lFAENpJjZwmIaijVRiu
8V87uNm+ow9BwfE+ty8LgFEgic/n1r15xKrD7O8qXgW2HFt1QVwA0yJVtDyQt+Qb/B4UTh7FgkrK
qVRKA/X32zTj3Hem5g6SKFOEVX3JpDs4MnqThCgiZHMptud2aDrvKKPsUnunz/Z6t8J3elsJNLP6
AvFjdVJetLefS0G2rk301cFsJ6Y84A5GspoPEpVfL+aW7ZX+ihbcflRJDhH4XsaP0zSLwRROEk1l
Qsat8VYyxIC4FUZmhuP9vFC7kdI1qgRPYt6la120O9/mhkYb0+/irSaw2S98FCsb7zQnZbAU1JA4
UX3FzrksY//0GlFL1S4wHScs1rJJP/KbrVC+5oVUE0wmmrGh2UQFmWsj/26k5myKqILDSZ4psiph
54YhdNgqygQhKpfgKPIjYAMMQNHvKoIumemsSch9h/D09fjd/g/lCUCaZsg7PVPwqvb+LqYTjXqQ
gLWZSNud8QcR9nvNdvkC+rG42oVP9VB/LZ6Z+OW6eGUu384RnSiQzbXN+v/VAErzL4gNWjda0gXe
+TsqW9Mir5cLHmTWvireO4oBQs73Cw1u7155aEsZz/XShMggL/6J2SupyVj/GcB311zJx4TgocgM
b7IheKQ2u/vLpbGN14gD0OMp8iY973GYpJmIaoTcqg/ZaG0WhE8wuJ/xepyR7AY7g2BAlpurx5HG
GX7kfaZGG1bBJ46noyQisV8vqKv/wTjRA4KLT+rPDsaM7rzjQLZhGb+sTDpRYq2na5//uABigTmF
4ZYV677mO+Nz0sar4hBbUFRk3gatFk+mYxw9zCSyMYvKXFCAShq5cwvXjlBZ00wuoL6z092fowrM
kReVVo/agU6VXp5DaFXpSeVNP30pWAM1Y2rkRQWO30/FtU5+mKrFD6FQrhy5A0XYJkw42SQyMlOm
MlDtgRwkPA8nZsBFXlU0twRRPkwGkagS26Fub2u8U9u3aQefWQbLlwwDFsfJ8n2at7QbXnySFi3Z
l6zIeao0EruNmPb7ZaUSBWJvf6s8zbL0qwQUQHEEoieQtlWsEftuR3U3QuiMY3AFRYnvi287ry+M
Un9DjzKbix/sZz7WoA4Ym+ieoQ5yiAp1BvLaGaKtHAYchH3nasPe7z0ydekpG1mEisXEEJzZLsrf
nXBH6Rgt5iLNEf6lBdUUS5ZSYlpd9EosxShkccop7H0ZNES9L+V3U0rnGf7rf5XQO+DT3HJnoDmw
Mymw3xkmCzYG76AcVM7/m8DZ588CMzlaSHTW6daEbtoh0sqwA/ca+rGCm4TXDrznItuGbrehdO5N
K7JagsjCOZ4ULdrkecmrrErnYqwvl09OOhp+pNrezUPWWDbiXbLo3rRaxbuuwaWHaf1xB3gXxljj
mdr2bvI75sav7dxcxaqJKiAV0TAYjyEf+ecYE2dmwUdOen+RrtsQmdkydECEqWz1EmGnzn/Enf/s
qhc2io4Yn82O512wjroAv+dhawMWiU8d+AZNOKoeTnOnmRgCiMPTLKmFZw88266Ol895mIGmdvk0
Urk4eYHFDWlDJ2lfCfR7hwIqXygCMOnnvy6IHgXvNxFrreh34gNzsiktrQUVDIEmlXFmpjMqN6zF
MeSs6p7gn59Ll/mRvEbdK31v7EBHbTwZ43DffRfEouFR+9t+eMlPdbeXpafDLuls9AnK7ib9ElCt
42CmeQWMJs5gostyFDtGviIPijN38n+wLK6f/YKrxTCAHQa4EJEUZNwtWPQ0XyXN/LGpPxjFlAfr
M3sZMILQM3vu5kyH2MVVvIiPaz/Sbsjc/g1lzNOfwujDi3e+9mTHl/TRpvz46PHhq5pmkVnvOQgQ
gcLYXEvmunT2cMuhAm3Z37OaSAQN8OPJqMpp4ALVXSp9TtryLiCRHNkRL5wQ6gSjw1psKt1/T8rd
BQToOV2s4iqNePIve2/R11fUycUg3+xHTehv965plEsvoOof62hjZWpPoxyO/RT8AEnduDsD6POe
EyRd4qeg+Sz748x+tWMWhq9DCT4ShX+3h2UivjvzallYYfndrLm7SnRtfdT6AKcMVVYcToPBtpYb
HQmbmy9ZflZJokLcWhs6KaJU0Un31O5TFJalSp4WV4SQwzn31TvdBjJCB7+3hKVpAJXQXrBtSxtu
nlr9LyaqrfjoM7UXnCVPyLgv8BVFQesHGv//eldKVBSwG+FqjQIu9cuvwxgT5GfPZEI9fN4VJybm
N8VVrbYVm8CMr4DtlfwOuFtfCCVFL/KRSPQ0y2bgR4p8D9PbOtzIdu1XCfWmlyyGqI2vJhwdHYHi
H3Jvlz//XDWeS2wAfImZaIssv1ccS3hDnLAwgxWJCKiUOwSHh6YrgcYA68Qjcq109HDWL0nXW8TQ
PK3KQozeZxmDbS1IY1gomUJY7e218lK4uSAEJIKISsfj2wHI4AABWrJgdr4YCAYIoT+UWmUNl381
xf3oF/RIkMJibCVRqcrGOrxDC5rviZuORkWyHispQg36RzBTMJ/KwHwiYnEG2R8l5Vxo57KVlaOw
evYatsHp4kAevXVka5cvkFClFodc4Xwkd43OfmuaqNP1wTYFYinaWMhG3VMNEfLgBghJuNt9x8th
NuGujRaGNFBNG0a8h7amqemOeKNgxzb/Whge1AWqyYMJNypLPRq51V6k/kmELLZB/MBAIKtHhA9v
V1UVQ8DneYoWoSCNlsoVgAcBbh/IhHPv7HaEUaLPsXHRSvqvWWM7/pGOzx6GfkicQcCOR3/KUWrT
K6+NHDJmHcgog/RTAg0ZFfU8D0rOK6HQQ1gm8p0WXVr9kPjxsArV/b3oe/hNuPf54RLAPTzPADc5
10jnPEGXk6y7H7CTvEk7q93Pdo32P2c8yhA/z0LKxg3KmrRIpCT/LUmTe+TVdgNvxht3EU9x+wqj
fiPQQNx7tM3fbgpnxXvOY1kKH+NUJVzFFHjnlOMJktMUHNvL8NIycONl25yel/5gQlLL8V5LIwlk
tEP/8bS2AljWIzvHA0GZBhURc4EdC3AeExdv0GXDiVGM4sfRNzf6qZkGA+pNMpdIkMOLAWTXSJFv
V/TK4Fx4Kcv3ctbzJ3ZX1yxsPMjuFY8zovPxv4S07OmJaW1WIWgGaKyPa2wi3DfBabNCzgG2aOko
twOkJtAnPz1+8UzeUBFk6+NSR0JMXihMn6iEJLKjAfnhIfDaWsD7j1khFiYeNzh+kx8/mVp/IQZR
CUy0IU91Qf5krkDz7EP3+/ZjFs9xz0OAN5NKiDTWOW5gDh+eha8utqP1V0qnQr2MayabQqaSX8IT
t7H66DRczTQa+dEZN6rvP6SJrOa9mOyZHri3IgZofZwTnbVUSSvkUgsRU8Bg7yHhnHmiWIKc8j3g
0YYuj/oC2XHsr09dxNjUGlDqGNqggnnmhR9jqSXGOxDhEWvDW1T6jIGOL8Qn3C79Fmr2DrkTgP1q
IQys4FyOAEqyJ8B+SPuQcCvRNofPPgp8jukFvDnYiYfk9JVg1iH2v0sSUt1dyHzsS1yfySWAzbf7
pdlq9337JcYBXVN//hv7Q9ADEVIuDHZ60/qJCEPpALFkFmYOPz8Q5Su/ZYX3uc+S/E0yNXlJHHwI
OBvW00+djCLF3E2W+7zMK/7tHv0j+UJi9u7CgSiQ51dwHvXWBIpzTxIz1jvp+9aqZFPKcbjsHcEb
hmfA0/dzNPGcIiJ56BpwuSD/W7kkgPQQuHn/5ybLtZ/xwkC1rCmeLrm8rEBw+s9e/EOmW6ZSjbsS
ps0icqYStkqZwu+hmEoIus1fWbFmLRzbAUFetoy8sQpFpw9tR01aCpR1cbYtTHxO13zqyUo/XbH9
yWA+tivY+6aS31FAi1HWhvmE5Cc6BeNxmlWe3qXROZ6qDtjHy33ap2/jspxG8FVQLIEpPtL3yZDJ
muGnrvA2HoTcWyF3iQ6hHY8TQc1BP7U8xC86qUfvdxpsbxQt6tlpmP+T4TsVO2NbIZA5gfj+usk0
/oZ+O7v1l6s8sw3b/YP0A2zOFQRI/6AbNV//eeZ7dYAKWx02rXXmhXh2PDqBHV38vNSREpm+tLKO
CgqMMATyao8cynsbJZgKYoYm6qWPA8NnjRzpduKYlCYcgirKe/gStMpAL45fHCwPQWC1VNu0SQYj
HLntYXyxRzveBB/2Dt/3vSVYiVkyZ9FV7qPyANfc7x2hHZ2l5UIW2gxODAJuopqV7xzhgGkLRyr7
JLesU6U1IvpD9aGvf00T5PVVERok56jCjbyUHaZDzKuWThKnlgPoKc3f5QNS71p6uU15RlZzaR2w
OwHw6xB3qRFQ7tb0/xdD6XlkrLdmhfwxwHRulR+z1CByP6lQvh7dpf3BkBwuPJIJiV23mxEAtttP
LeCSeRIXrMnjObfX7IbtNmkWzRq4dqUGaHxrCIAWQ6KSJPyfpZJTs9VoCJQ+308LVB/WKJSqSjt9
JLnSeMGLUElqwaTVnfy8c8rETujWcLqPV26Jddf0gFlBceEAAh4KJu5cdhGRe2NUrXhofyChascn
wnonz6c7VKfU+DFf28M+nzMu9kfwX702wQ5G9rPOUTMvQg8jY2oWLuhyAfTlkh6Q4V39bUokUcK6
7Qp1Zvu+YnzENyE4TxK8+hL7GDWa2lhw+QQqIxVV2jdJePHcDnEgSRQ1Q1Fgo1P+Cqy4cIEzy4BQ
5nvtnebcEoMObHSGtB4E2RlI4/ArNpl4Tq/7uq3GEK7KrrIJW/XmOT6UpEBtvCjqdl94eMqxFbbp
OrLQg3gvrnPX5bM9Gv/SF7GxBQt17dj0FifazI39Vm6p7yy4bD/yE4Z5H+JKwFUszLCp9TV9wTyO
SsnsccFBC9Xk+1KPh3/TFr9JfC7HW8Xi+0YLrGOr9bOivCKhpckWhFN/Yw4PI77XdEF7SlFjJV3T
fW+humnppBfTJelOPljE0VFci/HNIoAR1niuEETNDiHNx9FBpS5/Aaf2g2JFyxalRDgcVOFufwq+
jALliF7waxaNi3hNRwr+KPA5xLWTzM5QlM8SofDu//1hNOsANDn6Mye1wJJ77ShW65Kw67dLSIzX
i73HPhujZKwbzQ3qv0wh25dgeY5EVvTNUZWr4ZfAbPhYqBY0apc/abEtgKkfSl6z61mIpWTz6AHZ
yLavISQcrNu7P8cjYlg7cf/vGAvioYQj2bElmgTKrAjTVY9Xv25Ma0Mq8IHWwENZ0CMX6jJ6UA8g
2nEUcV+kB39Wp20P8Vt1Cb1nT1GkvVRX2zQg3RPIqvnbabvi1yvRJVGjZUW2FKdzNBSGcvj9P+2W
KhiaE48XGPc7DMjhLl9givxtZsPUvUkQCLxXXqLTAQafHePxUKoGY0h7ASKIM495yE0C5b3gddUC
XKiXr2a/4CIo/0hB4FWa4UAOk8J0Ott6Un0Mg2XMYj5Neiy6zi/qnwVonC0b2U+mio/0AAtmcPAH
EnA1Xz7/B5m/cMjxLYcjIWRmjpDDpkdJyzWEePg+hTQMCAftFbzQgGCKYvfNdNj1PHrBpke43aFV
NQmf0wnDoHhyT9kFJb6ZiKp7HapgEbhPGU7Pvir8pSYAtjUr4AhhuHtnIkdVJKczQGTqIWSXgTEo
/X7dKdT2DZzdYC7jZlVYjLHNViwqCe1Jfz3YqZ+kFIMs615VqIJYsgTg4290z3jdebdGYxBLseN1
VyMn4ahynNV/HGamT4Fi4YtInL2l1C7+bS2E6vN8sCUqGtfFGkryr0YPKIaCAAJU9po98C3kEWP6
BEdp37xfblrxeOYj+zjRd+WspBWGCjI4K14WskxIKoYMRyVZsecNyB2i/v9ihbcbl1XKXbwBacA1
sGIAzVXUXhpgLxQsUNax8gW//pf5/h7ltu3WHvZ4fXC7Kmh7jZgxJem6H1BqLsCfK/dtkx22cplh
PGei4jNFQn0HpJVMivDoZqr49x/d9xYs8UyKD06Vcf0GdX6z2a2nclCKKQzatSdmHKaCg//RgHG4
0OZ19VmNmUMzOMpk6ux09v21AKxofwboPeBHzUif0AraaG9Oc+wGJjSgTP8xOfJojIveWR+gKEYd
cK3dyVAvR6Vg05Q3yDGgQyn4SS2+FDXsec/f8WqrB20+KQbO5YH9KOqc3H1IIr5FZ3q6UizFV9qT
IcSo0uD9XskSEZ2Nw3aoeLkh7fsnTR89+nTt11zMZzacSict2dG7oqe9Hx1BYYRJID1DOnJRrySP
fdeDdjTOBXB8oa5fWJzMb7ZzAJpHQaImtICXmVe88lSsyky1Qehe6m2mAfhCsCo5H0pqeqJfcJYh
wQB7euaeKJNMqcFjjgkAXg3tbAXdyux2iq33Ud723YeSmid3n7QXTtba4wzAjxeOa5iOLi0nkK+S
bnS94X8NDP9yTpdSikMr+FBbEC5MMQD+hbDVBDKS5RTtRk85KwXO5FBrOQxBw0jdwxagqMyMKFo7
9SWkBWI1g7n6Ly6IDyi4Cj+nCHIMlVWS+DGILviP1AZflGM2Z3Gy7Tg7ov7pDIeS9pGqmGYwaaAL
fP/OPkMEOOxT2Dt5lPQizlatzxYDRg4Z5n8JAJQLGnhJGUI5k9NQPwbvhXZleiHWKgzwfIpEI9D5
zCEX3kVYFOPfKds6J0VzCpbFVcLuQi4wo6uKsAJMyv06ujKqkRiyXqzXWVsDmbHrAfWFJxPD2ax8
vN9vY1A9hEquRJP7KDjzmsdlnk2l9K5WBptrH3qHf8dQzVecY2wqAJ4zwDuglEJXFbQmMmKVpIVb
60VcHUGIKoOucI12vgzkrPuY0vjELZZWsytyUuunfc/GlG+JEd4cy/Lxc5s5wc4vCxX+bjmO5Qge
bFGAAiwswtaEymzmxIjr0Ib5GnOW4H/nyRqx/vUCG+0HCr6TilLDDSeeWRapsOnnCNraUyr88F8M
uf3WMIiT2UcV3JKtY818IcLLNllnl14czXEMuBparrbniczecsCR/I7csuoggjugwhWmb5l6uDU0
p2M8j9xOG8ICsxw+w3Jzvedb0d67E4HgiEFi/3kFpImmY3roeoxSGOMi0n5AjoWCGM3xQw2+s0WM
/GBrgBQi3GPWej8VQvVJeBpo4dV6sk7x5JMHvzWXbIoPtWQ7nOARkoJmFhjzBO3gaz6o2QlbES+y
ecnqwKY/926T6pYUBXAPUDeANIoIqlnWW+t7limdqT2GXQnjtiYH649hCiBBsnU5xIXTOpcpa/u8
OkGTo69RIl2pOVIBkUUyo7cbpVzYstrtyOzMGk/nqVpVFtNynzFpiXWeCPSRcvV3g2QLpjSx9cSY
6BvBCUo/A6kDhnvzh1ns7HIqXBIGFkVVsdV+nv1B1PxWdNdUgfoPLh0X+9tTTjz+DnRvzb/VxM7u
xQIBhoOMV3LYZgK0+e5jfQ5OSuJ/I7g4BcWHO0ZyWplLov1UgrIJAK00b+11E0JHhoCrBWey8u+m
tskOd78o/2qMa2QqNABP1nMI6+fAWkWG/ObQqND4Kk7oG3SCgbsXTXUhVhJQU0uDxBW+4mEKV4aK
YWo/aiWsIGtgGCq1dKB1VRne4Rs6XKfByj6IdZ4owyNSPq7atm2lWy1l+vXgI/IWrhv/AQlmVFCI
/RRoaCMKCqqQy0dOiYDWerba7Z3KCeXO8WeZ0VPp3heAnHdn0yzStxUmZF2BlMmao2zNsFitxiEy
KAlSwm6IYiQwMLGriHpW/kxSgI9LHVO332YaCT3OsYuabAr7Y0845pbIcAkwslbExCiKHrcPQe2I
GBOUKK/N+Papipd1z92184WjK5IfZ6SPEgr7CpKEKE19tFjs6E1K9anrSMmydNnya+1hQaoCMXhh
8PK5pFf/OJ8LYSWrXfKgMHNNSwQRlbZEHU+ZMMTV+R5bGqHbU/6bCviRBwUCjZIyE5YJUGkVq7Am
b876Ie2IWURtlELvlcRg20y59iJAOFxrw5QJsRK5OQOIU95jISBE/NpFhfDvvkTQf1Gn4MBr681V
q4T+aApGM4NYwqt1PCKComWoM6DT1x5zB6ngd00uM1QOheloKqfRXKUj+kVkO9iG72/XKradTqRH
9VpaZn4pCH4QcdYGDPbQVejZqzqsu+Kh9hC/0IJ5hvQAdaGvZlPX9ivlwZTZOjlNbyQAMYil5tDu
9OOczqRT+K1YKag9e0teSr3ERb/11d5TubBxa5tM5OYCsP1CIZZiX4/6al4e3DPQlQ2dzwZoufce
LTu9Rtf3bHD9KUIvrn45I8BMnSXHmGuvBYMyi0oyXgmnynUXY4/krM5X6vtPTTb7rr11N1LtuMiq
bi0y1QGD02Oy0dSjoddi7maqkE4DTduu77qFH3RO2TdHLNF++F/d3io6fZMYGhzMUlRn4FXNMUD4
4BxXhX2FD+sFw3X7Yr3upjRuXnTeI/USMklp4VSDShW9qiZSCBXd6U4DWTm0Zs2/TSnbNYV71aNS
YnNiYSWl367SjQOiDGYqS/o9bpzsYsKGNxbq9m4yviklMA8ISfPMibYz1SHL7WOeiNLEQqzCAt3h
U+gN3VFHBdbN8JNGDclLkTBrUojCHwuD6enQCccAfuG4jZ0Z1l09+fMHZ3rEn7CDXf6xD+Mvp15l
ZiFb8nDMhszl956T5hdQz9otVFApkSlvG9hEnkz6+PsRaLXw6xbiUaKKpKA8Slta7YSPMPBsr8Cr
gc1SffSIVMSS64oKefPsDSFsvR4VfrUxV6ia7JuX06rYL4txSzKljMax7BQUokk4HXnDg5V+S5tw
8nxS721fMQXmudHnNC+gtDUiWCoIxToHt9siENlowreH08WCaUYXcnzCYnFSct9/BBgyt5FHnnC/
rFSkfUWlmUpUgX6HNkdDIhU4MW/GgsgVYWndgwsGzKz6euHrSrcQAg0x10frqE5cmxFcsE/D9mlG
maGn7xdiJtCvM+AUl3vR0q4JGfpNCVTWZKijltdBeup/Qn3qPAQGFClnXRqdRQd6kkmptGcaWxRB
pShZ1/pJLa6HaD6fj9//2zeM2JCIQ71CArNbqEfmvworEbdDuGxXZO6VHtCOSyFiSrXFeK7HsRom
wMmbB02HJrrSw3uH8h0qbRDEoKAiEyLI6Npqr3/l2xGKyASt1c++ZzawxC48ubBm8egXcC315SGD
Z1aEgxNg0352jkN+YtSM31+3cGcK25Y+PRTPYUMz20RcWs4npiMLKvApkmQ6s0FvebmwBRRVTqSx
RcUKrglikwWaUJjYe+jvPtX9NxYoRkAP8kNhTkZ38YYVfLz0aVl7USRUX5GH9DHLItPrOzHWMTPP
QQcDsYg6OY3ot2h3JxokQKVTRvfCbwCeVCf9NDPkvucvMgS8HReRxzcOvG95llJRguxS7VolAsMf
JKONdlWB6RkiUWwOun8gmeSPwdKhGNpN5yNdcyHKoBcRiwHpH9X/c/AIS2ZHUlj0oTjjoUYBQ5Af
PwviUo8zePDLHJkRRlmc2ZYFwTWNkAQwbfXLSFbIG2KaNkompCLWIxZPX+llHC+ymid2k6lRAZt4
9H064hxBqk5p+Pasu9i/F+LDWRW5URjuTEo528lz0D2JMt4tHmzAJMQtPNPCY64K7AGcpDx1SIO5
X913c8ucytM+LRhXgz8e5rwY/9keXaSCTkTte18Jf9I+hwDsWGyxlXLRUt6XQHhMzB4iC6P1jyt5
kNf7UwhS9xMHs0TPZx+/OuQQHXn/ySBhcbwvk/gahZXxNEK4KItnHBPK2j3hTReD21pLz848rTk+
JPHuC9ennwDIma7RYK0EG7OcHDkuiXKFu+nGCX2ZiAJ9uwxyGmN5L8RbMulX0eZfFCPu/BIU3yne
znfgPFkK4S7cPOjNtitZTufLAra8hpZ7TMa/7+3MULB00JxlKWqZyyD2cz7tALG9jEhXpl4XioHx
h3twoOk/zKThpf9q1R4GBbJFYA+n8RyUIb5TgQLfNdc62qvDwn0rEgmMpwLW8CvQCeIdvF5XE6CV
UkMD0ehh63uUB4P9g8rTUwwSkrVWd2RdqE36jxx1DdyogH/RW96jHOi10VYBQOGY4vdE/EHTSMQT
ey7SbLkZClsiybWkTbm8lTBb93vcoVuQNxaUoOMMPhCVwfEA1TKWurtOnrFW9ySQNh8/QX2c9X1R
X5lqWOc6T9hSHFy/y2ASAQeYz5Zm9OZaJhaemvR8pg5q0L7paCG4dC5I9a2hFrrxsZbu0GYDkoKm
Vnai7ryPzquYSN5MiIjMtQ3CPMu+wA7/EPhznfMQzU/Gyr4PWCrv4SvSVRZXkruqJMY17rKLKP/d
rcopJRrgfUApzZ6/JjHlEqBrw0zZ5keuIg8m2PB+WnYnXECaHupKUkUEH5y3Ok0TPuLQWjnhTHck
sPcFUioD2vm2GNzv8rVXSWQUjq5O+yUMRDAaAiEEWrqH7TFKHcVBAacx4v79B8gdttMOfeigwkTr
GvHEwR0a2XwVWmdbWPgnKMt1oxaWO5MuJQp0rHLM2XWI+jPpA7UPHK0fHzO5UhlFjFu9zQhV2hny
JfIFLdljjWlNnO2vyByVe0pyDPoVadkUEDlpB4etUpYQ9ArT2PZiSSJamrT3ztvfoMwDquXnI4kC
adI5AXneNeb7/FOn1qL3CUppD1Ncrg63kqotK4A29YKD7lCzoHdKngnqIlgYlI+wafBhzqjnTIPP
5Aob3jMaQ4Pip1FE+urPhgzhHx6h8EWHeE9vSMWznik2Fi9LfMGNCMrTnDCwXhiLIFnopDz5sDbK
xg5v9rE4cTi/A72NbPqNxdCh02YZDpt0JgYUO2G23Gj9kxDNr3fVDIhm/taWAT8uT06iyw1rR3lD
WLZqY6Pe/ErfGz7Wr0LzUGr1XpUpXt2JILNXqwwBBVS3/NHgY2roBDo1XmYu51q02ktfNWk89DHF
bp9VHAbRTuCkMA2//nhh0XNtyOmnOSZScx7mwdQ9vsBAhxOXIS/gyI+SRjYh5P9JTiNJyFrfJyPK
1NiyYVAQtPOn3q8uOxzfxs6OPEtmH3ZC50ydruKPsB8mvAFnghM/zOuni7YiFC6QD8+FyDQHPRSZ
uqKVely25N4IY/9eEyIhIl1h4DGAOwmA6TgauXjW+Cv5EzRlgp/NG4dF+n9Nee38GBV0dARiZ3Vq
mvQfLziBYruVNPaMkIf1LUK5Tm3D+XOaovTuF30rta67CkVHT6xnHfBacJrq8YxPSj9chE3Kmcrf
SS2oqkX6vixR3TkFmMj3GScK2Y9fvqrlRJByOX5rFsUm2fUbIv7CJtQH/Q2DG+PNfvxXqlKFR8OG
MytBStOXWmE2z0haHsir+1ekmefMTNJIny3PRf9aUfqRgeAWQxfE6wKBIOx0x+emHW8x/0K8RD+f
lOecmx06EsbuMr6k+pS29AZ4ArgHwLsoF5d16Xr0wSpyg+xPOIfcFu/PXikB9GqvfRDzYsaawlyy
J+ukx5gFl/9mg5MImzRbvpw1ObrRxCCefT2Vwa8O3JYfTIgjFex+Zd3y2Ei9IWXug+j2NKBlqcVz
eAG7fZJosJ5fE1fMVue34sqVFeMqS2icTB8tXOKkg3H3OJdFEADGz58x+8VfroQeAgW63U8JjurA
PzzUKB8bMYN/H+zFDXiYdD4GbDFx2DnQqiXNRrUNNCGrufTLsT2hH9Zf3NaHmIUnqKpq5wh05eSg
XDxE1MZ8RJkn99pX2QSNn+cunHDakNOzUlH84BjovcWc0Ekc4pCTU6ZVQgYUO8rH70YzGyAsWskE
RCq3hqGt5BphN0tWfPLd0VyomLL+ffHo5T6V/zO5fCMLjPwWke4XDZHI5iORzd2ecKQ+4e/YPH4S
fKOqFw6B6QkkQ77vLOtspuZmezigORxjB+A42G2pIduQ2Xoz7C8EsQrbE6uSyaHK8TxdG3A1REIa
ojzkPBtFmS31oNxDARtAFVTNFaH6ST56Aovw0bfx0dSKsjAX+I/tYybrXXcNJPtaPHdMufK0NpXS
EYe0njhvNjfA/SR0QpGCkbPmGNMAB9fdaGj96VXQTtm3B6X2BQ0UzcBDF3AJuahGdNE8sezD9+/k
Zdls5nmEzy1SCPzJxSrUznqgIXqFs5HXrxqXEBdvd86SSznVT4G83yq9BlyRxqgUKnZ5ZMG1foZY
etljhKfZw8R2w5ALhBAEgHgjOdVTRiYFJESqtfuFr7cLg4Iy21fO6juLrW5F1r3dj6sZZ24vXkUL
Glx80ZOXJhAh0w4sAq5RKcaOwMfleL1FNaCDwMa4txCdRRZG+9vfDXOzZjCiirfGQpPcEr39JazS
sH8J6UNTFF+wi3e5k+1AEElY72IMlApB7Y7XN16MUUJrwWHRGjIrAd2HrkcuPg747GfaOPhZ2stv
XNNieHWFGO2pKF19/G8HPP2xr19fTH2BQDONhzY04O7CRBO3KxTRt4vPi3/Ju1Up2TJLLQhHEnr0
GGNF00sIwNyNV24CUgLGofSuWgRic5Ed4cPk6/cLeWmjVkUhwYZzNBgI+krsn5I0kLq3ht7Y2l5H
kINH9M93ilZesEQfOyxKjm1MTvufjlheA915OebYaKTQgscwtraSecx2AwVBgcESW4Nbso8bOkyL
0QqxrATNHaDwyYHSXzbe38wsgaLDS4qUeXvt2lqeYf+Qe/vcQvzzThg+F1a+4nHWJ6skoWWj5QQW
q34rBq6sBbSAyE4HNrVB8q+L7EOZd51HtFz7xIt13o5McFSj+4qgZFlVWgMJ89gIqMoZ66TdCKny
ye9azf9Xggq+ZmrmEiwF7oISOeKxMb9N+AIX1uCSCw5Px9gEfmBf1s/AWScD/507wa/77ObTDjaB
u8xwkO0YgpgglsTS+R8Ok1kE4alS6UJTQwXSDewrJUt0XoqLblzfpCcGAKOPg4Tnxmrxj2YO4fvh
MCzgVPya4yNzoCv/YjsLW0A/MV09n7Q5Mks3XF2UPVHzE8JarWxtzuTMm5a3dFZdnfsxFSxQ5xYT
M9/EmN9VgzyDPBaG17N9sBurpzVhWpui7jCjGVT9rKqSY+p0RoDLqRIfKfq7s1H/aMtTASpk4cdU
GDV0nFXuCz3hs4r2WXxUe7fUVgawTnvd7ANVPNhYMiHHYHUNC3zN757WgNOqwFYt2iMLfRr0hpVH
cCG9tbETjx6pj5xD3bNUC7AAL9HaWAR7a+UWzB8JHWVyjQuP9cgfBR0UFFbaDgqLKbs9SBffrgIV
O8e9pF96BH4eTq/zhW4Z7pGdYkKcXMOwHyMWiZnLgxWkkjI6hccC0TLPFARjnfsHDfCGbwN/y948
X+TsJo9Kk2S2VKo712zE0DLK6YDIGuC1ImH3ZgrKp/rwjI4xVVvFtxNhnTm9oRKzELlFTZjsK1iE
ZWab4akdkI79QNvX1dUlu3e8jzRiY72zA9MSeajR/vmaxL0QcBTN24YeBCIgwg9YMuuPRaPcSRFd
fv+Icd0G48eQrHt2OUyD0svdzPmEV+Gm93mRT+ab5MEKzhtdLGNNwRGgJmAPCvH2V0+39mA+5R3X
Wc2/VhqBURZnZz9FP18j9hfqIz7/iDdaZI7L7URYhIcPn3RS1OSWP79ZZVwWMFdQylG0dP9ZPhKE
iZOLcWNl1YV3YSxcKDLJzNXyxbcQcQ4Kx8YXlnjvy/AJUnztjnkmVPjTrOyv13lAzYcd2aqEceDH
TsOjo4Dp2qnRbQdvezH7ngRiA7pl4dF3WkZvS2Gbe/LDVlkv8fOhx5up8qjL+CTp9y/jSryZob3E
HbI+6wRQjGDd5Wo5AHulYq9a2OC0xiLVEaUPanGmRqtjU1oIpqDDuDrqwcAnlLgGMrZKPTBZfv9r
+l9dla1VGEPWLJzAvDkORGhgUpdeu3Pxym/TGTCbC0Lr2vB2IRhcjyp1FSOBgz4vauabiEFw3+zS
NgKWBYT3cJ39siFSBE4sEKEi0zhdhptfOEDAWVsR9KxezAHhDr8sBtjRzuC9KM73I8q5+orKUzLk
ezrXA1jmU9ibTpsvgheHwEn7YL8eVaM1YsgsmxUq2FfGXFKwb9w6JM6EV0ByTIcjzxtUNYA7A7Wf
9Jn0KnCgKjcQJUqBlVk/+wAQjZqnO+JBB5ymRFUMqmRfsACtLmACSJzH77feaSBqpyxGXG9nz3XO
KHh5w0XVYc3IayEKYxnXc4X/l6qpZUHZlWeEombFpN+lpJ3E0/b1o6R+AVv96VMjimu32Q+ls7uA
K5MRVjTYVq0UOOGx4EaRsIVI1wUsApEmY025NAtRHqImIQ8a3OnA1CD7OkPv/gCF2qejcGWg9z9P
424qQI7y9sZJDRY5Mh++LseDiUNN8rzeQl3nCccANtbcu9Q3TP55vdp27GbfOovVEDBwWexgeNFF
QKJ0dFBjYf/mGTCO78S4OG8qFdLgjs3gK5VGH3BQg7swbWEgAST0MrkHTiEnHw7Z2r5dB0Sr5WeN
r5//C4Vdu/yeFDOEmBECzpJjo3Q5amwX9faD/BRGl2GwMjHzV56VBeM45qcuVlgxZTUY4nOZiKsd
1HyZDMytW5JE9quo+B+EE35L3k6cmczTAqJLpS5e8Is55r6z6UUFFTiGG1zDK4+7UI3ompDdbylo
p/Yaw+vcD7s1SxGtCcg5IwQOJzUy0LeOzcHGw9jvx63P+23qYA1vO2T/tlHIL1ipO5zJb7ER65cd
Yn8C0z3kMBjhjALhykQuNhL8uKZW0Be3LZfc0AjoWLw0tT3GhXBLQEpd0fPOradVC5E2STrduQjm
eEWXYx9xKkAQsJHwcxlvDKXSnMfoJcdq09ipoCop6dgTtZjyAwpTF9SiZ+s7Fap/jSIarZFYFDfj
3OzRbS8QBUVsi2YEa2duXTf9K1pKYDgEerHPZxqUVCfMztcu06JmQjGAIDolOetdYgw8qtQw+Qca
hZYqihaoozYTMEex1h5m9bQ3LFJw0PLdDgyDOmQnsMhdKpI46BCofFwjBvinYM+IL28uGy6vu5kz
rLThtYJ8wpTxfAdn5X0ovJLxwh0FI8zVjclutaL9J5WYzeKrHKjWzsP4dLnTmTZVzAa+rTroV/IS
QR2k0eSLmHFY6KfMlfg9ZE9hUc7kWWpaah+zCgXy22f9VZVnstRR76BzbW9JTUMjYUeZpvDIVmOW
BHjIIn2iFOJPRfMshCHiSe4Kf+4Qrq98DtjTnDwOhG1OvShaht+SKFq7EazdOrjD/H9JyGCMv7zB
+K1gXwpthV8DYacIDl3jbQpARUiulXTXuTmGd82XH6aXdyGBitO/al9iPyrGT7T/Yc6xjSuRND69
PmIZNM3R7u2O367VP5axhrRv7bZA76Q9oJBEzqYaFUDUtypb8Twq3OBoxHKREeNiIRxxYidFzyUB
bNH2eI24D5G9oM6hUqOvgozmidUgqb8bPE1MhhruotQa2i7D9rRPQY00Tr/1WSnSRUQca/olTnJW
T/7RyC1L7HLHv6GMLof+8P9S78AjI+tVtFnXP/WvBjtJ2utrZ46jjTNc1xptrnhgsDaQCDGMV4Zs
dq/dOyDz7NtjLz21csewzNPF1ZFVqJaanxE/4nwZA69dTS0knBU22nWKHiHrZhATlLzStC/Thzsb
QhJ/HatKJoAVET7nipDgUwz44WWOI1tzUK6khyVJUaEuPEkO2p1OOoFjNh3NzhPrBJUDEXq6EkQg
hMskD+v94cbpe+O7xUWrHLkNf9XzWnnW+s0cjQ+eMScb5wkOFQN08GFamx1emMsG6t4q3KMKiH/L
GITx5/Olx28pbefCX9v9g3sFnxhk9qvpz6y22X71lE+uWePuYJu/ST+atBot59BNbj+Y8Td58pGl
q40mx6dbodcxS/inUt5XmWx1q/oZ+kWGwzYAFi09wR5kSZi3w/cupaKYAXVgpETR74/mbqhgI3jT
Z5K36cEHFfwF5zM6Nh/JTkjaVLxAJ5gFAvZ/hDx+3IJ7LbmsMbx5dobMq/Or0yF8TZOhRJLEJieK
AUmimrLID9l2YX/hpxnv+wKx+e1VYpBvJRMblfDvbXTMyl+CjGa6cfwACYsGzL+18gWKOFDcHMd4
pn3UOqRmHzK4JtfBJkaRUxSGX4+KO0JRX5TCSOdIEjPQj1q4kJ0CFTr6drs7uZ5xanXsxpVKsF54
uYEEPFO/3FkWg5rHkzfm8oJ8awEjR2nE+aZFp8L6DHk7T3mN7OrtuVbmFOw9Ej3gkYB1i7Zh2Md2
A+7D3vDbD3Ioa7WY1LhSeYSTUc5o9SNEzOft84WEIw4HPh8p7SHuRHReejq1gOsCshysSyV2dZog
d3CGQKH+cIBXYqeggMyqu+Hn57L4+U+ni7XUqzzoEOsMC8Pwf6n+e5dUHAuXfo2iLwazIhp1BZNN
+G3zJ188hZ62yE0xNRpiDMtHfeOEMsqXekMw8aENBqw1aXQGfiMuPSSEzwPHqoVsf1FnGWyqfyik
A8K2Qd09bmF5ZcEliq5Ey+MBgcLCuk17Jo90snmo2QgdAwzxVFmT0dYGksTQhr2e5tC2/NKDnO8S
cII+aVSMaZJKMy+gnSnqDQoL9SoBQdxTpWBldjQLM7Tgj7DiMpsR8nFvsVIijIfZxko3taoXSR+m
SDteYYj9Am7fuM3zXOdMRm7fMW5vD4AD7i2/RFQjuTkiGeqg5IIuNOiKDfLCkaTWpjl+wQEx4Vf0
atcc+HRCMTQuVUlcdwmxECe7sUPYGeGYxQZyir8V3UsabRWUQLXYm1/puQE9OOhu2jcDW60wkSNl
I++4inblgPQsr8lopwPX+5S/ZO/V/jZfsJKUaP5AMkynz2jQ+OhusH0Bm5BpiYtpTXA64UXQt7d/
J3JQbMLGhVlgp+05vfDrGV3cp37alRoMlBdEz4JDbxhM3uPCF+p+c4++MCNkrLYRluB3XALCMis7
oNAwlGGc8QPK2CMzFfzotS3I3UZxGjiztx8PkepVHwdPL1kC0mRf8mNICxyB0FS7F9nsPLy/4DYX
tPXzg8fSENZnnaZIpV3wJLy9TSl6Bv6KLtRVyaDe6GTcp4uwdak2V8vIvr77sNUsHvAyXaMWtJoT
Eyg8ljAYGDmPZq4UUPHOx2htCmdyDp6cC1gVjLMdqcyxCjuo+JIgvRm3YNYPAYzArhZBcH3G0ppU
VAx1kSf9AjOuJMwJdeVhEgOLQbIYgd4vClYfWgUXkxvRcnqwKJX/jk8SfbZ6SYH5B+a5dn7mvact
Gmf+Bv886+zJa4Y/f35gFoN2TzltnnHLdUPRVRmo0SOZG9iJuGVQMa6eKzFl+FZ1Y2L7SrmFj+jV
u8EMZRWsrGz9eVRsMsLVzZD0xTc1F+r4r5HQDVXhQkB26u0aB1IUQsvuOe4A5uG4Z8H9eCjJOG5Q
A9ysLR7CGqmFs2fJ8B4kye7QEeDYLObcKtlAxhfQdtxnW3gsU6idXoUH0725MPnn4ekrENnYHIyk
pb82jkR9kG5+xX++6pxo5e5XOEpxugRDs3anBBedRQClXOJ+DHar1tMNHsawkE5Ww5CffIsptM9D
gtSpY1PVmWs6mruKuouXsO7OOofBu1eZIpXJ5685HV9mWI430HPcfRuhMhB6nVP3aZZllYo4xPxc
8XnXgQihVZSaF6Z3OrL5xnd1DXoPw1LALeVxRBIDKxVRew8Qjtnyvs52QLR1Oj+U5/A6qhMVCqdY
BwPtDlo+89cjXXJTLM48UayqKMcwL2/8V8wmlDbgPIEg3tAqjlGuqh83y/hizsBTdwM/f8MV0DWN
XHT3vAhv2U8oON3Th4/B8L0U8YOLCM9udOracDLDTDmnVOXJbHN7aLDTANlLMmlizKqf+DtU8TGp
ahVL+bJQ1eK8d18o4gnu03sKMMEc059IhQb8OmhPfFMrJFckrjCvWkP5uBj8NeLwqW0S7+YZ9T8m
QX7ZgqLVU35ZJJcOnSZt/y5svFV2BVmYgoVch+OgwQM2Odyh51T+1Mf4w5lkQWca1WSqozRWqxY8
wxAtDgB40uabx7mB9mierlUMrYUQyTJuIbNtt1MSWICNJZvRmyVXl3uQwYBHTNi+uUtgpq6F9bbx
8bmp24JQ18a2FsbuOKDwQqa3VgFuc2wRR3/6/trSyjQ0RRdWXpae/QBLEoMYzvlQYC/RqzQoYJET
HxlNyhbTuHUsjnV/PfCRWfPvVwxkcxl0PH8QMZJwArwBYo94uvFVVNv3aPi1qGquDcBpJyqm+x1L
HrrQZozWli834Muel6TZYr+MK+Lwy+zQt+2jiSgDCFQ3W3R/pn9L26fJC2YPqw26Ry2aago6t1ZX
cgb06AayK0T6+Ck9xaPyZf9RXd/9h/Y8vq2ftK8keN2MwOoftJjJv4S5HONcrd14tp++t5O5nUQO
QX+ej3YO1FZrLTNdv2HGG4NelN2v8dCZ1VCk9qbb+nCThDdM3uDoHczdoAbXU/GvR8nlL/u1dh9A
iixZ6IGFWg+2RbJ3mpU/Pn1frUKpDlScyHFyi/vqDB+U9+0k5lPYomaSnXwPvoC7kPfmPTdYkXAE
98vLVe68jGynqdlMODOyS7cGw+ufwPdvRurjhpY0wZFsEn1uhRTj7bCod2Y4Eg+YooR4Vwmh8ov+
KjCqyHyZhl1BHKXTqnLusPf6u2BTjE4OPYyhn7DSaELUhw8FQVCith88Gpp0j3ogYHzcmZHlb/5G
i1nOlzyQX+CN4amFAtaaOzn4J0Fg4t3ca9xgbUcR8Hy8dElKwkwhOfFgf5oIHO8eQm83LfLeGbsq
HLyk82g72qHz9k0CJuumm2jB0CDUlO0kSbymEXPiulV9y2bsIA4S/SXb6x8eHjVJPjyeJ9ASWjoz
P5UbkJNncXqSnICoIeak6RMxVBMJojO49UUN9Ocia8+VcbdwvcM5tlMdJ9Mjb7vLjAbMWDBrHyjA
ET9IIJsMsQyruELFksmPTlD5/DT8aCsJDwLrI8EQn8Q9Pz3ddGskF3U6IMMYYDhVjAjR+NDLHXlo
BzDtzNevBh4BrCCIPPARV3GnOH9pxTzB/ROIyRdPiKlko1sN/aF1KnUjYmrzxlZ1x79pSMtKuANo
1FJ0x+27owq6rdtIw3bnLtOX2kDpvWaLe3uFQLv6WwEVgj9XBT8s9tF2mVOrRnOy+tCAsdisbsN0
HLmV2F3NCdy3CIHA9oekrC6S+JNNgtZs2rIFhsZxyH38TW0m6OG/WLsUWOwy0vBwccDnuZT2k+OY
GUgAZjt93WxpJz+rOQI9mjmyTU9NbaaRXdu9d02s950dDO/s210pvpXbQAJHiBTZkl0K0Tfp7g6M
8+1NYbF8jTbpsb7QPRtNP/RwKej7VWx/jhQH2SkBBiCDMQlcjPaarhKISrWe3xIWeSWhRgQRMhuB
FzUQZW6R7EpNWXys3PMHI2y0vYTfgMk21nsXWDRQmeQ/n+88PrvUUK6fhFqF3z1Mv5yvRRLJJgo6
UbDzptzS3WBDituNJr97jd/o3SyN7RKwE+DrXS60xjIEuOpKn09eJSZCgDkQU/rWlurf1ANWgccM
z+30ArgGUAJNNZ6/kZH34J2HZVDYwULcLTjM+z0jWMsS5ieERCqvcEpPxcZjkm9yf979rV/vZZwT
RNRmhTgk51VwizxWzc1pH3gb1QJxr/BTenkrAaix1J7EPWAsofRuElS1afUDm75/+06ZQlaPMpmV
xlyeDxg4hrl3f8ewFtOtO9a3vRNn1uoU8lFqXjDc5OqAy6nb6WsN5PGFbvYmtl0LkE8R8ruJewKT
1+NSLMOcpo2xdGyl0ja3gXi+uXW3V4lhyCzR2iPXRIv1Uny9Ug/qj8vF0QnVMh1NjAAeffZlaW8R
Zs+SP+b8qs/Nwx5s6lh6li+/q2Qwk3U6Tv/zHxo3YuvaZewOxMVaN9lNccH3kph5Rh1JN8u4golh
IEXnQJeLXyJXQiTKUjPvh9WBSIL6sdQcCk3RmqS1g2IHjVMp5YWF+KK4FIHnEU783zegatja4cV8
bgvgNO94o7sGxcYSkhOVSCb19FzQTRyHMIszqOvH2E9erIZ2aYoLwiF5GRKJ+v0Wy+pAUiqvX34a
woHQN2IfwcGEF4fjyhf7c20GylzAIh6Psa7y1IBNiz3lVDRPEFYhsqNYWEB0aI5gV3oxGuXIEAnE
/6+HDWAv2zBnR8M0DwW3mn9gitRQjv9IDZ0AVEOekV34Hsxzul2ZNu8QGlDtH9WMd1RPVcjxNISe
53QEAfWBIRprJbAZp+ZxsiqrW9B07sV1t0SVvj3obB1TZE0f+JausnqahvvpclFdwDISuNdLX2i3
Ch9Ac+UXX8uVwv5wPEhv7CK9sG54xuyLi+h5ZyVwV5OiqyMyZG380DhNwC5hzdRzXzpFsTMMFGFU
HNFYfOW3NWePQNbTjsXnPvNnwXEdis+JN34yUuuhTfav+IaIMpuntDpI3/i4fFlA2OMeIuyHikKZ
v/Ayqx6Mdw+PVQ8+nluCt7bK9L+aUbmUq+xZ8xQdiwVHcTWp9w6oe5SrXZ2BAT0LKDUxkmoLdprJ
pZ41Ox4qJisJIsAjJaC4j8coBM3hCLuGm6akj1I4+0y6OTjskowxCl3tXi6s8iYVCb3a2Tog2AHG
TXkVWR4Di9RLIMakwtyZEFxIAVEM5vSvDwnZYenrPgIZTePPfCdHHL5PoWDHRZpo9Vhp5uR8t1O+
rGLqaaNXfOv2p0C+KaaH6s0kIfGkHUAbuQsoQ8CvUNF/H//FmylrNJvbz+vxgHHGHKGJpw3YQdzn
MxoSbr1FlBa0CHOk3eLS6tej6C3Wahhdk627gUcBCfynq9atsRXFHsbkWF/5Oiqg3cUhVOKtXHp3
qAfVSJ7gN71KSg9zgvJtTUJOie5O5qnTQC50LTA00FwWJmxmgSNNFzjUfDzDuN2G8HCVHedCHcTx
OYreJltrc/6YywpQErfRSuDsBT6m7apeWsa25FsIpUTsYc5Ra3z5b6USNPiAbVqwIc2TUQrrp2au
45fezbKdDRbKauKgIznrJaxXOT5HI2vFbXi7XCDur0fvCA9gtDy4K8XUoLOASs/iqTwoGNJhvDZ3
k+evj5i/cESPbnKQ1nhcsQIPTqENTV4tao8NrrzxZ2MswO97Jhv4I1qoEg0caNNk6ZT+jBMtLa9g
+9Nne8aT0ta39j+eNt/e3/I2FIRh84bMzgaF504b/7xVnkF/Ps7qLGIaN4yRFpahcSNItaCGSlkb
2f3mf3a1VWCV1TNTePF5Q17rl8+uifCycj7P5vUG/StXLuTE88Xa6pCDBEVqTpyCIFveMa/6qU8z
ZZ9gEoDXlDxyZXY1WjT2ZdrmEC+bylUy0QIll0HK/HqhUL+IkicxvTdfJ4R+aVDQfhJLUSGr7wKV
EdA+TBg8x2te4SxasyQq6aT2UJA9JZ1fwiT+RW/j/fCZofe9gMC8AXdIJcszJEYVNgW+eiPeHTHv
lto7Sgyt0nCmduc+mAqRfyrxpr75oFm27q+vLii/E92ckxkibnXRYl+g1AIIIGdDlULgHb5g5YLV
1vErlmV/HyM16aHUIFUhHop9CrxpTBGCcPP6yLz8lX/RpFUdetwwdoEtJyBzBorCcbgBwIunQKjs
3esel6hz7rgJL1fg5UzAgfli8j1R3UsYSMGj0zETZ2CBEE8B+vV2HmpU+utr+kbtZaX6maqeoCSX
0u2nfG+TE5q8mgJP33sJ0Qj6IEq37abNZYx3PbwZP+eMYIBHNxEoY2GOv1KwY+uf9a47JcofGc1P
HUq+CCKCgwN9XeCljeVueUoahm2ugL308Hr+uryDGO7mcd1CLfjxtoIHrQLhmAmKHyUcEcr936SH
8NMnUo3Q8pjwIcadsflSdyEjOztQUzQOg8kqUZu70l28TxVpF0tsUr+2DyTUyjICb4o4cNx4O+vg
kzriEuK4iXiDdTpjywd3btbECQvsJVxTb+osK0sZaNnOh/nHfXhOvKciqW5XzMiLnL4JYzQH306e
YzjkPFYK6Rc1UzBMSycLQ8kHN1roQnBMzAuI/LrCmOUN1grW16XSSp89SaM8E6wuYINPKo///fnS
APp9bsTp5QzyJ1vs+sjUghmzfGhHn7b+nmUjhZjIbLBBt0k0p1wEVALl32KCfARXcqDY4e28fY1q
C0k8aF4zHVgTR9PrngIheXuj8x16gNj3RbtOJmrWZ2dQtQxzYsU+KwsU3u3l1KIcz0S/6UcLJCP9
yesgWdDH0uYGi2xCq5B6QWLTxzcQEM73nYiDKpnKD1EGgWMgxLdBuATOjeBrtTuSes53/aHuQwd3
6N8vIxiq/e90CzocZYJhprdv0yZ0w7J7iPO3nan/apKm/1qAhAUGgeWWZgjxmSjo8f+J2UZPPgwZ
1Hsh7gJp3UOqsWL67C4ZSBxPt9ke7fuIiKKgapKXtE69tYOV8V0xDhYC2xpMDrnBp9SNpuhOc3SS
rfVxbD7hMr0dtXkWRWI01CYEfC/udDTS57lTMSAyZBqkqmzvHFUU+swWDQB1X2fJn0YnKUEpOsjf
p41VFi/jTmkikGwcryypGWj+auafoe9NjpEfgwL7WBcHoQpu9Cl6Kuc4UyfUeYw/mG0kAuX0mLoY
dSC3oRb5HkCgpc4Hzum0AUFCKBv/T5eGPNck4gA24FTSS8uuB8tPnJ6VZfngyvJoYvyd3ms9Dj5A
03t99DZXCwL709SUB8QFdN8fVQTLglYmTItX+IndeHpIC6eIqifKD1qSGLs5SHP5hs80rdQia5jv
gRdi3694kRG7gGbwkDqlevsDXviSGrJlK+9gtqhRx9AOKUso9o7c2N4qiFWjUkfCG9N4QS8tlPCw
y8Sbxqk1CTEoZXGhVIRpTFsgqU7tit4CPMUxS2qa5vetr0TtVIe0LR5MYpOU1ed99GazVPjDjipk
+4XwP/3J6SgpFRAFc9dAQU1Zt8hmAKj/KGeRYb6xBFHLC2u4Fyy49X4Oz1vYyW2VZ393Mly174qG
tXM4/R4bTgZ9PEch9VHsG4GoNNHZ70nDxkDauXTWA50nVGUBxOP6aVDM4kmtZhAjrjhpzbrdMNyG
xYDOrBhbZ0hNzC44kxQS4sr1xiySpPgH+m8imfLn+rI8yxIZGQSV8/BdSDKfY1g6sdSRkcyklKpc
LszJ+YXGTo1JFNdlO4RWT0JL8sqShxhbAp4hII/dXMOdyuH0cnwDD8APwTefr02Ka5dZXAnHPbOs
/gO/eZXk+c7Hni/44mpfEE9ZiIghuE4AZK0Z3Ff3qmQDlNvH+Ba8lnfME1iP7ISsUCon116Jo9G5
s7UXFWJ4jK7W1tcYS367l/vd7J7X5JULh0oS6TbiFchfI7x3OL0+1dduKcU/J4w02wigByTuis8P
w/3BQxF3+IFA6cFCGM2vsEoXTBBqbTGt64U2ifJb0dE3AulP/FMTis8w5bdnWNpJW4QHGdNGoavE
zV9qkpHba0bxJTKgWiJqZ/kJ52OqSkqW9tJr4aH7OzgrCZY7st/YrQ24dy/J0I1LKiQQgPvfZIdp
ZcjECNE+8u1hY0uE79llEtBHncyob47PSVmRtTVw6q7VoXZZKivsPgYXxahqBG4E5cThsVfhE3K/
WDcYSfxwwMQFGZ+iYas5B4xD064VhEaK97m3692UzCNHdElofYBN8iIz82U5OJidEDfKniW1SKwX
KcrlxuEPfE6IxfajCd1q4GN/8A6nkQBzVQQx37SVA2CTgBW1Ft7g4XNbbUbiyo34OZXIHVUFd+R/
dT4xug9arZg2JgwkPWw3OSruhBjapagYLZFS3JC9KU2JzOoLgXDtCM6XWnO5o9HsFDxgVddIxgVO
Hntzw1dvry8GvRzv+Tzw4i4AzQKF7VCWNE1TThCntQVizRtVqt2pHAO1EojJNGkrahYE1FCKklAy
wfHfl4mNKGhJ8uEKfRNKYHswmkv2mm/Zd/zcVpHbLDPNnEbHta9ra/d03dkThKBqSDXs9fSgY31i
cEgoK121IJSWj/nVm91S3gkIb8Lq9GY/6WFlt82ZbC496sqSqogEi6cq5YSeMynd7xEFHwhHgQEe
gMZ8LqHq/SID9e3Zc2NUgMZjduX3f2mEwjfkXqZ9KCtKrM0l2fkqLoeW7lrDrFRDl2/iIzv4WvPo
goxrgqIQcwbtv3vn+uRkYX1rEG6OuqJCK9eIsPhOfJSU10nUHI2FQqtZUqEiFZWrsvhRAPq7WCar
jHCiXOkwbHXNBWbeAxWeviV56TGgolJNAB6bz7Z+nI/aK6to8EisqgTiHEc3z0drnUfLruJXFTmM
kyY5nJHVZabZ1Fz0c5+BLRXOcQD8mcj2JbnU+E3gg44P1kRHLCTSv7+rfzBRjesh5b467EP5eLAH
b4W1eT3Va31hoiHdfYFNz5pbQnAYANDgji+7brF1VdzFan2d8qKXAxNeai+QiCiUCuSol+oOj2IB
rJz6MM1t7I/BEtPkt8ebjxBm0CaQlSIG3xOWTSmXRSNjXQGv+G7LzGgz5WAt8jCqZVf5rub6Jprk
94pgYbVs09EP2KEovoXonaJHC/a2HpMN/LwFeXrePaTn20k6ZOg/p2MeRXW2J9SEQMw4ak+YYM/E
vRK1YzpAzGgNbZyzUNsh/VvR3QC5BYb+TDYXfRhLrvaWC1pm4oM9Gh4DclbIwkTSqXxaDAqre5Hb
Nj0dvJCMzbkLvB5JUEvSBmQgovSYs2BAZdoDa0X1TwKWoSWlSLV3n+SYH1ech7b+tVcPgLKuQUTf
WelYXS3t6oKad6SZcW8OPfFiRw4Ftojg1tWODg7Y8U8Dk2IanqLb6rFdMR+xwPlIA1wWbqgw3rjt
Qrdw/oQawvFzZ2rCQkJBHlfdvOGlqDzo3RGQrFiYSBnOvaaIAb+f3Vf4BSEJkWPZ5o9dY/K/jYXj
CaRJzMqLMFZ0Bdpq9aCpm+CBP0qlhL488QHCJx4OfTeLVQfzeDsALBATMQ4pb0Q8Bg/qG5/HUg4S
t8jsMiz8MklBunsp+dzwKaFbIdVKknEUYhCZ/0y/T24tIhM485RWOGkE2qnb1OAiie42DCS/2n8w
DH5k6k61nov7KrYBARI3p8jVIIEy9WRGYfSYqd/9y5CRqKd0nIxUmU4kfRVy+1gnupDdg4CuY7oE
ZzYEzDZ75Nw7uVtnLn0eIXZNoiDwzmQ0SjdXrEtSBYxrXxG0oej/y/RONex5KoqJqv/vVswhckd7
e8tjKwm8OfWPcd84l4aSIEN/t6vA77oMyTH6JP9DXMyHmd3UYweHdI4ffKcbRIStiv8ZG5m+5fuE
J0eK03j6g8pqUsdBuRGytV6kURubQXqNHuLjjQsvIXP9Rh7eF1G4Qa70wkfOSpVbeZMln5nJUd7E
/xQx1A32aRY9+EbU4gJBRkvaVxW2b6rzpIg1BXb+PoqhH6N6LqPwlQ+ESJRXSo6JQmtSBun+qGfh
GxAfAy3v7hD8HamD+ISm9BfCX925EhlV2baZArwgsjT69QTZksSPAFvu6dmueUWCcZMopvYBvetC
DRRRgjfdTwNq8TqbYHUiryxu1kQdTphBQTeSSNhjVD5OtQ/cx29sylMpAgJPZFE3xR0yBxrvuwM/
aAtc/k8gXEDiUeviWs5FPmcdbXRAEhhIP4pVn3CkFppkPbdENMiemCtGyhZA06HiIQl7TXMZaHNa
7NMD/zMgL2FCdVsJpsow+Ea3UepP51wulsqA8fGjFI2u6P7jqNS9KtRJWXA+peiAj6jOaZt/j2Aq
tTvTQQwWXWwqKkylXkefOjpLZXI3wGZ/njloeE3MSo6l9QTp/0fFZPt6srx7kwkljDS8pN3TgMHo
mKq5ByTcFJDD4Z4lTUqmaITpr+9nk9/HLpoEncFMq6kYhPy+jvVbSQ97O7VR6A6YANXb3RB/p1oG
d+Dj1mbCqCpbpa5FNjxTl4qrl225dwVhPMSG8kvjlLkCmgkGDWvpm3IWofSqzi13TaKztCBgoAA5
l+N6y1lJW3nK4j2mt+fZSHocbaRNAw+KGlTcjgigN2Q028eyit+pWEsY3ujfS+fNDYNREu1DZ7wv
Q1e+F0DE9jbs0FYsKMwQnS/2udxNgHROcYlmeULlUcpzkeGoOZpXMqPZYyNTAW+hBmjFM59RyPzG
lfDPy2/YmdNs/W/iusyz3GO06jDIl2i/zjprSFrvoFQA0imG/dG0FPHMRILVNqCRUosYVuDqsk8A
9X3gP/8+efjjzFv58rFIulcMDyw8ABS7FsQNzWgRZck7gAXjBH7+D6GKf0SFpZlMbs4QUyZuASo6
RxLr89q1wdck9SfUd5Yl6dQ7m1BkyHEek8XIvw8+nnUj9Z94xLvSz0zjEx5SlxgIBYF4UIDHLdRd
swDMKrZCDUFmmPDCJSYSV48xuHPrx/EtHi5JDRKVgAAzYMAuinJnMAoDcGpZsgjFm/hjhE9ho3NH
ZaPMN2BUXNdg/aeT0OWLPFLcTgwdu9nb0vxJCzhH+rg6uXn8eio0bjdNic1qttgy/gciHpTue3f+
9uQzeRqzvEu5NN9qw0dGIH2i2EuNwUzcuAHaXntxkOF+mnoT8N3u05i6z0WBL9+FSvYnuQYEQJxz
9g0M/bE0xrwY9p32Tgodi7gqj/ikKPNenfTw+pYFDb5eO6dNKSJbfHfh/vbsUUzmnkBg40axoF2h
nPJuL55l9VJ2h6mfIQBGWJfL1jlID4fS79XDF9HOlaFTMbxNT8A88MFvH6+09Sbf2csHQeEE0dAE
zDVZyjjl+B5kgLiZfQtJEf1QZ0+vhce2InRYOcDcFR67bftZ+ipJmUjytO18U5D6BoP/Xe+PzKCz
xig6ZcYCcpkW9mAA48BY38sZ6Y+QCoaRs8LQ0glbgGmMKI7xkfcWFxDdOIBqIg63AzRjocrCqeF9
u9O8gQwQMXR+n5NdDbGBZvFp0SYu9IODG9Yuu9HwIOGv9YRv/z4x5N50WE2SCsKGqxp+QFzKkJ7a
daoKZbpennQhUBqrE/DhDfqk0PJLgbW9dbH1xBAd2h6CLRuTLP28WNBVzIPuDhyaXKC7kJtXNfPt
tCDyl0Ecu9SlIg1Ky/y5aAGD4Bvu9bHs+JJT2OJ3lXrSfUsXefAwLZAxRkuh2XOh0RoflkIrNYID
ohPyEW7Zs32eZz5MgcVQNZEOJkseG2Erge78+/kBVgmtSH+UbqqZo2mIVzOQ7ClG2z/UkGS26OhQ
g8Bge+kmengWE/Fzl3OEVp2V7aGvn1J+4tHyg3h+dVxDvz2+VmMc4HAlphFju82Sw1ovfKOZn9/g
7idXXxyfMc1fg2pQKq2UNShYSPzAvACV6LA4B7AprrjaJKYn1SHblkK7xKZ/oCDJY8lIZzjjfeWq
ryvAIfnUmM3yRpxVUr24o6zfJztlnYszYuDD7BOIC8nfxQVclWGnKVUd0x38X6y/Jkhat0LSVXva
NfeG2dde16DlSceHVXo9Rm4wgB+HSzo+lQmwPf5MgBaJ1MA78z/Pi29tIZ7JB2XWkeTaKL13K/eK
Fh8vI3LXuj3YILiam60xvYaUNpQm0F39atdA5s/rtfJ2uUvK98buMHMevUROY0yMWF4KDtA2fUFl
XM5IgE3MVLWa6vviAxTvjw2xipalhAWZJLJetrkFLWZttYxE3jIoYy1mIuyeqb2t2ClRYUqkbyhJ
IHLisyR2gw2xTpaCYQmDNdO5PCmYwD+vTsSjiE6zois0oy6UDGeVXF6Iu7mjeVK2nAyxVzmHcwSC
QS7kDXNUrmXhfNnzxxzWOCAGdiGDC8th9BnIFho5qACvSk9XUDjGYmpkBlPRX+7D/O4d8mlMKjx/
5R+mqBHjC8hEp5pi2p0gee+/KrJFcJL38r5tWXJ1s9DPhO0JirNTOzJ2XBuNDpj5rOAAAwNvkJuM
B5/mqkKmEn2rc1/xwoYIA4VCAXlaqUbjqzzw6SgKHiPlGKNKcqnCFAOoCbYWXAj1Cp5dA4TgfxtS
9laR0ekzM4gVDC/dAVBwu53UbOJ/ZEOr03TVPZ3ji/X/fko/r49ZPYPVXSdY+yb3hr3R+R3M27gE
wPrZt5pZY+gzZOAD9fMGvytERoXyC8KI1ixQ+FKxi2d7umBM5v40G3VxPabAhPq92h3B7H9vH4GQ
QV5bTPWwerTUmune7FdBZC4Kn6bbVK4V28AejRK+hUgiHhH1qmvo5X7HdSn/1eQdgO+7yfGdhMR9
EAVGus8fKtj96tpC00MJHaPkSLnHvseT9Gy6gxRDdf4RDx3/2wTl26x3CGRItZXmGKFD5fiZMHmj
8z3QDjeiYu/Jeo+BXeg+Pq6fvgh7sveqZJjnDbS/3qPpI9u5jnZHuG+RryTmLXLwJgxpSs2IiGHn
DbHKjsLicDvbk5KZBDmV1EtSLpTNmYarW83LLdjffplyUhBa+CfE0m+dxB8QrsOnL0rW0gfG3m8E
1RkDPBDBpvBAHEsfheJndNrBNJ/+ZZGg9xn3GH1tGrfa56caa68bFcPSWNMimnDzdNJhX4DPJ67C
AbPivQoVyHyXAUp/lxyzLDA165yeMDoZ5iAGe6Pb5AvdvyTWs6RBh542AFbErNo8pS8VV3tOJgSP
dzVGvqe47Z0lqCwQP/BjQIsat49zri0bABAZCMMqIDcjje4hltOgnqGQC0zfu4HZyQqwEshBjZBE
7zdxHqSIDHdhT9XqbtAytob136e0HXelEOx0vnSRYSUaifO56RhiK4hCzZ1HVlXAXHLlolm0xVBs
E1fWDrKf26UFdHnMFGdWcsj/MCrg0oOzaHilnamVHuw8cNNRkzeYkK3wnDafWqZSPRxQBL2pSs1c
iOqYPhOjpRrfeZxACmyI0QO1IJgj9ttaX8+kSJDGEGsEkwjBBX4wNvjtNZgMlTbVaNCWFf7AtCOM
mjcxQAgnFqOOanga46Nzn3OpAi48m/9H88R4fG6ZTDbUuDcAnEY2hKby5Z2YbXN3y/ETAjSjWDF2
8QYyl/A9ugNH5fNowD7kRWfmUo7z10Rjl64r3RsjNF0is8OHqkJZiRh/ppPWCiVQ5FTEC059F1kp
PVuoFc0GVS5cufcK24lc9K/GE6N+/Kwh4IRTUTlx2rE++IAizZV1Ovw6V+uMEmFHFytVnLV5hEA4
Kf5I1/Gwmtbmpx6FbDZRBDhG9TTktCIMzENZr05zMZhm1gZfaVjb1QGq1zsyAzsVoCikEBIMSvAY
rf06EQJk3Qwj/s0dDOLNDgdPFmGBgRETGn/+JeOhc+RDmqwtgdM+a5Tfu5213Ht5jLtvO2WutYFm
OOj0yVW5vYDax572KseNen6QgHS1L445BdDfKWZlF21fK6YpMs6YGh5WTbEcr+9lirxkhQ9ybDUP
6pAbwzpF3xlGgC/elNUzx5bIP5ctmNj0h9W43dd7Gmk0tKlhlaH3QAKd547XKcjpBB3+tCBXDjVK
4ksBmBFbBybE3OYE15nvIp8to90T30x/m9shYp+wa8QJNoUCotwSE9lR/6K4k6k7c/R107sBdeQo
+S/+MnEin+LdwBHmc9EqVWaJzb5WTrE1nE8ey2H5DbfdV92yU5yR3zfax+CEOMjej8H+8Z68hDfm
ZGikBr982wyZibSUCNk+i8koLd+zZE/xl20w4Tr498Q97ld+SIp1WPOh3CX4pJD4AQPWhcSCqsXF
1E82J5xX57KPzHZ2JXyoxSGSoeLB7fgt7q0pfblBtMRwz4hH5r2ptghzGjvWC8TttItF/lTjIRWv
Nd0FJ775RP36+E2/wsirJ9v36rsqKzszuLHKOt08T8QXpxVvpczh7dutSj8Q3lON3qzCIQcOZHpU
0Dk1eJ8bluwB1QLL9PXoFAvpk91lFIeB7wcqLPc/8a5IOUzfWtcHVaU+uRkmqLaQeIgt/hdG+9wE
Cu/BsoWicJ/GbfeAlttpWaKFyhFGV6+8cVDn1mp6oaF7FFjoTl0oiIQyu+jnp1xoWWAKa86ghA/d
s1ZlyWWj0wn845DWhDLJlrtZC98p6rrCjTwMAoLdXRIXUG/yaeNpxF2sAbghOScwf46m9O0MpE+d
5GNNmRlWNlTM4p17caF69RVwkx+THeJLgTGXjjvQFqO5HYEGg5qvbjEq6JVz9s+tnBzn7eUfmR2g
9WKp6D46T9aopQcrR+L3hHRiLTm8ra09WAeL3Ofv8s6zuXph4LUWlS8agFHqTkPFSrWRZHzy2Yu1
ffYQ+w1ccitzhOBqGWaSkcKZfbvC6G7M6CFwk0hyVPAGtVVrhkgETPuYNwEbPLZYf6zsfzz3uxWY
Sm/oNc/6e0d2hli2gl+iZPEF5ISHvGjLKC2oFNQ7VQ3gs8qdBZ2pSKHWQp/+l5uVtQuaEH+KJN+6
sSa+qf3sTSyWoI8bfl5QOKT4EZhXdvWlI44zMkZRUvtdhL9/uLxNLn3dINcOgZb0pxohML3UYpgt
k3Iy0e3l/4LpgVpCQFVYOnf7zCvmOJBDAjgtfZFUfOBY023ycum6f8HE57LQ9YPyBST7jBi4+0ug
e4ajOMtlj6PfWPXsntcdK+Fn5+z5dlnRBs7VK3qlutTsegIhmKngkdkB9ctOhAjy4J5KZYib+dau
iz9wxhN67hgdR1jW1pzlaQNQdjKoUrSgK6bROct5XduHAGbEwQLjOvilFIx5SO89q3P3311H2pw3
Z9CvmNBnA425gdHB7dlGAze6d3IkIdY/dAz8KsGreg6DWydRbVuMEbDxwKMoy1478tOAg1wICdL8
NR4Zd9gBTvf9/ZzZWx83CEJ2EvKkyytc49vY4Ze+5p/zo34pXxHaalj9TlGXKa32HJzT4USF7GrB
Nlpj5YAe4Uo6Q1QZPKC/S0LnQDZmFnLMMfoI8+XlSeNioBTxAlIrAZwqeEn9J9S99PSjj4PaI2yy
Jv9jnYjc4QkavO+BrJMfIdPe8KQxE4CndOALBfs9+UntF8E8aH6igUfjmU7OvopBKT5WltelwGy9
F/0BLirjQJIEOHcOovXY8TISxNkORNDf+7K7JfBEIfKngb/Y8sIOegsbSJ7seRhGMPFwC+m2ZdAg
DJ4N75y/gI0OSNOCWQUMs2FfA5uYBzPqzD8HSsvhR4/xG/XZN3AKMF+Xut5Anai9jw+zeQ5GaTfx
A09jT7UmuP5SaOlBqRl50z3VRBfUCEtRSXTndgaUKGSgaM+bEeMAfh72s567osk7Dd5OVpw3c5bh
PnIM2RjROOwPfUdU3s7HWC1FwfAJmUUj+YAOiki+mpzylLpgRCdigOmJ1D4UCQO4BTKYLZwqzEnx
+ucRP8qAIYyddzqIoMKd8v/2WdzrTcUvWXLkF/HCZNP44DzK5+qDQQhNk8fT/CjVPpvMKsyQJ3ii
zIKWAbEfaxqDj+oZDb3Oh2+vRm8OG8+qF+50P+xbMpyLlcyRYXEXGI+hmvziI91ewMztWnSnSyMl
R8aAHlfHAWE6W9fyy13UYBgQO6MlWid52efdTTvIxckCpE/8I81ZhOKf+fX/t3A1i35Xr6yHh3/R
7iptjKH6bZEVKY9mexZKfnxDT/1YPabxIZX0kc0q5ud9gPNlz47La8IcftwrkjX+aRHjzbxoKoCb
RpR5rqrkxMGmFfhX9jA+eEmMMW/tr1wjIz+RiDru/6xQWXa9iXVIvten5u+hFMcKDz1WHZmtyD+S
qJZgAmdqQeBxRq2CpPpTdWh+nJVAqKiRWm00Wqcx6AAZkuKY1bzt4huVJetpu4mbk6XkSFw4GgXz
9eqxJCUkxV4qvQjo03dtZdm50GSKeXGhnBHfnFl1DjM2+w0c9QkzAJgCBbq9qeEkmAAoS6kv1juZ
Ezi4jATKJdovvjuEqMLtsfOzKQa59OKyF2nwPI7SUnZNY5OOdT//Kme9Dl6k/E9OZD/tB6ml1lvt
m17yp8a75NcAIFejoFgDOTZ2AbhDwfdQa3gk6Ic8BgE4DmUHEHlLaHaFhTLImpHFPf3W/1FZuRks
za2OpCYRlGFrNvGgXQw79Y/KaCeCrrCgbb0A6nQhvLIfULvB5tC7VdsPkSGxx3RCfy/ET64+WDDx
614+kMkGO6MLMxZH9RsxMgqCKFL8zdmEINZSceNyNrmF3ETJt8dSzaeNsFRR6n/kyxEnPiC3Ni1E
6PK3RC5c0VJcIvpXMxckFds9pxDI/dCRNNjmgRQSMmXG0BwMGKxxyCeNYYXUR/tlRLtYV4xaw1c8
1OIJy6H+ip3kewO/azOoeLiUFhPPk4NejizQ+yap+g1hdZk9IPccHzdbXNReE5mJF0TBCNrjdHWn
nGKJUTpD54rCxJNJwgb1K/Yo6aAKR81RRWwF4g+nEEyIuQm9wiovmhFYoZ5TBKPQkgSS9bxEEkIa
lHQKzGNprYFoneEk5L+MQX4/eOfXF1FzbaPcVeZfGOFWk7F5rUwrHViZKbiCeJdruDx+6fXIZhs/
g6fsI4/JYWDUmFlKGGfeDP6SsZSwP58aCWC1M+25nfqJVu9SW3owGWCYwL+clynTZ7IP7x/wQZdZ
GcLFoUHj1h/aM4RbdCoxMpS/TzSYj0k2BGmMrKvKErm8IEgxH7/QTEmxDoLgZzdWsgqfDTBEzuum
HfGX+7IJYOJkvUuYSs4SpYn8STRrgK1IIjCcRrTMQY0zXkB+7pYzj4Y12Fi9WNWrtYWDbbXHxHrS
q8uFZZjUdxIbgzwreFTyCHlVMT+JoaXW+aGZWYRN+fwNBcqKW3K4IIz6XOg0AB45CKvTGJ9bTHvz
XqaB/7cuYqATtzQflqputIytbVbWF4t0mEQV45UG1VHwBiE6WKdizjvFiwR+3VGt/8+p99SDT2ij
gKyCDdqvSjXi7LLadcnhucQR/TS7NAPInYYAz7aHQcz3T12eNyJpBmn6g0Hu6RCcyy+hYfQEhp3h
aTljbXV/Ac+AWDIELdtdaOwMY/4cuwnRUzACgbiQGYjwLGlsNwc3UDDSUNlFwraZ5uALhkg9+ZUP
PXxw8ZEmsMCS9NcHuR3wKZGf2M2V4KFZimVkkdRPDit7FicfWasEucaMluMF5bjAfLJupSKkpgEH
ZHc6ehBYPoa9a8hbUm90HVUCSzOcSJ875AgTPTSv8NBX8ngtKyedK20vvQElWdhR9+pRzoKlGgn3
crTKIPlUwJRWybmSs11PxqtMCTs2bXShtVOAHKeKvwgz7DoA7r9O9iD/2MQd0OL2DDeZOiSYXyIg
aRbkiGe+zvCkreQDhnrOmi1HjpvUQcBZTK58PPNpMfyvn4oXmCa/ETyjAOW6DIWwnb+lVAyByraV
RzjqIbGiUrbS5V6z8ifrwkH/mUgyQq1UkRnzPQuVrNU05Da+WYY88Zb0ClNtRDzT7bpt7CiOvExh
Ig06do/I/oqG/ozwQ7V/NcH2V73Sr1Py/ig6egdR8ym8wjio50SBgkixcQInjwVEKt4ydLiTmX/G
DIstWxnGKKeO5XqG3LfpRpC52r4CT45NHFFwAIaYmzuJL/YIBwZLCLbyAs5AiLwtZFd6divYZiTb
j7Dm20l/Suk6kiX+P6jTVYSuCHrAC9qPn93Mc8lGWtjPxtG7zHplLa2zaY03uj6hM4RQ/I6jFX/A
KoTAUIMgpm2k0TR3QGS0NaS5/yP8geFOwckui6BO3X/gPNuS1JgOz4ihOfzuTd09bCHOPt6jS/1x
tWSMRIpxsBOYD59t6gidFMhdc/VnYw92TS/nePq+rDcuWqTsuq0ZbB/xVy30VCROChs9LrYlZ3LB
LZNsZlDNsIhR/aSU+OIQu2yFWZYbz70moVy/p9UDCn7w3ZNCJTjFLAF607/Gj6qsdv3DBSoi/08H
DFM0Eu7Wvmg0+Exn4SePpRKeY1f7PlC8RKOKCXUlCDCvpv006FMbmO6n/UVdz3R87lv9nbO4yta2
8gq3r3ADV/wwbcAl97epo1m3TjU51q09+kKTOIhJX0lWRZYgj3UdxptrngXLxVOgfIDmovdX7BI0
PgLoBvvTKHMRVsmg+PZy6KRnThfJDs3ks9A7tEeJJ6vz/Uex1b0tQowpGolAQUgaku/HhFJkoNjL
vhec3Ii9w4Wip+DCsBl83JSHshOYX5eZmfM0u9likOs53RMxPsL85RsCYSLezIUzyuz9aJsAXgUx
lCy6PM5eq/rlKR+i+X24mAUvcNhrrxNFB8saszUu7o7IW3oABhP5Y9ixbI4sGsFWL+iAgUERMqaD
74fypGyPm2Fg+WhDD7QKNADS3WqaMzzElG4LjV9cd90FRHHy/EVfNy0QfIrNoeiFvChBgUEYUWH0
dNwRE/FFq2OjWnMZRC55cmNfFc1EDzZSz48hYIZaIh6raTnGL2MxQGlAIIr5zK/qXc+yRNmvDRqK
MpswIJDrgGlmrapjIfRt8yI+slye6R+9cCTrUOT2WhceXLdcirVJoS5ZoIzu+TYg7FTqL+8An/Gm
0uuB7HPbseCl5HqYIGp/VtRILT9kCEXeheBU5WKCnDqpI2zgp0GTU66Hbg1kNWOA6xRIOSPsirrW
KJi7zX5kyCQcrV2y/RFlGypUdKP/L+1NZh8Y610EvqS/1ia2dicWwpUIrLP1u+kxYv/1hTlltps/
hELccUq0LgAnIcDcqqWWaDAuXPoaqEChNVO5LxOpU3a+1RQyGvbMO5a4Z2anl+8d6vlHk8ELfRqh
ACdpE7vc0Xeuw8RPSRZ9aWYPAlif6ltBBwDQbA/g5cADIUaa9woPPwc9qoUVsk+7JyuBU/5WzRDD
3x5Z7qxf/SZgZ5lm3kxohRWtfUvtc88znDWe8e8TsxYI3DhVEZb62weFCoAYGAVIvgkn9qDJft2D
LN7zSuIM0KxcwElz9N0og2PZBpR1zxRL+OxNQQBgXHxIMfSWUlg0rWA3YwHAg31sqSmIC1mcy+vU
pxQxKOhPtuBkYI9PDLVoWEVDlol/0QhlXKJMKE+Lad7t1/GgRcPgeqNqObXxyjLC2/bOLDoCls0K
ziY1HQw/N3Pn9SM+RtxgHTQzaroGfp04u2RR+Q1pi8o0qxRzrEQTSCM+YtNuWCvfrtOvs+DnRLWQ
1DVXpq4j0LuoSagA7PM82gzUHT3nbQ0+R4w9VrqMZFU2VzsVpaHrsb2sK4Nxsqpo+Q7l5BPtWWPf
ytsFxPacKAn6nxMbvxKlqeuqG+Mb9GtpKBHpllzVcyK/6cwsk0ZoarsEhtliFu5FPK2QUqB3cn+O
dKpdi/xi70AEspOUGFP03YYtcJdaOGV3zOieso7/Hba91obd2p2OiGPWxEdzWDsErGnbeyGG0ODq
z93H6RGfh8nLmmr67UL5WxgMrIq41kXtvjNcCStWB6CIJZONgxOUUT6ZQqVIpfmtu9d4V0etn0/T
bf+9/HgJiBfKrO2oGhInDXS7QVSO0GV4dYfRL+L+ZsHrr3jtyCKkZ3/Spnq1MUpZBklTXbZQtVlX
UJPpIUdX7kH3/s8tFgUih0QNMXdsnDnNSZEtWcYE9ardpsANSlW0U/A5aXkecDeCnUwzQO/bCDKh
dIWNIPsPhHWbyPil1hHO7vvcIS9UTNImOBcZ1eWIWGP+xleK/5r7IntBVlLYvX3PEkje+tXon2my
dkUVO2kbzYSLNsfX2RBHTJAIcg4ZuSDTHP/hTdi8t8FGAhbT1fuY+Akp1DvYfYMTBhSke6kTYnQO
B/bb9tiq9niWY8HmXfUS6FQcKnDRR5VEuixc9L4paLIieSxC+Tt21qKIT9iSpNz6tUDsILAwJIae
87dSUqiwRS/FkB3MT+aNkJnpiEtsx+iAXG+iAwj3WkNichYyXqpMMOE7lG6MORg1cQYI/ICi77M7
NSdCGRtXW5Ar06r4e7Ipv7Bnc9eh3kCWPFtVdCrakDe7i3gRl7KUx8O0JxLDIf12cuxQbAuBVETK
0BV7Q3O3Sa2yAd59ePCxMOyyf8+Li6kYXkqmaoOwvI1G2htr7FdnQXO/vIejyTDOcEPJcFBto5vk
o/9Qa4mNPxd5MmxmoUMqy0IXBS9gb1yNts+nETyTUvBNxPZvmOoRTFlOCfpG5jny7auQJGWbR2Wf
Qe/Yzh8CgQ/FnfznQc21ocOQLCSevY5GtDgAGB5OPsnElMKi/Bv4gBgIRHc55D6syzvEkgBz0H3j
+c9UJJUGkp077MM747evmhONiabVvKBq9oXSemgWRPMEjzeW9JCK2HnvUNLrMfKcT63gfNW12d5u
jVnHBVPi/wKmwFITnVLxuQac0uTeL01gEsILythU32TSPLnrOxJa1sRG3H2zQqErYK2cGD4vUV0o
JJAg9zcO3NEbrR6MoNCI8HK6jvj5y8gKpiM/N3OM/6ZVQXteB28D1qm0jg5RPbFERzf0JrUH5B7C
I/dWvLgLav2vl7bQxMNSGr8JlIWMin47h3rBM5nNPpIDPXkstUVMe4b5W/DjaveUtQnOv1OpRtPS
wPWIx+B/zS/FGdS3EYyo292z9SjpQ61l00679ZBsxj7frS03bK4BVVjUGYRdF56RHwv16aYbnedH
+CV2B155IZnM9JhHy482KvDB4BkirmTYLVkrcwrwt+X3g6NkuGvPD1FeX1ar6v9R1yg6Zkv+cyWE
k1ILQKYFcciS0EhKrxBu9rveqkxGt24noyvtrecbkh9o6xBj4b1hoxByKoxHTLofRgJTwOjmUGpO
adwodX8MCt9FeDX2vw5fr2Wn5xTCRXT0D15uuveiXxPZAApbSMq+RKQJr0X70kFpWfC5nfnN4ybt
KW7k2evEM0zuKusDeF6h8DJm5OztgFdkGQLSnXk+Wdp9r0i7pEywQ4eH/BZhSsuiLsNH+e5vapzJ
yFpCY7fdAGNIrp7ob8+uolI5QmR9cz6WPyjoWL1UpYBfqnnv5a6SSNtXbHy9rz3DdW4OCNlr7tth
0wLX+WDqlHTw1m/keP2ppoGuSFUjIl+JLmRpXwRe5JlLFPqZjeN9fN9WpG+TfYA06Mz7jqhKS/mI
9wz27Oll38JtoBl0VaZ/E4b2hvygbyXJDbvbauDQq1RzGNMFPurAzO2cUPosVmm0iRTAiEdUpmzS
8z39OCRb0RoEud39xRUktuNaVfi1fZ7ILZFI2cDxXcxneT/BLQyTaUGVpkugqYoL8M1GVOUtAKrM
4qPZ+vxfth5lnaTMF4eQBPrh+HfVTXWZafnK9Zlgdh3/NUKnG8pC9bXlzZKqIcwDyPsquZtNTrzF
+0d4AuLi3C75V05n+h0PWdquHjC3F2TclXQo6+ewcdympuRgIUQp5qtS8ayUSc0EyeAvvAt7kDo7
3toewD2YBTfvkHN5i/9WZ14nqHbuTqt0DPaw6tmvMP411vjvpG26A+I6YMmDuTJz8+FWITDYSCKc
QfT9tJb5nsDpZN2SIuPvgH6MdrCXf2BAV/MhPUKvwMGUBOjUF6qgn1c3NVUshy1L44oPcG4vCIWj
jkHTjGfXDMdKZGv9uswkr8AzrTn83HKePUT5j/5CM7mioQhMGS2OOS2mLBV/ThRWAP4w2U5XEBCc
hnn0QlL4UStY01cNAzPCvTSB3XueFkQGWVEmk0YtFroIxorNo3yUqEjQrmdwrPlcGiQeZO7dY3aM
GRUDubD3zVQtALpNed5ga2V/GgKTOHg44G4or9J9mDRJT3ytowD4sz02d61WAmqUnl6gVDXSJohP
xUx7oximegjxFC4OYq4Ej/+DuNuznMjdU3chTML9/zjO0uqKwaviLTVyl8JPH0gyuvcQonz35MXl
DKShcIlDm/MDelUooaTmnJZrIAHc8IpsLLE1IG/CVE2thHcwx8fbknFHRIvuFYNRCZ82bssz2VK5
jUBjnX2F033lJUihVvdZZSeAaGW4BHyDW5L2LIGiSKZwHBGJ7YuPChX6zLPHYTuYyOKRT/vSWPW1
yEcM8RYAFJO/0kcRLuefhHEB+eW9jpu5D0itixq6ZgesWDRQhgUt/Vr9zBH0PonLBOcmF2jmIZU+
424PnhjCzb7fvCYLkuekn/qzXqotDju1XmCegkv7M5s++V5lVly7JTsyOkrWAeFnrnvHGym1lE33
9e6elgopHyTkDyUlwFIXqXO7nf0ha3TuTWtBqY05xKwShtbCOhpokp1pYWk12hnh6xUFuTKb2QEQ
J+dKmjqProgz4jmGX+hjzJddrL1ab0E7KKgmfgcmnEuYKJRRqvm7ylZp4b5GPdKOTXfOZ0MQpLON
EjqCgnVW+kt8Y+R/InhmfpfF2Ec4A1ZHZhinSWCS1BKpsxn6CEcDVmpPSN0VFQokZXs7R83Z2KUH
Z4B87yyA4AAlIqZ4wQwVVR9BYR2hsZBmajh2K+zvR/qW4/nohrVw4+fYXvFr63IRht+UTmEJj1uJ
YR3oUJ01uvPi1XtgkHNJWCl8op0Ch7M3stTD63wuT6Y64v4e31FL64Bn35m9FZ/NE9trBo4kUDge
JtG9loIfYs8plM9M39AFE25jeFxF//umOVPkL41hTPZJz0bYyorUXG7A69voOnFVNAdHCyhJXcWU
gIJuLgT5NePkXnbMqZIODJ1lyoBCVnbLP6SYI9FxyDFztmJzSSIdPP+bi7MmfjeCnmsSMNBiuyiz
rnGgIxLtrGMPc3+zlCxNzA2DZ9LxryZHdGEry3RKF7nojajubVNH1dwWcOnylSzgFyT2yRTH6/mj
Phv++Ia9dJY0hzROsItCY4VevxPP7evwOr5ZIepVJ1QMFAyKFEEZBsxMCAGaNofyHHc3YmLMR0gK
ITE7i60GXFgwi6dndjmDxJRpESNTHAUsAE6gIsaiXJVv9pWR2A2UkhuhCtsC2GCEdr0fqVHhXsKo
WAAhCNShyIUKTWwqEM0o27GYSlG6qv/kxjhXtnRYuKf/VmpHyNZ/uHnXxxA1raHZMszT3xAWOOWK
R6IpzNmeXquw3RcCvUrtdSLQ8QNyM6qLkxGoLJS6Pt6HEuXuh6EyaxkjXq/j7RMVX22Jj0iDePEK
jqOwwry1A9XevdhqCDwnNuhwBBVEI/egdRZoQHM0FHy6TQ7Zdi+utOomRsnAEw0+zzIYes4ku7EJ
LN56HbZtexvB65crSSbAblB8yB4UvleNe9G2ZxZf2yke8WgDhEGaVg3Y9V6ThtaBZgpIXh//h4zu
JkS7NTIsFi+R5E9IklACjsJGyHyq+oksx8lIrZfWN4AVQz41dMoaIJFar3JDuA4mXAsc/VEKE6dj
NAbczqRhlZxMKU60jIhPz4ISdWropZ2x1Qypda8JNskgBSNfXoJthrM7VzobrkiZNnz22QUaSvXM
BouMze1y+8MpEUKszsZlBSDNZUFFp2pUe7vPeRTtc407xMrCPKNOPYXrZ6Y5u5Bjxfy9GIEDSK4N
uvugP/yd9sg6tgHdJleWB2msCuvr0XaZOhdnlS/6anqmHH75mfbk6DH8O+4bwWaO7r0SPUXAVRPj
Vx8umfBUQ5o/MyVhCpt7ehhWx04mf9TtABupwFuj4UkIGSm8iVuGisucuOtuxwP0rAa5wdHlGONS
zzC50LjEjySGqBA6YmSfKHh1nIJK3pBrtUh5R3SlSeS+y+me/x4HD08yQWHkgGyIO6f1kbK3t+ne
YuiFsu5Hn+rjXKoaw40K2jYFlEKUDfCWAoCWD9qESMZ6e1WDjPgPeUf0PCxST1llKvPFjWA+LGnt
jAWTHg7TLZnQg3Mocyvp4e4Zv+rA9mHchs6naHWoVPi069wExZynrDgaWPJl4ozDRmBh6VB6XXBP
QpiPcaNui2JcFRbJWKoip52weuiEVCSpzeyLJfBg9QlYcEtmy5IUABiKdziC2sFd6pvFuWhFORUh
2nl7WXbkvULKGq79vhtFml+oiKOmUu/uRAXmrMdYDg12efRpEIVVFSQwGxdQeAySH7aKtk2S4cJR
uDCqnWkeZghE3N2PSalXc7gjzDo/TO+JCbY82Y+anS1DNsLhVvujFLkXPq/60ZktvsDrKLc+t5tC
iZItgYy/EcrcinshhSscKVlUQyK05x81JxM7jk4bgomlGP56YhSl/zKX7N6pl51G8f4zUc9myL4a
0avht6mXd12oNZ+5DbUJ7nzSErwV7SPci3kcyzS53an9Va7ssaKS8Fz67Jd3w/qHXhl4QSdhGIcb
jBYs27ii/EeB3+k8eh3StGFco7gruBp4lyZCM+hy764mZkFs2CLJg9UA+yvkSlGO6G9bbg6mnPoX
a6G1jZHpNBekiLqP8mrWfPaBzoeNp8n0CkJy5O1wUaf/WqLUkXeWLz5T17Jw9VZNMpHbgxYCAQN7
4qQkc0fiuJAsk4e2iihOX9HkS5SBnKvqTKQDArtCEFLRNfdLyhClZ5ZnRjYxLpx2jRHdGybmQF/n
t+b7SeXNxpfVPSmsihogeeX+UPev1wOCuBniWKhkhYVow2eNPrmTNfmMT6RIwMsxE8r3YefGBhGD
kZdWRDJ/nR6yWe5+PVYAtKCxlKgCDPQBQrbyNDI73UFHwPKvaUnRX0Anqr9p7Tggkag4b/xP6lEo
0pp8xx1/rBSIqp/fYnrqRKiatEw/HyobpYIdyFEVXt04PX7TsUXrzjNONRcfpAOvx3iUPprcuYZb
jvpA61pfqE1iAfc0ULVN7vlD6i9EqXRjEbFOcTFwyueW2XZShYDalYM4ksC2Vu0L90C58IlTmDnc
tp23EGGcx9lekOh1Urat1uR49+8qZKlo4Uwy8yq048o3LpPNWccob70tslyHbNuEa2P/hB/BWNus
Kau/6a6+D/UCG7OKWtUEtIcZxI6UISmb+2GvSFo8qnlGNfEcND2y7o/ex3AUNFqwzcQpsGUZohe+
GZOkNPMwG8FhvlsVYfgKd2SpeR1bz7vdzKDCOXV1iCAx9XCdrRoi1nFBWYC9N14LawqmB4UVeez6
RPesoryIGYFHQS1MRzSC/ucZ6OaK2Hx4WrRR4S9ZhmWN0vAbqmdJ7/ix7WKo9q0oeALX5G4TnAGC
mc9O5m/0x3vhtTUNCRs7bf46I9JOSEDy9H4gwxEHtKhQUz1bhBT+x0sG8+lPsKQk/YrSo/m3AYW/
S2Bvyz+esRPQYffZ5tMbMHss/gJkrorN9gK3M4MP9XVYTfO2NJA8R/lbmCA7cQVW3rpC5R3XzByy
rkfXxs9MbYDeSAF11CaMGKZqLgRAIXViWDW5hvZqvoUf/5YSMqpGTDyo5zzSc8wlVSmgZib3MBES
zkieUBTGtos8E8ylBTRgShjNr3HUicrH3MhXzQMB/muUXCZgGhi7MO+CocUidAFbrGm0tkewI6la
BHwyqe3lm902jjpXWyyQmeV7W6zm+vuMUZA5kv0qUlSpa/ozoSBLrm0mBXKK6Ci8wDXfSerRz29Q
i7516Xf8bZLXAwsdcGuC06dHiNy+Pn7eRHqNn17/H4mS3B1VPuNnylJ3B4GenQkJu7P5G0BR3YXS
eOmDXg2YAvOYpA45gH0w0fyeAF+WtwlwzTTP+5H8Y0p/rb3HeCLJjOIyATPypNzlUmzbobBqkKds
7Tsm7L8UC+gLKv2ZwzSypv6i9PIcOFTmuW6qSdk2W2pk3j/xAg9H05+MVgDY8n8izkCBlqzleUG6
aidcLD1CiE6RP0+AswfXzDBgG2lFgz4Vu0neUDRgI1LJrmneWgObi1158acTNhtqDbdqFbjp3P6U
66uL2VDMMEacI4+A2GUc/oDmRbcF8l0k+FYjxJNLoqmtagknQGmpq0/KmosZmQM8bw5rA/4Toyww
rcRmhBR2b0Ww1uc1Fq6vq7CFcgEicmbnD2X3mHoWFAD6GE+YMuBxSG/+tnPs28rkuExt8AxaJe6d
NsXAfH4P5wZU2YF7r8T4/34UX7MWhNzZ+APaKjd59E0jdSgP+pejRwE7zWrppcPH/xicAQAM2qmk
AAQ6KJQk0ApQ5PRr7ooETri4tFxyfB4F+nvk168lc7EV8/fbvYyEv31BCuezZ9gukXzCL82V/pRt
C5k/lXiMYLV7wc4zoknXED5SIqVk4xG8/W1hISoe5gRgh2M/r2e27Ru/CZdyEABK6ZV5kLZucnGF
uiq4oFJxY7GiZ6ejzCXkS+dZlnH9Uq69zrRYW4vSgiWIIHeskMyZAiV2gmvqLf0SZcWO4SqzdTIW
EihOZ3ZICOXnRBq3oRFscjZaeqw+4eB1nvQQDBjZxPJL71GhOE7lS7ZiVbWjxHxXmfAYV+0JeWHc
fcEqgQQjh/suo8jc11lG9Whg0QyeoEonpV31Lr+Z7bj39v2Aon+uINQt2MVWV3fzDXgB/P2BoDYq
uJ4C3/mOBCZglHmxYeKDCV0MHsOGf2vbqEVhCMhHiV1wQ1MuUySSRqitZiO02ggKNtOgNwWlE4+j
7Kv+ov1gtU0sXcUM5M9IXBH0RxureBX8meRkF/L3qNEmWnyu1W3jq3DOx1dQxVlmD0gXWdw7KMbc
L5C2YCL48XjLCDPN90uL/1ZZ4qn8befGglc5b2KSzEbHRhR4pOAw89Zs/v+ONaGUazz1zBFK82FQ
zIJzZzc0SIW9KvrhyhcIjIGrgMTBnHKhLNRoX6kxkLyPwHj0wm83UAGCT58eq7IpG+AS3LxwGVGF
/uO/ztDx6nu0mPi9B+Hso9nLj7bXXnn/bxwiPYJUNNv472TBF7d15HxKnuJwH+lwU5Ay5EMacTu8
iSYMmMvxgF9Jju69EyZ4XROZ00pWabNJXJ9zBxfs5snwy+T56rM3qlzsKmht5uE1yJgQxBC0iuqF
u/hlzfPMLfZwe0j1dPlGc8tclbHdGg+K0csbF5o52zv67UDNlfhYjHfAoG/qSAhgGzcqMGcGrDfB
WBS/NXIK4UPh73EOvf0douV91QY52EUlTdGpuzru+5AKrx0xLRE2tTzFD8aft6svyKdqi51rgkdA
ZwnPSNxPUavT9RQ4SpB4o1PFGuxzQdc8XzniTRBvVqw1nZMoBGvsy3OYDLkG9ikGtTmVEqdnLmsP
mmwCSadQV94v5/7bKL3RSbqC589kPQQHj5FX+EoxFLtVuUgbAgjWwWOzpmLC+NULhE+9+1+ubc3M
fM7NS48P+TPaJctigIt6p45UT+JUNaCZZ4i+idBBTH2p3bbCxvwsnpvJAuz7ESHtzXFYAvBTgkDp
s8x0/bfh2HsbFnBCKzrLjXDjz9O3gWxdr8qAxLixUzxf16uSSVaQ50vnl5fr3cGxt7h+fRRkLfdR
FMvv5Scz6Tn7MbJYnG6u0mO5h0DvKUTZcy0p2D3sPeLR/xcc5xY7C0lnABpU4kARpsqE8liI6ePe
lob1rYICo2cjVl1e0AVqeoattezm0n+UQtPxJSVTfendNxu8X7JLNAFflY6KAU82sZ392v+eRd31
iCfc+FXJvVHEXG4jD5mouMUxwk+VUwhrBH9hlapdOvTelkVyud3ew9CC0FrWQDwIiBqUAdN8XED5
J0G2pZvKV1G/UiRD/vDbmgQT+gRDYdo6i7Z1rMkUbJGQ/2e9+K3a/rnm7zyiFESOpgsqI65euAtY
P+KrbLgsj/6CvR0FIXQeehYENc3omCPgp+fgkmbSjejvwgWJoRlEZ6JZyMzEjGPs/aqEOSJ1UHvR
07Q19bTIh7pP0h94XLQP5h9EO5hFOl4DwGqiuT55wKUiIJ6GacKfGfsW17tP8Dc9ZoNfxD1n4vU8
0k8Qb+NTYH53LRRbkLzyg/R2PtKqESydB1UIy8gUAcKCtDH499XXNeRDcOpZxWfyL4YW9B+eFCJN
Q2EkH4ZDq877NQcKmO7H0RJ/B701HiP+5h2dgd70IGstwxT9lEWmeeGRE9lbq+YendPhbxOiobSz
lLwmolz1uCIqHbOIufJXU5U4w3sVVWmvilXr1fS1l60nOx4evKCgs1yQamms7pS+4YUjM1nU3DQ/
Dgtrd3/qizWAk3lZQD+zrl5gJ8LUNvg1XroSnsQSG+03IQm29V1sEs5rVRI+5TUo+jk7QOUX2HcR
2AHxBY+lBwMuxsDs2Vln6fE5DXk8YpBrG13DOmMGd/G5Sxf/fCuWKjQmf+PDQs9qAwxP0GRNDwW/
r4mLlDDezsgxwRxvH8SgYRZdS3knIdJE12l7Xx+KNdYJNNvWJmwt/B6prl7JtNjvsqMt0dkF9IF8
/JlnOisvsZ0sblx0kJVadsyqfajn0B6nlMj8oZDJVfsjVqVMIg8K520hq3GpL7q/E2UroYGfshdE
4UxmwB4nqPZ/0ZbXHwD9odq2NkWAvfBPIPlyK4JeYz/6kllXzyLmRqWo56rid9xn0+5vpHbe8+OX
afChoYpKK/4nqKm6oBy/rjWjoTkh8WaLOkbs7RjOzUSsql07tAwaef7w2kY8RYDA4IuL9p0lTV00
LvjzR5+lxhMntJG6h/GLbS2A7Y9hFkW0djmZdtAOyPQE2Cz9Yv2HLUedurT/A5UiAK7YCWLFcQyn
5P5D2ChzswSkLtBCF/8+zDk6afQlhlpFRSSUnKSJUjSkox2qofNli4/bUFRIOU9kfTcwyh0s9gUx
k2qz6QRi57u6yyZH2I2jF4X1pN/DE2oVIqAq5zwwcP1/Vy1/Lw8yuOdm46ZrUOEuXUj1K5IsW08G
M7rY6vqE9UhkfJorPv/2XRoh9IgnRlWKs9HUcVI0NWNFkFInjrI88uaw5V6IpRVUbl7pyPMyR9oE
GpBDQP0pxavTYoITSIUFZOClhYogczqDomjaC5IxMfNVmUHzE8nR14UUmKg9ilzHa/CZ9NcZH6Q7
tYG+vosnVLd3GXrNi0gOwYXxu+iHMsEJHxkYGC/vHCXpxxTSmgnGyLJbAopqOwu+yttwD7yXSGwe
puUFAicfbJ1xZhzEpSsicLqEYTgqb2y++6Ro3O1LtsPLWIUT8GQhyafkR6qX9cRu7S9JFnueEaVB
sNZ9P2NWgP0qSPquvQ/QdJZgTupPkOadUTEddwzLVsSH3ZbNnJfA+dcC32WYSuyaWTIc5+QrGsfo
2uKbQL5pMTLWySlpcR5iNzS7JFGu5T4mTtuqVB3Hsg7ZhBnidzuRcu0vljEOXyg9uc6WAxOPfFrv
IPcWWk1LbPDJWzJ3qu670ebJMA6pkL81F1YE6rWLZMjTg3Q82X3eJBqCN0tsB+wvN08iPEmhjFz5
HKxyWHmo551q1RNhD8Fd6Lsi0yKSWhvrJWeGn3PYzMw1XPqc9qr9Cob1Fzq2NdPEMSmMvMXVEfH7
Ye6SLftf7N+du4xZh8pK7YBmIKe9wHdiz082XmxNKfOLcQiE9s0rWDlIknFMBQkM10gTdT98rYhL
eX7KJZJiIEAKDIc24+bRzj8V3kIqNxWdb+3Q74aZeSFF3eAsiHv1YwULWhFTtYJxAs11h3qQqmJG
YlAdd2KDxnu13EGrg3UZxGVZTUOBtYD54pxwfhfb1XuMnrv1+jKmFu2CJOOrjIAS91XcRHPE9/2b
GuTU0ikIt86HLWCeRfcHfmOwjtUIy2TemfpQkOPEMf6gFpZmSURhmBExRZ6ZxXtS4qiwIsYCec7N
S2YatOJ5zmu34mZScIf6FNRMKxjzq87Y8P3CleKm00zGX60ZnDZHA0PiWlTnqkWX/uO9tZdok9z/
FbWX3JdlW2DcFUq+UqnZCgTkYY84+w745ED+YuTZ/vmXNgxgKKCNTzaRmSK0N3RDtp6XykgC6ESO
l2ynd6FPrnBACB/w5BSUmXGZfmi8NHbHDMftNIK43WU7AuRiTSAnjykufxlW4lPwmoTisZTnU9X9
nQm5WZzupuRjqB1gsflf/cB7rwAsxQmdfQp/xkwuIMSvsRgyQojNJZP2R/OgTFu0Xpyi+btSgJT2
QAhL8cK3y4KGM4L9cVYG/g/DCv2ZXYYp1fMc/0Xzo5DrLsoZpMXwcz/bRJ+IZqZE6GVBp5gyjgy1
7C18B0SKTLjlt3U0OaUaduzNrJfFy7gR+raocLdiWa41NkBuFLRRgWbj3Oxy+uOMEx8tc3vdVKpm
VGC/+pVE72FSBSuBGCgxTiCWj/05P1LHa2ihqMIOeosu2EBM71dcHIkUOV5GKS+7VYi+zliA02LY
lqQFuAvfVyb5gu2snmWmHM7PjxmxIA0xb9vNOOCgeg/6TUpYccToxGD4fDgkRtmoAfLRseKnqynl
H+eRBuD+/s3mEj2G9iGg4MOPHsKuGuJU/EAWLkKOYaHbC0Dl14+Dtru7PtvKs7ULvPodYfy1C3tz
DmPWcc4DZzGZB48IsDAaTg5lnktDOLj2HSyirAZYZm9xyV4mbnKy5ViDY1QPBQr4QLHq69RjALz6
U6q75Ht0Mb6XruweU5vo0DYHM7U6CNHBr7MAB35wm4KCOefnPN3wLYtTrY6dNxWNLAioio7udgpX
9Vow4W3/bu+GQN753gB++9j5AlIpu4OaoHoZDO/gj1sF7SqsjxrhuvpM5ue8gTIh5letRFXttioU
5vlTlttnaXYotgeYmdiYvgexw0nOnTjR1umelCCBExdhVdg79mwHg9BVviQ0dUvJhHhgN39eRyfD
lkNnXn8C71M7FpXE35qKLk7YBRfw/6EFb1ZtsIhxG7mYPtcmM2plSZaK3FQ9YSkllgxaHunimg68
mVan+UdKlkwQJLSQ0rI2ygAnfM2SwCqhcrefsJ9AlrChs2gBXjBFwubTi+/3fI1FlPSS8BTAhmkf
hsO3bjaRfGO0z5E5GJQBEpGahfmLw/lMouLeA06fp9X0ZgWkxhy1EKE8lRfzQ0Uw9wNk33tDz0Qr
D942WFpxG7NsZFexL9uIxGVmCTJZOZcjEkeGOsr8k+VIMq7EmfA5y1u6kdWNBPim6fsEmMpOEwpM
lBpDhx34Xa8EiCJYql6+wmpgyS4FuzO6Gyege7aMSQWwrDu6LNYWBgsCIRni0zT3SAqbW2sxPORp
dK7PwFiuWFJOKtDF69tQ6hyPk5phQuIFJHt5Vvhf9V5a7EgTT4AglWtj/EKeiGza+82Hn84crwwX
NHurUcsoH/jLB8RKBJQK0SorGPyijLKe+Jhg2iw/DweGxk1OQMEEY9gEDsUuI/vv2EWgqrj0cwnL
A/lXT6MoDVrTHpjFvA2W48s94WKShlAzsIm4eXvAiqGOErnEjMwB4lAz3fdpTEdxnjsQ0OzYrXGh
6cdCL2InglAq7OiB/vLTFehliXy9jNVGTquc1Mlzip+akrZFrXvxXCocAleihCKB7arihcqR1Ppt
Ok6SKByJOuYCyMLa/HoqWWc4+5Dzv1oXH7qXzHQFE+a/sWs6/o9gjtsWMf0Co74+mHfTDmgjY3NP
3+o6HPWI/n1aYTDEg1gM0lOMbWylcNsYpZ5nEXrcma56YWb9milZvBSTAS9rvC+opdsv02dwpIA1
0EtAY5mOtRgQv4reufU2XCAwweBA0vlUWVSLsVcVQcnJ3Q7ijetf55KcSi1bwYJcT7h/dnxe6Dbj
MiCI0NXwfmH0EWZOp4+6Tn1ivTWvvSATA6DJrgYm/kpRnC7+PYMqz4a5RikrXHJoZAmLJ/62g3fH
/0LTZ/OGSlEUVuSyAE8+OgzpEqO1gHMiDQAFOw9ir/iSIkBGWIJrb0iXxGFXgff2ltVS2CnwiLz+
oq9qjgVkFw/lMuZXdqncuYPqs+nYXbDs8NJOfHUOvNLksOqzhMAZ1YGlDagIpcjFBdl3qB4iCp3q
xhrBUhKwd5iHSKu+MTBYPXE/b5TM4ZbQ+Ll+6DvdAWbsBGd7hBkzWmD9ac1sqUrq2tmjNS82tURK
aO1ywwSQvgEm2ig2ZVFNecogJbJibUSuE5fulkXitLmPlvGORepz7D5ovqDJr2yIwpRLf3GM3qjy
j12YMQBHaArXqZP88Iu4PR7dZrpPMnvyRRVWPJkMH5+TbOsFuf3bAhtiiBbaSsavTARxXoOvkFI1
SQsNZltnRzlvg9P01YEzMO6HpQgVQQxEVDw8GaNz0xwbOZi89QJBDAOOSdSbruTXOBl+9eiZvkFX
bhOyEC4ypcNiXVSglcmwkIuxAFUd+8RArqWiAYjYexEE8qm2zJpuA5kYkAoORcbHp3PCV0YKP8fw
2W/pdHUTSLBveEU33xsPaEYUmAM1pzeMNcMZGO61C11yQl0M7oHKlDor3DPgnhcHuVTs19K//gyx
zvOZPIyeKaEEJZVz2oY0vtj50vjbZpfpXpw64BITcpTPbjdRw09Etxt2Va0QSp/87TcpXMrAiIhb
QLYbKY61UyjpYsd9YaTHgqTwPR/CTa6E4FAwfvd3aGJWTU5Es2UYJnXza/0ekwvb+kFc96cIz+00
HS2wat0wmXyngoeyvLedmsE/hT2RSroAIT4bijy0zEf/Ijg/L8/xZFoIbOsmloqdeDCUKQSV+tEg
69Q2PmsWtJJTp4M95en18BYWd4EE7dPuwSSpIPXuOlQ1DxdhCriERD/B2vuTDa65Yl1YEld2/0gi
Ymn6sUf/wELSzDK7VDh2u7SDL42Y8qpFdbLVTrzMTB3X2cYACE+0/TNoXkjBVgfHOwKybxOMZ1kR
Y9JJ9t0HaLhGkJ2ZXXXFTGMlnaEZWG6Wz+vqxBBpONiVkR8Q7VHDKvKX82klt3meODhF83B2K5cY
KguMN7A8TMqGYkk8a+OGQHP8+a22fwB7C5+wDr0WCC0Fj2DiMD8pMHP7unPFwo8xGwGH3lcw+afu
msRHDLEKkpGv8XClQb/sbAQn/2H8HqTyXF2smjEO9XhHIuiE5GxZR0sJUMYQa36YpRhYKktRrvpo
uBjOjaq//50zHuS1R2fwfgGsrj68OtYYkLWw+hqznbLiLA0LuqIZ0C5x00GH/R+sb8zXae6TF9rI
e472+SsKBJrlV0wRkc/rCmVGW+1w+lez6uJ5ghNNrX4k+wryz64U9n3WuH4lqQkn+WRSWK/+hs3S
AtmjxfLgtt32Hxyhudc7A2BgBFPi6dGhR9U8m8qQ4OvVsFI7ErsWCdVtb++R3zOPk9XvL3H4IwOl
BxAnbYyKM/FIjGfLkDDHxOgyUrGPIcP/09kLExhve3FARMPWbTUDiYlI9uSj1H/MiStsJc/OcDxT
2Wfzib+J9Dc+PiJK5soHhhjgdY45aeW2rPuQvlTTJtLF3AhXS8CAy+l4SPYSUWdMxuXvjPaLyeLb
si9/aqEHkyYezT7O+m5sUb1VXb9X5+tSE931bFdjJpFr8sLNgCpO/UVbmJQseYYodI/CmQ3KU6Lv
aePVlqYCcgNHRP0rku3dEiyvCiPrUAtYvQQKqnJlpEA6UEpW4tmFBg10/NfIj8ikN3nROpcaZ0s5
U7j54PnuPP7n+dXonnJJFYo1aZpNhVDWwIMBbxbBpBUVJAabNrMwsUEKB4Kn3utTlZn34WyDYmwj
Rm8aEpKa3x7SXnvG4YmaFzqg65XpB3IxBl/breA6+92CWu03hnlaAcf9+Cr49ykdlzNB/oghc09k
7i2JDK6xRWT745Jqb/S4kR1ycJEDtKmVNPRL9aPZEf8BDcQ1YBRpGpb2B6g7RJhtVVCMi1Z0cr+P
Vrj62JISeICJab9hiBczfpwqETK8L4XqSu0E29zW5GvOQK8DWU21GW0WjNKgq7wF4j4v4l6bfCwf
4mBJR4fyhnpLX3IvKFN2AQbr7R6Lv33VhRVGsSmwViP6adXZ8ZhrMJlVV8vHNkUdhw/GSxqbt+BG
+WPkBlMEF57uodDOJaTHQcbkLg3wBl1hiY/GVXdvjqlZE9gaItqOExraTuVljsfGy4jx+PjGo1i/
7BCTgf99YuxN0KyVvVJyGNwQ52HXR5MoY5g4zCStSZrBncrbzr8BwGJQKOZNukhMrv2cPnYPuyQ1
ZwwMQqafGNn1KycEa3lQRuQqzA3YeZO4Gfs/dN4ZV7boQoDgjzoiJAJpW9yG5K3TjztxLyr0xNb0
i+z+q8qrTqixHV1+xzlvnf+KYeloWB+MMma7wiY7cObH3XOV1Z9BcyVsYKoaTLPhLsLQP0wEsAjF
IOpGTp5DvhFqNtXWH0ykkdiTXEbdiQ/x1aRLQu3vwa7aY8PYcXlUCs7zzZPhluFHZNx6ezyMKR46
MvAUdU9d5RfGqjIwk5gBAr7IRDrfpXY1Z8gNhXOTKO9Rn6GIOQ6QL21X3qZV411AvIK0ROXJfOzM
KR8iFCcyUQ/2llTUQ1upszERkjjJTyEYp07jbMEuexvScRdedtWHlF30BHauCXMe+gcAK5Y15xae
0WudZocKw8bKqJXdc2EeON2DOaRoWnECzg6CMZ9fIVMW1rdRBwBlTrEuiygP/uM4U/anQRnDhLrm
HrFgEgM4KYm9KR6Nc9Z9meaVtfe+hNN0/0i1zV0QGcKx55HJqqpm5hK6TdEm729x79P6nOUaoK2O
V95ywlcs8BhCnP4CVgXETGn9IRkDxaskvQlVLyJz+PbhU9fpBf6+P+KqQsRzzXd4vAFHl4mfGooU
6Nv0kB4IKkHBJrLB5gkA46Z92rBb3vQX4eVicNSQcBu0hCC3DxbM/byJrIhJLZxZgLpNkgw7hQT+
nVH0TDdoBp6H+9SHlKJ7C3kppFyNZK4+XZsq3QubFPSejljmMA5F7M/xxeCCW21EqGCYWCvIr7yc
HMXASAPnO/DzRlvd98XeGd+yAl/pVXdUgjQWHe2zgnfgYKeElNtiLELXIA72zdePcpm0AsSsRSZG
EF1+FPt1YqPL4PU4rBjpWb2IRbwHgaLWORSxDqWVGO7QkOg7M3pGH8IPMcQlEwyhXM4pzjCba0ju
Mhd35YvcwL8LnZOYgWMPX9SULeGHUfNPoLKdqZyrn2ioQfSB5CvFJJ2I/cShqG5gw4rsxyIkEYWA
9qkXmLaPFKSGfAmNJuSe352NwCdAI9hW8vutIERZQg5nCeS58o9OD5eVmh2WBrWRN3Tvg+SJoBH2
E4FcXfDKfa+i1M88a+MMCBQSd/Sbx5vTPj9eh7Ymv68cPKNRLIt9hY2MKrbuy55+pkWVnsE/cdV9
WJ8E+XCbbX/s+tKZigrwADD/YAMkBAjdAUu3TNlTdeHUyTC0DlMT6EAXi73qGXJcGYhjkXdAqMO9
SpkmGiVv3se+x6GO7mOpAnTw5Nu78A1VImnwXNp754VQJPN+jrNPUeLuv19/2o4Wlj2boOXculKI
91bJA0hnfVyd6ar+qs53k+8gcAoMnSE+uHGvFe5ebVu9BBpagG69K5pM5/zM7w49mS0/fnxkSJIB
bpkBWPJTjISm8LRkMqJMEGZRGQahRo845+KeflJByMHilAzzR1pWDccedNfHzj1TNXFfjIF0zFoF
6O03legW/dek5qItq0y/rPDT8MyZLO5GnP6f2ypfe5xoa9OBF4Cnt7vOtWe/0/EDlwgWNfHl15Tt
nSScAI0eqfZUo6yQtYTE9Fdu/JHnxAjETic/igxEST0M2o2TwYNNzS9/15Wc2cFRO774FV/mA/qq
50TPJtlw6EYImmiIhve4b9B2zPEa6OsNMvs7fMPpdDZTCjB2EIiwLZdgL3IQk/4T1bViM+R12zIJ
JKqHACw01tBjgcFUF3nMD3DKRPzopN0alm2uU4JS4+yusGHhsEz4/YLOJU5GMpr3jIFqIZatQZdO
3L7EajvPimejMmJfxZeS/+iVx96TXLmh8FITm2exEyI7bxNtob2OgFAkPsOEimHuvj4Ib4SxA1S0
1MVT0kE2eRtDZcRgvAXoZLL6SYM6yc2IOGrSK/rvGTUvDdhH9KT6SkmsdRVFTNqnYG8uqL3O7/pG
O1ubDOvp6AC47NvmFO5KidBByhvQ9vE/oPnkkf+Fiin94J7my1P+QewmB0MwdSFOvDVByqfcHWs2
soi7aFjdVUeUV1EZccDGqSQbhgdBL0uGy0VCu1H+4BBAmVZZ89n4x4Kzu6grPzxZy9nmVWI8kLR6
fPgSiXDd/tokMt4Eta/D6ikrWc6jmQoqR1QWE2d+pzDyM7oH/6NZ0pa9hBhcV8Ltl0l4ga4u0yPS
pZBMsUgPka/1ZjM4LeRy9Huh4O+Gu45JdO//jCvVpIkTqyG0TaKlDdHlli87chOjCO+p7AJm07K+
2ASwp1BLRNVDkPIUQnJEslM94jhpMprnxAn0/oqEcKEz9cOCmkjX5cHKmUaiEfDtXsm7nS6RW1q9
/QmjLxMlhaeKRHOcQNNnHEtS20tXaXaO6ZfitOaHwX1Po+YGvQwY52fX+bmlnCdOnmYX2xxmXbyR
U7J4nQIDL80V/+IrJDwNLFK25S+5NUCcVPMcPncg9L1L06eIEEuc/NEUARoHuX91M/wyEjHnmtyj
TLyFwG4enxJTdZrXyTyHEe3WiqFpC8V9JMgCy0fSpmunI8lDoTpE4gW7B2rKNRnHy3yg3pSUab5o
LjwPrg/TTUCS+v4aPsuU7ikalTJdxXvKT02bOtfiAtcHXwbi3TDn1xmJsyddq+nu1zVQGFgKFcEh
N8wiD17tPlRX4M53fgKMItZuP3OYCfUW2zAXiF2cmnNo/VWGxRN9YSFSX8E4Z3V5ahkXQkKagUMJ
EG3mYIFqB1fCKhk4l/W2OCNveIwH0hud05HIZpqoPVBuMZoEFZi3fpqh6i/ALr0tG4vOXPcKLSGn
alI6WeCV7P2kAVpR4y/uYps+R1CDD9i8WI5k5M6sOuZOWj4oAbW0oBhORZRv9sb6m4zkGn+1blQ9
0H2htnmtFbmTBJDxMOz8ZkrBV2liqkcpmXrpvK0Vg2sJf2iPXiN4XM+4m3o+jcltrPpiCvPHBVdV
b/pOhA/fV46S5sdw3tc3bFSTJGGoeSHBAMuQLT7/jxRgr5sNNdbyxZf3wTerFan+nLP17JSRew4E
EU1V0w8ooTDlTzScSShbHdpJAAnwjs4eZOOmQ6YALMK+hwEJk2GhV69RsIoXZjw/h4+VNWX0t4Wl
9YUTpR5LigNQRw74U5q8wA5tE8sgfzfwDWuf5RxgNTLAtOfle38ek67L3KKawMoTMMiN2oUPnUY0
dTll1o4PsouJrGUWK+nx62T512lbvfJ6zXa39svsHU9y/fmGFaUgWQMpB3jFJtsu2HAGOPaj+2lJ
rnvcEa5T9lmkjSWugtIHK2x+BAUsj3PzQQsDsJLwADIZuRgUf6aaWWTc3qyOs2JIOI9D8pqbezd+
Q6eqDjeRe0Leo1TDGa8rZfh7qiKNuYWo91A2+jlh6QuwfdN88OgLxs6VXYiGTUhazacXHQnMnfWO
eCHXLfXD0oTMznWrC1xYS5iZXkJqxFcVgKuLRFnd00X7++URNzvx2ci/X35eOj3rcyFCfaNOIufu
avQIkhE9Nt/P2bwRM3LmJ9rcUoHCNKDG3BeRqHWfW0xYkHCZMkXMs1zXqflf5bl/vSL4m8MxRU14
pcOdbBM+ymlTmUrxEUZr3GVkW4xfMxEzjylGnp6JKDhSVVth8U2IFc3G1o/s7ldjrdlRN5JanZuz
k2SC2VM9wVwPwnl1uEw8IRvw0mF5ngPlgaS0u8V6aSAYMnUVaq5XVhxbzNiYsrkrQM5C9vb1U5R6
vWbCUXSFeTA6Ds+SR0VL3VYWgasM5Y0SEnIRKKlzrpWY1eD5hqwoEj5AQCpENYspeUplyobC23Bc
qTAoGvCPQerQvy3Rq8/D4Wgz6hv2Gecfgi5hcwxKsFAss/UH7jODC6HtLnjZX/ZUtDyQZBRrLUre
JvnyOuAhTYtn9aK9nvydnH9we+avsR0R6TI+RCoJGWOhlITWCdy5f9A14HPONluNsIAqqXSErrIV
1bt5UjDj0JH3E2hm/rV3+b4V42MMZhlcDwL/eCRwgM7IHsKmmMCHXj7Lbj6S+hocMa3dyqjcqp9X
vDIDYudbcs3vP6e0yWmQCOJKA9z4tfdBcx/FxYS+BR0cpc8uUjw4rCQ5KZKbU8qJE1aGt9wFqQ3H
PTrfwGXVFuQhOSUz7YDseAeVXCkr3vKxIk9HOhLKjHNobrd0FSNh75NDFLo3KOy/lPiE5z1cHENp
ulU6o2L+5V/HZbSWwMYlQ/BBOBaAuQLWt71TFkoFcutfeNMiWsAlOf7GpJUzLFcX5au3FbNQV6VC
tfdQqZuRyXo4ID5dTpx+7kIIpwsv/5B5UPz7h39mBW3Vdt6zlFqWakLQEYb/7pEzNIHd2dhp2D3F
WRNCvxJJo0JbDp0+glHIkwxT91zZSdGMYNa39mzR9r3P2WCehv6etBzR28Zq0BhmLL+ONMu95r4M
uyoVZjqD4Fz8Qa4aTGiMJ8VowGKOZRC62b/k/xKZ7vRF5TrEU1b7Vm4CCdhsnx+0hBh6q/osjNsL
IWQt4sUKXIv5lav2qSAZIjXWIIPjAlDII7sD4k8xJ2Ab/OF7qIYgqrPycF2mt48ZZc0BcB+L7byR
o2V6czNB2iVu5rQEhv5vw1lyK8moS9F8Y1k5Wdw2u3qjFeYFIrZOPEav0mSnZh+FpPg7fd1Ly65B
y6c4BmbL60c/xnnLn+kYRCwTtjZ1jGVOCs+eARlMrq5LSLuT3beGBbF+BBFqIjsXa46V7H2F1wGp
f3XbT7vJYKG2KAySO/9CRJQvMxrtlRXXCDmVvhTVviWdxB2YmX2uOlOHT0dL2nijB8m0bxrxa75r
9ve1faCikY2pA4gXlH7Hbr90SRFbdM6KEeY9rJR5IuGx4dQ0xvrWEwAl+9ZXprojWP0Kj9xSmzN4
3EHRaCFvFViEqwgVdeqhEhDxqaKJr+nnia0uZyWAFQ0+3iyiaaigHrRVJv+QgbLFOA6LhxtpEXNK
3O9Tmj/PpMP/BDfoacJg5jRHU09eScC9Tv1qaujOsBjiwONwHAchh04+iKP6nnvqkhqKnrdTctRf
fRMTGsivt0uegecdizqzyihp7wFSLLnCm3JjjZ5TiFvItZjFSZUCDH8u0ywhqhLYuaaPn/uL9gp/
oCFdJpbmH3GWblTp79bs2lho1KFavFJ1S70suHKZyMHeRABcr6RbQodLRf6wvup2BCcvGSQDMROb
wsZNPy/r+STKJuCKrh3ZFyML4h60cVS/f5ZkEIDtCjgwsnU4IPrax9wT/piGlHy35l7hehLU3pQn
ZKSlyoCYeqXJV35EGGbMpcfJCCY8zBdY2GqxzZiSkJUtFNjWguj5dLiDGuqBqrFcs3C8vB0EOiGu
2GD/zhnqNMTUQzkNj+DhVJGatO3tetGAk84IjMgzdqWFfkK+0qzFJDUuTIJbgv06eOyfils82J1c
H9qXy2+3IgrfLFd8eEXkkPn7tUlqjFH8OyAI01KETzbIeUwWKdXSWNh6jiRfJgTshhyFt1bdGD2I
+iwRc9GQoV+aijGLKkfIp+6MJuuJLHtlg00z/MPaSvW7Rg0Sbj1WTxCsbUpeWWa1SDF6wcVqBSse
72qgzhz7HBhHnWpzwIlIL/a19Kq8wfzEshdG99kCUHjTNGeSh/o9Dzl1p8r8UTdsql71uDjg5QDH
ao9w4ZdVhLX5H/6Q5SpmPUrewIfliXMf7l6VOXTrWEcICKF/jwvF75vz8aKfSzTFHWx38TtTeGYq
tZy+hu160V7+CjnTaaM2U8L8QxsyiLPbR3sO9oTZicJPVr1qEAnoIcOpuAczex69MBTi/KG8s7MF
8DBv5jR8eEvLJmE6XAOhMO/CASaLVJuRKOwQm/obIEffNXvhak/uMoUHRAbQOT8NWEL3QopCoU6v
bk+gZhAPetxAI6Oj2UgfyZWDuuAO6m/JhnZydnJlOH3TdDf6/Pden89+zj4vn7HyyVRqGkVK2kGi
RvRXqVYNTy2tkxoSGqdZlVmhepHw9F4v2asUv9I5E+JUJXMlKfiHJIi/xyE78T9dEU+UxyABUa/Y
ycO9RmsS/HriNCq4D+d0NOf95ojyJcQi1MRJCIHHyFElK9XjMwsW+YBMccX/IILPIKAJl5KkKAYG
toxLmsrgOnK2puuoWsmPaNmJDe6IYVzTDd+WZiRT/8ydUgPzvTx3eNhI4JOBWTRr+yphgCAthG/d
TkbRPKcclp+gK37RFN/JnyBSYzH70rAL7wHy4QgDU9Dp8tBza3vgD/WsSULVUlnY3+OzrPj8ZFOZ
0taYaukh5DvbXzNGGaHTPOnTA+dDArVa7olRTvXEjn6m7sUge7+lvkd1+uPOkykn21nJAbIG4LPr
0g0yIkMD3pi3WA6pLBFPPTv3HfMG14d+gqSHwT/D5wrDimS77uxwAtXwODylHJTqNovVIOoVK65N
Tu4tBRefdRMvkdpOq9+2Nld7UiTN85VdInpRBaL0b84jsaHc1vPXr4LxuIUPzF52Breggj2CxAL4
1SuloaLUD0p41886Wf1ewk+o1H5YX+3m+NuoG1DFM3ENy7gE/fA68W0El4ZDbqXpjKEoVlX79RDY
avQxsMRJUlTQmsQKVRHWNzRqPPfKR4VF18voE9RGn8heDbvyk4S4vXo042a3Vi5a3HLS3U7/TLFW
lfI0K8m61Cvm+4bnu8KQldjG7NO91Cy7PWd8E4tQDwsDUAJQaQqVxmH+X8P8ySiEyNnoH0F6AsKD
43vYgyzdxaAv3rMbs0Szr4iHWfcFimzSYhUtt51o4fTl0TYlsV7RpT3OZ8xzDrvrHOCkZx6eTNbJ
u+dHC9InJRHbpPI6ky+PGRewL9UOcNxGrXyIwJ/4QEd3bHy32EnkVrdCLpBEvddfGVOIMKWUVIQd
L5Coz4VQiM4h1edu/Ugx7L2sj7JFl3gCfjnb84BrHaVQFKoOKulpgx5OG78ZWsjCT9ekY+Mr4DUH
k33GcFDysyidEo/u31yOOcFOLGy2PE8AFUNDKmKUY5mFhRz4FUHwr/XaD+cR/1aiqnG6a/d8Meey
GnXkSja7z8Sl4X9G639b/lfId5JJF3nHA0BrM+kcqHJxGEsmbVYUc6P0OjvONuidCz41p5ITSgAh
EyvbOFg7s8Sq4Ci8knAiM7GmxiYw+q3wJOcB7crUW1QSBRaX8qY2E67FjT/LwPTPTCmq2I89nvRq
z0Xp4BTa0Bw+vdMbss39p1zEpANY2UcO2XgXt/rz7S7f5i6UJvEGxTcXE01cchSxa6/X623MfgxN
bY9k/8OQ27530Wi416LbGgExXjgG/SOyU7GJho3bX9WsUtu/zvHHpBaAfpxXtl6YaXjj13ENWDBS
j470D7Ww3OV6aUtX7l+rN5J01kR2kd/t8uEOntwhTG08fcpiJqMjvIKbjWvjUWmuM90BArsJ1n8D
241DHUgLinVG4krrKeyX+x1AhMQ5X5lb9U/QnHnYQcz3GotFrvL7K7+AHRfRrg4eYOAMtLg/3lxg
ocXcvCQKIQB6tqQBrhO4BBCd/uozWqzpFDWuKGxwBROqftsoCAtwb0JZSTeK6/LOwNufbbj7cjMo
HSCg/QafO3YvZQnm/LkZoTAcZJdeu8HuQNOWR8FJLtoMLqTEKxZquGazqlUX96/Sbf3B4ewM4BUD
3sQsXtmyyJv7HgohkCdRVpQtS1Ejby6OhlpHSTFp/wQh/2C9qMRGupnThMcJPgJZdEEGj5j8xANq
ALfOpg/hgQRFeNOGUiwQfgkJVZ99L3bJTGJhx3d2bb3Ja8t1PCV5cBpu9zxVH25K9C4HBbaMxCFO
P+zCetLGAblU0QPkPHy2DEnz99OB3qBcPmhOyf/IxjEr03hdY+5l8KwJHwz9JN4oTV4I9ERomoOx
ELPMGR4+uw9W+kdaSo9LTeIJzGXEVRfQvG4gdXyLYVU3hxHgUOlizBySRyL+5quLh4lXaL3BCljY
gyx0azoFE4uZZTYiTgNLPn0lAsHBQ7ujhSnTVX7O21xdo6geZdFvd23RI9vIpCaQUVDkn/rbdLhh
oDGqHsOewsZ1WDMezgvyLBhTrHTR3+LM5nifjdgmZlGl+B9lW0RaFKNgOA2ve3nu9l9ns+crCv7z
uMOp+PZsD7MZP1+bpTD5aq+klz2o+TMpF0ftDOnCyQyZB/aRKHYu9pRYgG5CMASwK0lIEohri+Z/
AK5ePh5CaTWYZ/FVC+6W6f6wzTdQuw21lwtukmtWCckb/jKtmhOaj8ZdgzdoU/7zCGxCvzNOExgH
WthnTPAbCC/Yk+qT0LRzZ+WW0Hd5cRgEFsZBVWTSGjl+LwAONbivjmW//nLP9hZbJRkxlR/Q9VQv
/S7/cBNDmly+IkJnj/trizBcUqPiyyzb/2hqGNFHVlNcZjtlXR6D2SnOpYBws+7px/P57GAPA16L
pQfu/ewoirOCcvUy5hWgp2IFs7IoxKbzu/dhBLS1odIx/h18fgEI+/jcwS5FteAUPNmDkDrbrpQm
9Nl27T8RVYRVL/w4fLINe5rA2ompW05/zY6QMSs8gMfmBZ4zsPo+79tnsdIUenQVxSeL0FYn7KyK
JYXf5xiyYy6WiFdosf7MW9UpzbMnGg37GfcVT/AC+hMKI8zemENOhMecOT6AJeIMkM41eLE6fCyi
8pjWaogH5CyxINtmW2IVAQg03hYpiJPClsN+VmuEyEpe/4Cl/piDkYBHR4rNoP4Zzx9OfuKAjKre
SfxorDQP9VyVExxph1osMlAOVgBuhLYcZ9rhlB29OXYzH5At/Bv8IzaDkwbnE9iZatqrIzF/8Vbs
IsgqnnuuTKzJbgeQF2omlU2lqI7E3xS/BWwT5AMReDINXksYWqsa32NPBKLnMwIGAtVw3hpu6tlh
dEFv/6sGGdeVXlEeQoG6MGKUK9NSFzStccpDsjSfalG40RdErgBdcD0VSe5Q6hkNZbkD0OkapDmy
450ZpVwTsudFNIMnYmpI4Kxv1viI4IT94iIYj5DdFPalwJUTSgZ7KTiH3hLM62OBcZky3n/4bgQE
8mDuTVPJ1iEcrE0Pp4dsv+THWut1t4MS6qOoxk25jn6mMFDrhV2J8ZZlgkTv6f3CC/cm5tffBlxu
h0JeozZeGNR0FX3gLBQABxOWK0CajlEffvgbcmUFC+t08WOxjVAkmdQefRyjWTLpHhaOcrSNAe0c
Tu9O2Rdc/ZpNra8qe4RzczE47Z+S7ppyAP58g2ajAgXL1AT38R8wEXbZ0wVFiFEfXz5RBdbxpFBs
Q4nm378jZCToluOq7lOpaURARVlJuuxLypq1YhkWhA4UJeulQWnfikHTm1mUzgyKJTswJHX6BDDH
DtNgkeee+iGgaUFm6PEK5QtOq5csKlWtc/oebEx9ZOg2jG2DxoBFUi0J5KVE/8UEHSV35n56fe+R
rejY23JbLeJ1lficcPjNMp29oPR4vjV0zCcwV0KHOIa/bcUa4hRjGFu5+LliuzZ1uOOQEz4OjKHk
enpXhgMT+Scq2p4szSpSxi4bhWBkmigQaCF2r2esBl6wOJ5TeoiFCpr4XJZiLwmlauM+PlBOJoMO
jKCSmb/zPehnbq43k97CTT/fc46qjqIi4lqMeTaJSj44sEwx9YMF9b9oYSEkbGggtcVPcTAxmLEu
YWIb2dUd/MaPJvYaxLUd6cfD7RRWP07nFdBTM5GlwFKxLwEFVzpu+OMvZGkbyL+jFWmfEQUNAgnw
VZRgYf1CfdTv/7QhTqjOEFRqBB+ycAfH7+0VvGEvKimyX5QzmfJc9NMsq+ur/Gqlnzm3dcwxYJS6
LO1gs9YPl7+3TQDcunovi708WmpIkbJEohHZkB6QtGG6HxZ1Dh0zNv7Ot1d2JVZ0Wc02mVmr8Tph
TuL+gSrxOXnjV8xR5lQWtX0cwhmDL5U35h9pRwNuFhlE825LaGNaYM53Cuo72CXeLA2Pow44a1EE
2W089PY1CcIfWBdFXecOerGcJP5PihahAC6Zy0pRG4cwdL282g9+doPahx3hoZGnzzWi/nFYRJzs
kiaq8ycV8d7ChYWtu3pFeM+cVS5Z5G0u1cZBmR3mQQhAvwCq3CkHQE32iKFd8JyfarvnaSm7wRE/
jkWm1HyUxRwh75vPe+Dp02uOXq6+/4GRrPNS0HCa/uyITtoAfB6SgTtBvyFc2OSg0/uLwOwAMz18
5Y21hc0gmuB/jFQqbDrvxqORqw9zL47JYyEGDweYyA6Htrw5Hg6CmnmDWVwSi330x/llFO1NvpYL
vynbEEqpTCBWVeS576jR6/jcZ5yBNQTyF6nj6lAnRNWFsRux68G4rFZugzvz7HaCoaPg56Ap8Tjy
2vbbB7Uz33nvAeZfocobsIGkapy5U8dYRdLY8FmtdsDDoj5jOPOSIJZy1Zve060rPQQ67vI1scmZ
7nxlecWYKdHiqBDei3XA2hUV8scolyaGVgDA0pzCkSA2eytqxz4FUGujEL73u/fhVK8htwgUr5WA
FcO37eMV2ff3aXBWD7UWjTHKiO9jLz+5kH6nOTqAhTJi1EaSDoxihfs8bUeCWOTmQX42VPggc5us
i9exLLWFtkR0zj2x3fF60WSWKIjIdfd1dJqsU0SsnXwcLRoqfuoq7SSGM5Ksy23d/CA37vr1oJYI
Zx6BIgzbtmSqO+3ZiPlnUsjYSTZMVNysKftL489gT2iRd/tUgAmYFUbgzBpynUl7aHRkQkrzN7aU
0jJYlbfP3wNbtmEDMp82zSzSB/C04Tm6aS97MkXfyLHfKlqO4EiKHizduMVzfJHFewjpmSStjqyl
JyazL0om5O50vaKCVrehTHlx85cmYVfpRg8ojF6FoOqqxbRIiA+UWWkyNdhk9dATaEpOoTiUD/jE
AUY3nbJk93ciseo0u/jtXaHJNI1uUlA1H+iGbGLJrWrY0kib8JF+/JjGjVSwfzkB7y/KOZSXZk9X
BcB0/SQW7p51CyEM0iwyNpZbfCCRxfoakVHws+HQ1E5Je7AoJbCVecOB11rHjVnOswNIHlPK7ZGu
W6JD3OHgqyfxNBVG6moLs3AodXCzYC074mD07u5C2j/Q6DvACmf5pXt1V5D5mi/8wezv/KRW0JMt
D0sCJDQPGxHqDlZLSdtKfzlqQJnJ6YgpmURwvoq9cpn6aer9/DMi6aKEyCCGwj3kqY4XHcY3v2Vk
7Kr7jqmxz7Mj3IoGqHhNHE5SfvXwkBBRpeqmO9RIlRJhV6zgJqTkxcGw7X0Hc+P995MuIHcbRm5p
zBWAexaIcImPEQIDk7qttMPbBYVNqhguRPQ9TlhET5qFUGJ5lLIdhrHKGuP06CKkmYUklRrlTGXC
vs1DDFlkR3yRLtOXaKzI9Nl8bW/GCW8+sROmk28RS9rR+AbQS284YOv2/ldLZTKfmHCnMlyFtvtb
7M3ykoJ1tJA4k2ha0nH9KpXRR8tvqSL6hsAg4Il/Li0ajrZtV/3dttExqooNMGFxhJqOtLgs+SZg
h4fR8ySFB8jQOzzVtDpZV/go5q5QFLVczgQRrfB/h5LxPB/wIT9ymzsTmnWSy05bqNDKgzMX8ETL
/gM0e37K1f1hW8efINepxuUsjPHZDRPkrXvTFuch4k002Xh7+vQNvNzQP8H3U3qGxlpAkIUIov8r
oZZiWQvW3gPk5bl4NHTQ0+ubdLNmqXJ58FmmgG+s83Y4BtXQacpmLz6uoYlCJ+7NkHiLFWPP7Fck
ndxByGexvi5R62FvX0EPTTPOuqjgcahdb9d7xn8BIpdW8sddu6QSDGVHMYvopehVAKroZ6UbRXZ8
3GYQi97ZOli4udSfh+n2Xe0pr/vjbTP7ZhvJamjjP6IcErYcyR2RkekKXwes168B6sFw669fc9AP
gUDsg39FcEnSLy9vxw1PV9Oed2jo67sE53xUNpIBBsAdaqP1BiAD6pzwHWLTY0kJzvnzZa33Yl9+
ATSyzwRsUvtwVjP+NCZfEbGav1O9jnwRDRyXMwjj5owrChkaikBlqzIC/vhuHvnHc4rkJrLfNEbU
uIwrjZkEqRDw4ZT03kZ7Xth3yf6ylf9n1jfWWKzWkr+SHGRu72MvIzMFiaWDS4R9y2prSjepeFrX
epFJHiEF/linYjSQl0PwNz8QaNyXcEaKOATBjX3XBIBQArTnREnW0V8zMsQaAAjDnX+rJulk3s0k
7BRs5CnMRJJXWT2Kx0ct5E0L/3YWMwl+2X28fBnzc9KdQ4fSw0bduFF7xFAYehlse+oq0z7bIyQI
Agn9vS+IHx1Kchu6+4mwPNuv23juaQLvn5ueOxqnfUFyhHAKXP6PXqHJLUwXjT/mfNHct6MbmtFD
Yg84gNX7ldA7DlIuRLCPpsKpcCKLON2p2FN4Hs0Ju0amK3h45heTs6FpMWQ3IM1Xx4ti2mOIr7yT
4T5jUCT+HwC+6eWia54oX+zUE5r9VQVba4PQws7OE0mP8QA38objpWvYEzNm121RcbdsADWdaGXW
y5ejn8b9BveBgiOIQqhyZZ6CYpmUJuJ48j9s9JD3XQldDShhWHB1BNcbeorqNLYembEFXbUmdgol
6LRopoY7Wtey2bjw54CKlROGYGy3f8zlsPpeYxR+AOOtH2+j+dKrk083c/7I57J8Q1pVKUsS605g
3yWBeO0RlUaObHOX2g3nU/Hdh0HbVCqISVWQA+ywBDfB4n76NUD5TUx98jLzn4JWqNI2/+AWeXTC
4wZrRea7jtEFzQlm5spAd3+wIsrrU4AkxQyTjg9CmMPF2x7Zk5+DIPbThdqEagZCuYHdDZ2+og/x
BYLCfOjrUaYgXe3kVZeOjz1ImaDsAcURUPMdEkUb4s/e8hkyX9QV17H9mJ5JZ1WtuI2NoYK0xlPI
AapnUT1YJDdnSRIIfurGjUuwAO4Lie20CHjq2sU8bCHjKpUDUwrUsknCvGNNYaSXPL80boZbCJIC
hOBumahmhMx4/sW3OHJoj0RxS/YyDO6w30XT2RL2Zk3z090sqLAcIZ2Xen3s0cEjEgDldegsIC4w
R9KWHTvFa5FLIH0EjkUHMa8uX3fgkVTF/jep847f5JMuFKPLO7YSsBEpEJEUDJqKfACOs55YbFMG
RO2m3IDoGOIxeb0jZ9PHE250AXIXNnmCSV4WVLI0sWWUx+gf+uQf0Q3ZLU6HEImBO4DrkHbhIfXJ
wUG9wolWqS0oa0oeopKA06POyVlLWBnJCLfrJn5ih6tpMoPP8/fCdQktMOepuzt/fPeAr8XOMnkX
7brN2L18IqxpmaM3Hb2Qfl4iJ2/fMsv88CHdYmO9quHR08VauMjOdgqmC2nayN2sn94/7DqT+AoC
ZHDHUvQ74rtljC90qlx9c4gi8h0ZmUzAQm+4fQ11Nd7CucjOyvuaQevZ2Fp1iv722WqV01xWyLqp
rcgnZ14eBky8dKe61Dol3FWLmQToZdQS1BF52o/Pwl1RoTEfLmSY5Rnzpy22QLoPFw8NmTbW7Mkz
lyD7F5moO2lwmYzZ2WUe5qCfW5LMh8hfDoDTeozgmd3RM6X6Zzp5fuD+3h/y83S2xrnvvvufpahh
CgePWzR1qWC64TMBKh+OR95NU694dcEB350w9oBDPD/QpPgV299GFCo/eWKKVJkct6ywiVnSOQVa
LZEXkwusq9lAquYQGbsL0ciJ9kLJbIAqg/uVf0gRNOjnhPjYTmE1odICJwhzsBVZbquZwqKFnaaI
fQoPc6rdBf2FgjD13cfDtRDThbkJO8sBO8WljlwXCYtuDNV4uTSoevGTueQawH71CN4Exr07eFOM
/aORk/hQNR6gl3ocsbUAiCtxEQrvgR8hy44mWdklyfSkfSk1wkwXFQ3SXGUPEfdOXiNlTHhS3Rpw
vEY51lt6hfPcKOLeAv5sj7f8fewDXaFzSkkz/j86NgCMuucDj0mWngWChtW4WzFHMZ5kBv0/T6UH
dAjeT6pf/JCYCV94+aJzhboSF5tprwjvuJc9ZVYpeFDmJ/bZokZD3ivatGsqA/eVOX03tAMglKn0
uG0GLiFtrW3ZZAhL8UdaiOwGdOS+V4Np8XhCd/MKpF7FyGf04GPWuTKV2QWMo/UJnu98jwV5JiAM
r2ztfg/TP+6AAFFgSnwtUhbQIJbVhgxf/tGdBr0mgT+7LBA3+hzK2oF8Ay+rl2bYDqWKy9EbxiKG
uGgAOjbOR7P4u75UhdhUv1KDAj8QLGlwZnnp+296bYsKvMvdY6/7BgcY/Akicga0as20aTGbmuJT
GB5aXT6WFy6OFAWQYjbz+B87w65c4x9xOyGUDrhm/ueG0kNwHEO5u6BJhMC6mEYr72PyFJAYTR11
JL/+kJG9bYOlqtVvbffM4h6St746PLeVv4rOtQV/Ssj7vyucdh59OK2/PLvzK4xo8ajbhsiKyz+w
e752L83kENRlX1ulSWmBlSKp2R7cMy57eyT6aS0AOTAw57KRqHFFBhS0y5Go0G4xIh9CZXGGcLcV
0HUvmSdOdIhOiMGw6ElWfgPMmQBMdslrMVY9rmpcjx4kvU/yvNni30h2oabPQkT+sau08EVCN3Y0
+F7MoqDUUz6CU6I9/K3CiqKjqUPQF7Z+X34CsJmz0SN8f7HqnOA5a+TFaJRtd0YG8QicOsVuUx5M
xHqbKLygWEzW1oBTXPOKHhcSZzPjNjGPH6hRLvjJxiXJAN4GsuWqRHXlBSzd3AHLhdzkiPpRGDwt
S5FFVe0h4Uo5BjU3gkCwxLhUloQAWq/wArnMYnrdfl5YFZKjv6xrmujTiDj33lAYKHjSzDdyrC9i
291xI7WnGbpDfYBdCqIN4JlMJ0RHkn55Q91vOCz5gex5Ede3nPG8ohz1cSdb0qb1sPckti2K7t8e
mrzkmgBg4Pd426l85EV6JkNZfH4FPvGT4Fucm3cSZg+w1GMBh9xLtVTwCfyrlNWMUG6+To7LDlv/
vRqoDjKcYtL9r+2grFY6pIOYNxxiuVAjuvYbOJbc4bnOaw9taEeUCyHDDzeKtgKyy/mVP7P3rojl
Alri1gms/toKnzsmyaalMcJ8RKGBaPHNJ3W28rMM14+9WzoGSIyEEB5J/PH7RiH4QSRwl2qROPrW
1o2KvwViGJaOIK/AK1kCYoaPkFH/pyUGERNsoSQIAH3V86X1F4AqmAzzQ7ikwpbzmRrfeVvgSHG9
gdDjM+blMtJg8P7x0QsCbQAYoDYc+oSVpfuRtmCosHSnNIqvQQVmQ1p4QXfmcbEtiphnrRv2LELq
mvUAaRULU1692lXTWje31OBVdp2P2LOioE15U7AWLVWghVI/tJQMHMeLA8ZJw9oKZuSqWop+5WWT
gDyfARyxzeHEHmKx0y6YB+WkPqyEWX9R6vdew2UrCIOU1FovTY7CrO9GDYfsnJ3e1Mvsw4GL8aew
JuRo7t5ug8RY+22uz1XTKVNe5pI0mku5e113BVhqA6KKIh7/Ep7pwROuUWacSL3D2mydNqZ5fSKC
gmeDWdIFEftH/DUxb7KcC/bXDpW06z68IKImvUHdxRLeVoloLaC79FAL60PH35V/WdIIeRvkKatw
cVejQJnYaYtGJKd+9bE0GfYrkBOKYhFcLmCpuvEZ2PvPrqlIOlHKMOe8I1OFybtgp4yjAPTqOTBU
v3+ksnH1gFxP6uwEQaHgLK+DfKwJP2BzFJ04nlwLa9yJSEb205i5MFH4kZZGcySokUoIb5IYH3WI
RbyW9CbPS9HCChKAGYTpCeDQKjK+0hFyN6OOBOy34FzxkD6kPpzA5g5Ek5RitZ+fvdXhaAjdIcLo
kB4gpk81hucf6N+7NnW8aYrQ9S0aTrMWk0JEU90/ZluDVrK9C7BHj1B7oXB87TRHNOBxw0MQk4Sp
EAGBCdNb/QanV4P/ffNfjc80J1nSUYGHm2MaRyQqa/ifXMSUdiwQr7Q6XqwSwyKdfuNHLXIV20o2
G+G5pufOKvPShJ/oTsSZTyaqVvhNaIVuI5UBvYed6SW2zUQwsMhWhpqeDszvP63j5mRJrBwM++EO
6evSKt1+TzLpF432YQCr1nY+oGZZ7n/eoO9M/F7+gFwpq7/PmCYlZBM0u0LCRWBPv7/RYwMxFJhK
Z+z0/xKw1h2kqvM2PmKtfm3dXWAmUHE/JYisTY4K6nGoBwyrsk5jQN18lRl5QWUQ+0lABeHLbJGz
zZ/QfMKGHIuTmG/NVT0rBopzQE1wxyjDpMM1VZdGYVXccGTKOS+HWuSvsHZOdYL0CR3cRrXl6xu5
3j1YjiQJMZliYCsjW9ETejEFJKffJpx6H2Pe0oZ5BKuOQxJFgFX/Mp/NwveBFuyYNg46vJHmr387
zrO/sEGvs6fwaUs63E1Ch/TCaSKJigToTxI8xThVuQaVN7Cu6o919bEgMzHvtxSZpK673xcrdtxf
d+/Tvx3YRTy7ZzLBhAxNzrJKaL/vPCr3xtSePH4SS1rQHTTcs7RhcJt23UQi+bbVp+sPUu5UvMTX
98ufCxqDT5TPmXtIXJLXo1fp3cYQeR5CF06YPBt5mryeuFw/VxvyzNbH4V6iKc4EwtLXvOnYnUjn
RiOGhJ0Vjmpr3mlVKxn7xMXNaTu7Qhd6ye+d3DLlez1jfQBdul/69PdkCSX4ra+5IcMJbFzE88b8
YP/FRT077AeVDbFFc87mvwLZC9MV8Z+ul6UenSQ0nilqJbHYydXKuvTnSu6fGkLMmF4lpGkz7zwl
mnP2yKM26Ad0gRPNMn3wzP0mRSL9Tc16Qbq99iufwyIqdm2lUYt8/VR1OQT5h+PEx+UUSSHf5TCb
JXmuLKVb2QNsyMSaqbKMtA0GZM3yx3zdhx+orajX18ckz+Y6IWK946JkPHEYlL4O2oiXP3O9BWek
9w6SkGzwYYcJYp6OaqxwwOlm3v1QZv0R7736Iw4Zuy/W1Rzj2kf+hF5ms9WK9ayUrQ48g5GDU5/f
dL/v7TXR6bH2ZrDw2CAQd+ZjPSX9GKN/V11ceXXjZHtKyU9gonISSogWAHNIH6NEgMvKKtucBksM
/VXlt9M3YSymqV/lLQI61We2TDZpxATuGVDIa0e2k6chNTuln2Y0FivEeWNvdSC4EfHJvvo5+vM3
8SwmeXKbwfdGsmHrwmDM9mfFy5G93Y9uppDuWxGYt/+lBwcG+o3+ZhdHVIQZ9ufvYo/ukP7FsPBu
JZFR1iCsAdh9sXMuRUcRgh2bJm5rz5sMHvwMD6Mf/R3W4JCqDqTHUBzjoI5nqYiJ5NLZEQ1RQIC4
VnEbaArceQeFTvAtvWDbFARMdAXhXghMhZ+uGiAd5r13q3noGaGk7+NGAi5p2bROpKsHLB5snhJF
3ceMg46I7jzJX2CJfJgoc+CwLwFZhsy/IqJrpeqeE5i6gS2hkE5xdttbiQo7FlV5cunNPGP/ZGFW
rbpfp3yQiQegextFYvOJgjsCQMGEgcn02SyFR2IFP6iGx+Zk35W4vmxTygjFmNeK9Y1mT84ADUoK
HO+P/1G/S6qyyJ3822DwwRJhSPJP976Gq8wC4kulEa5iIE/zJ8X77j4lRp8Y1xDMcyPzRSOkx29a
eIUC/yfsT921sHm/00BuS7aWl0h2SY1tCOjqPYIfqbB39zxuPXkKVwzWTRNr2n5swSfshxtvnjBc
5MVGHWFXy4X5p4yKhDxh2vofACGB34XgnaUgsoeGV+Uc/6ZvHu7W6gs8pj1Sd8pwDt5yuDZXbrrF
zTD4o1udrBR+8r+rSZ3YMlcq4vd71ikC4pbjaG5jQlwwVLWmyg3mPAWJBfTdudgR8IF/mRbvrLpc
7yPlNnUXrcEODtnF1G6n3fF3CD04wJjX107888S1sbruvr9uBjxrGFbQhe0VcLiNVTdGElBtAPc9
Y25gbFA7+YJj9G1ENiSCxtciHmAqRAelz/+X5egI48ozK3ea+41ZqfG+EBpWGK1n3/jdYftG3HAq
SD8MN67tZ0g8zvomjXt+EPsFOtUeKTgNMHHZQu7AHTMSOPPdixai8E5I/fisgKMFEFKfhMfjrigq
VaFSEl1Gg6rEwBq4og8z1kqGRD1niON5qGso9RPo8axhgueZ/NsteXdycEOAJCv/a9utb4q6NMiy
CtJFwOjpoK1nrNZMu7iETEyd7D145eKiNMBcAUnSCMn1X08EXNHQOpd15eWHINHBe998AJU0r3zk
dhFvo1BYLjjGRtTUUe71Ycx6gJyMFSr8pVVqDU4oRrjOuoNHBBPannIbN+CoawsX1lKagCOL8kBJ
hxNjEcq13hZHYmKStdrtoC/vArpMBWGQ45MiBBalUZoaJ0Nn/ktQUwn2Yvo9P2WmHBa+NxwN4bDe
7wl1aJorcBmklGynaYvsNIS8kBeYTCybrTtIJ2a1Q1V+luFUZi5CTOWnQTMQC3b3+LK8SQQEiHwk
4IZuAVuSaAmVDwpuy8eyBatOL2sRiZfQwWgiwKulBajCZYyr6oWINj2SlgiAlukUOK2DxB3YD+2j
W484pkt5DVbberGCulY8ySS77qhNtGsDzzyVzGsNr0AK49XhZlObOK1LCLXKkLSFk7mAcjjg9pcG
m5Sf7R+HmP8lnphwjX6Vl3Dpxei0IIQWGqAzx95y6ats0Wc1S2XMj8AE0PnBd8GuJEDT5Un1S8HG
IcCIOGruR320qLhdbVFED+WN+GP82yiu2w16tr/wzeyhjycIXPDs+VPfMWddoRHxx1TH2I/reE5m
taqJ/2UhOVBhYf5Pj73iVdOmS6HezUPBkur1bNuMRlF4MX5yO3/XM31CbVntUBWJQntdXMhq5W14
hi/dklhA72yiz/FAyAz85qdwhTYTMrlErfTjazz/qZluYVjRm3evkanW/N2cConkUA7W67pC/4XY
iUOzEB64rSMHSkO7WKQJ6KUf6spFm5yF+n/MQz18tWwFjwonJpRoEOuneng1BU3fbHhYMxkDgmfs
2dBQZZxCk4zQuqfMDRg+6WRP1ZpDKgMje542Ms5/NHFlRQn6s0Bb9db3k/Egnna6qZgOdhqnFcYj
1bgk3KLDcej3sKAqjeKLEfZY1aCIVjGhPHgvLNpeO5xiQa/6gGidD1TfKoIL70+dMC9GCENWBJJ7
jT88Nk2CC/D422NyiCb3uFVhqVTh31LWPlxMa1igUmxoq2lL6Vnfd4bjeqexYltsBctqCiiSNVeL
8P8u8h1yMLEmLi52LhwuXXzFzL2p07cNeXbhDz9tgOfAjHJAMM2A+UlTTDNDif8i2rnJ0UdyMBfY
symHqkxdYbFBq33p9Q7nUg7DgnNyJENs/xGbQMIeb7Uv41Az9FsAhdS3z1qa3aklrBjPSghMc2gy
qj9JPoqTwsGtBCuRacaLmx94N5MqIWOpKepF9t8t/TWV7n8CYIwyiWk2XJJd4cXN44S+8V4f5YHh
6hJ4OJmpv1/VlA7GcMPB/DkAsHqTrC2Ry7DYw3aEiKfeboqfnhMk9G4i+pcKw14jIU+MjHYkyjXj
JmCaoLwNmB0POlGNjK1RDcNP49CURDCoOlqiRkOq5KnVK5DBsnkMt6YPP0BsHYC4/xswv0FlSJT3
/BpownTYFGziJ0p9ovR+1rWTPG0wKmEVItzyyJ6zK3o6hTWc+WYXHXeWNLkShmykSi3G1NUHkFYw
edwjOwHKOjo+L+dIn3JoDU3RXA8lTPo6iJDOyIZLwVl45qXf1rZrU1yMBzKUIsOLEkAkltAczLzG
bmw0DBfpBhxeOHfGczYuwwrF3LC517SFZgPTIZPUkBGejo2htlvh7SVk7PkK7w8NBaVFs5riCWY8
pb2/EC+MkXNIUswuK928TF7Wxq6HLBqLJ6P9X5UyXLvE7rf4HbYPrxF6bWH19Bbx7rnQaEk/LB1F
nsYHw4WjCMApdUsuWTUmBTuONK3cNCTgdD5YgVv9yap0xK2O4Z3WLbrdAbq4QU02IapTmWbrqZ/M
9hs6dtrC7FTki2bLHB/WBZRE6FBLF2L063Wmm7nXW6gFer5MoHX7hlYNrqOce/KoALv7YgkxHsw3
bqatSLR4OxXvYZCHm0ZwYw0N899ORPVZO15eJOSF8+ONL/Q2AVTU8lYRNBggfEgd5YkgzBUfwHYU
m/Q2esSVI2uY0I2kxcv9e9J8KIxBTw5XNv7uiYHN2CZsY26Kx7A5yOPuK4GrQSHI6DCcvfk8qiR3
O2vkISp4DKrV76pVUobWKCKdRVoDi119Pt4w3TKDdxc2eKFt3zflkn9DvBeGKUa9khw6SlUnl47V
CrDHMZizJl65RyIMgurMgHKJZX2TADqnLBrfonChKn1ZKHtMlRlvEaUkUyKV6KsUlGPlYAaRxg3K
ZVIBmhBwy+DCrSWPcFOtti/rg+1i5fSKvkM7lyOf4Q8bcsZOH7cKesCX0D++j4Vjpq0ZpXMQkjyY
G9fASFVtoTuQwXUtLxHq5A83Lb21vcPHzYqhms6yunEF/9Duu6coNEMx8r7vEhq4e+dCqZEEWd40
FZoarvtqJz9rzS/8l0EaLPzkar5mFezU3uSTusM5sRGvoaNb9XcX1HnQ+rL18dYhqI6hKppRYTqB
L7DtkYiFVPz9Nt//WfBtQ9OdwX6t1yWlBAMfqsV6NHUGKTnQYGVkEV6XxdHhSa6O0BeK/O1celmT
tZELN0Gn2Kp/jm4Fm9j32uWqc5CqV3oeISNXfLDR9o4m70WzyMqMa46uebheMXOndFWlJC8NYe5F
QC6tgznjeLYKZs1Hmyx23Yh8tA8SgipB6ASk2++pEbQXYN0SYy5epRrzpZYIHrfFFb4EjNbs5gNS
Xu9R/aeF+kEM49KJBTtRLydrStiF2Si1IjNfPF88t46bakGUktuCxNLYbcRSIjH+bFMfprI6fjRB
V7FMdtefnjtEGkh0YOOwgjZhr4WWAp7FmMvgDvqbfCCtvKVnghTW3HFfPIylxcm+3VwpoaHs+m75
XHybL8HmCjZ7FnYSCFUzeDazJ/gsZSWlTz7+eC3Vky2IU/U9W7EiRhdjdQWU/Dq5+o1ZNGbT/bXy
BrpU8PorXXYco3i5i0T7W0T18EZRTBvxf4YBdzgMdgN9rYWhm9eglNj6dn1jSYBIKwBv51UjsUKn
AAmbXzfrST5h9TkhBH+Ba7FgOUD38RaA2B60yCshwYU6iY6LxINoYzbNnIFsnulD8DK81ib7FVKx
KhWgp4vNg0eB3sQKqCaLT3levMZLGSnxxFNclob9Hu1si6jdGn5+4uhbwDAQQhE2zhWTArPavDD+
guPR3LQ0iPtsMHaktZ7lQbK0TvTVvh8XkkzpNIIlh/G8IhgSXBW7P+uCPqBQmXaJLyvAbBlpygbB
onVENRFi+FChz8Yqi2tM9cr/lqqZrpyMUYoBVUFpEe0e6M7HrWsRdGhcF4dYiQmMbvcBA6uW3aVI
XrHse/oxB9dM9a+UgLES2pkHTisudIsnjTwc6HI3oe9LWp1Yw5jmjpsbhIEnUHzk5YYS6DKV+QcM
EdktX1f2reS7hMSGKuDta8GVoLzEmB21MomNGKnd0ayAQ4pnTjv+DIpT2oEm/AkKoOqeayEXoqmF
FRlWzNZ89z9+cCz5TjejY0DLLN9Wh7s7aEnNzdxZOGNDIlDtnxEzstR4klcBQbXq/DvAZ0hPHbKh
ByuIrpw43G5/L3KPwWFxZD6Q8mtpCIuFBRJ8EeHDIV3eKWIvmy9rxXqG8DszOysysURfQ+ZYlZAP
Uv507kSW1qH/E2LtlLILzXmBbl6Ng7PY3+10bRcpyiEoA9pm3ChqYUNVg9gkYeSdqV7rDpzSjTdY
hp91BNF0HWhf0oR+MLZgc91Z864xeUGtcgzxC3Pls4u0s+e4Jv2FmqP4ze6gzXD4mWaMTK1k3Dal
031q2eirtUk3GyT15GDdBNYuDfZnmU0lcysPCImoIOeUSTscYNr8pPLXGJLPe0HbBgpk1c5UGsqz
4v8QuSaRSyrLplOKziADLDf2FVrQQIz1rDTFMFpd9SjFSMZq3+r/2Bb3gUDSVGtINM+L33rVXoq6
VLaYuSU3jU/EKLmC1GLYrejkLwe21i8RJbnBkOshwilCY5ScTsMgtEdPH13GB1xJIlovO3atliT+
rTbQwWR/pYuWCEwcyZUn1s0rkg6ygN4ePMY0ti/TgQEiFSAVA3IJeQJi99kQWQvQ7BBknndVi4xG
VrRJnrgy+cqnLZE60FGOIxHw1KRpzfyvvWlsn5o4L9WZLYywzwqvgHf79JqeU29N5EXzg4pJMEt2
Z5yG61WtVmIAq4yWkxrRUU30obngAziSmdq6iVMR7pW4am1fEj5sXwdiHUY5EXcNRptC6NUAe3R5
yBUMs2sIhvJfq2nyJbAz+Rx60wvkI4U/aXnZYFAp81fxt9Uz/FJZC62g54xThciR7MTFVjDcW1U5
jSfVqtfnpQ+DOqMAfyHTnZctkiQuH2LF61T2J891izaOeISpB8uuIDv61z3vTsQFmJHT6zuAyPTF
ycH0Ah1dGh9VD8Sg6J8FSDB0Oz6wyKWk0VkpZr/uiSmEbRMJR3QHHy2Eqh0KlnIfhjxmYKFBOCpq
OgVctFlFJrmR+UiRm/gZxqmZCx30kdoBGAY1Iv4ZdizdY9KvsxASk1yl5YvhDv3a9RUn6UPExLZu
UGh0FeV2E1CM9HRoQpI5bLxImaJSUQ5V1Fqn45fhKGV71H298PlfJxbPGGyp4fvSX1eSRsj94k4+
f+KB9H7Dwp7rWumbNh5Wujt6+bYchSi/BaMBzKvnuqi0JUXMRO5MmuV1i/kvXxQxkKeBqT3QGmmP
y6LUiJaCHb9t8srllQ4vScC20ftxuoGzc2tpz6q+j8zeot7TmHVbI5DIhO2xepPke4vnndYkkI22
lmYJg3Vo/9SltY9sHFVYZlHhWewoyuMJK68HBz9fgm1woCTM5s8sKz162UVczujjmN0nMgDt7rtB
FHcMjGkh6LbsCihqkydqFpWI0t6D7YIJimsh3oc7QlqKTCTxJY3ArASLTODQzENXbXce7VqpFFZD
R6jfCfBlNMBxLehU3KiumBYiTdyyRk/RjoQyQTbzzM3lTH6kxmFspqI9v8RTFOtH/Tz6aT8YtyWs
PYFAbWGpij//PZBkFwHpKYnN3d7UQp1+aJivFS3HwKqEJ/7h9p0/Uk/qalYSR1knY7gyBjEwuGTN
EIAsELdsp36EizLph7jmoYODuIUZm3rHq5jAUTiBabn+OUbLYn9ZgcOkirfSHuXVYPtoSln55+i5
/7GIAu6Hp2StZYdWy1Qj+Fql5AG5hCQRYnx5gKbBsQgvYvmGrgmeKBly21lyQJXeU9g5zEew/GMs
rFHAIZvSWN+L2pZ7fAJU+ozCQ0GO1MeQG7OKEfoclh+rCQ7FQ0jfa1AiGiV9cJA6FY1tpCs2H+bY
dJKkibdGRxu7FIrvrmqlv11nHlHBv3um8lE1lpxEC/RnsLyQx0lWStiiXLujqXjihaJVWnXHq4tj
FhZYSsxWeV0EiolN4mVQkG8Bo2U1r461xXB0zl4UBNLPuifqIqswUrFiNvyjje2G7ekpfO2m7rRm
NuiHXbl8O/WPqtyE7ajzsWdcPj8gjvktkks+47cPQPsjENX3JPAxVMfzriyInCMnEthO2BPJdnPa
eCzfzV0JLZxiIH6dG9MNBczPDXxgKZKR1xM/cn0PBSyY8U8Ac9s/PQzVslJ8HRGQYnC1gUshPU9R
iljFE+7uV67AfQviIwIY2RdXQzDPc0OWd4l99RZRhCtoUjx739RXc6xuONNbtxXs7F43gKmxYMTu
q2MF/MkSpDKwlCNTh/YVk8uZOq8bJ2gaAyOkUrdFhVxDUsoEjBXZTN393vdAmVeu+TyyRaEnFQV0
EVt5wi8kGmB3FMYWHfcsOq8xIRh4yXGoqFcum26a3uosrs47HwM8FuiOMm8GsXW3/wGLdRCyt2dQ
YNmFzO7j/Cjafm3inpnpwh7ZO9HLsqCSvmBjOv4D1C27cHAehCVzE6stxPJetpgDn80BV59WT0da
f3b/nFARJtdAs/mxhjSONI8GSYb3CxdvzJkIDA4xdwVIGrd04PR3vhpiGWAcsVlbs02lTvq3muDd
XcAEqlN47MHSa4XmTiebogSo+xHuvSFZcJOGysygkdSFNhpTTQNcvfRnbHgMWbT6IR7RpSMO+cH7
dgjmHtYSk7MOOkbM4hpY9xyyM0gIkgnr2lho7v2ZKu0ONHhqsgcki5rONJvjioewsgCJuVnrGVRq
d0knhnZSqLpiQWrI3PweiKwY7i6XVQmeSFgTC6wY2Cl1sZAo03ep+k8tTthlsmvYIb0u8j4KTLSX
XNPMQUIx89miNOE8c7uZOKfLChGT4GputMPdbNS18FMM/VFzrcbk/8seikX78U3t0RsG3nZvkjXY
grKE9dxzgB29GoSwGT8tqfkUs6v8Mvmfca1dQslJKGPboH0VljQHa59mY077fK0BM56b3IqDIFRY
hgYPi03dI3oi/jb9to8NJoIrTo+vibbxApXJiK5pu1iYz7k7HC4/FoEZrSAZmkNXVHPfpDG4psIb
6LXgIWDsMJjxbtQzj2KGNMJ1xb3YXnja/Uf6ml7lb2qwQH0JqVZQEA66An70RK/sVHKOEtwlPAqt
1P0lKS4pakfd6sPQbgOP8MkTazXHTm+I7LQhS3XVf/CaeYHbuJf6kQjuE3Zw2uIqqjfIM2x5r0Wo
/4KipVqLbcAX2UCoev8OMOcICk1g5APs9400DMSxjoYPXysVsJl7REon4nI9LC6ZdRyPSIdMkYGy
cgIjsSWQLZDTh5V5pZW+nTqVJZhzuEccyMYkALJyHvNeu6touRPhrUZsE1SWo3XDSJNH3L23kzeS
xLSSUgk883OWo2iVMEguf8ko87JrPAKSqyNxXX2UIyyLsPoXoPueL0YlP0m7PrdqxkxmEKnVwUEZ
7DVefNrqmNyvGald4aRJg0NCuWgUB+vH307oFW96P2r0yIiSw/AfAG8CE9NaNezP03xBMyCAxXXW
wbZ65rW7LosNUp5g3gMtHey83uOEkEVlmCZ2NZ1KnWdRF6AV3VzH1N5RCfcS6HVuNO9UhVv+nntJ
h+mTfQ6HFTlWWOgLtY+1HYlWFUQNGVEXHi2W6Bsp8rmH11PakWHBmjTOLdpdjQgA7USLXp69VopJ
k/mlZ95/FGp6TM+XD/TFUDJ2euJ3M1p4wuURlHp4N2C5385q+B+zAbRj8cpejv+a0uMrg44pbEHR
2HLXHMr5o3NN7tTCinO/hyo2cpD+NMrSrzxOwPioDVYxnXB0F5pUIqCyuK38P6ExizSHM5bfbXow
LBqGNtvvdTGAN/GKOV/jU0nNtMIaXrTdtWFoTlFYKONwF55YfXz0Y/+lORXRNy4oP834AaPpBi9Z
ahWplqxkhKG5sq6qFcjdBwZGKWg46C+FcXIjMYEmCTCoDz0us8fxKpuuLDyKo9dMeW77WW9b3kVQ
LGIKA2Dx1lCC9fUWL9nbYApmzTs9dv0YK98K85PfwwVkxBMTWixEC/BaawKiJDcHuDEWqIm/1lL5
r/lT6hpXBqIOXHBxDA7acdEhvYw/uGnZlbQvyoe3eCmpJib/XqXJ4RhZL0h7eHm9d9A6mdzX3Qsd
Gzulnep8OWpUR6Dyz6demWEDaKW5UorBnYGcwXbR2Z7BD7BjtcNIlDg31n4oA7NCSuEkusEjnpwZ
ZwBA3xrjx1DTGtJGMwSaaVtVXnWNUqBjPcMcI7DaTM7n4MUnLviyyuP81XzCQ24ngHAs23A+Yqzf
k5v5ZEk7BuOfBa7nBxYtdWrznc9Lkfs0xnvKTmD2eKmclsKlwMg1OHlCpCY5ibiPIq8t3ytged+F
5ssGY1grTKw5SUUZTiQUZO2WEZLRODEupVnM0olGq1FJlYz7hFN8NMTFsHcveNMJ1UawIG9DS9Hb
y+lETDlUNvnKkCrPkDaf+JHXdZ9Fu7PzJZhnsPIxkZNYUdiAD76gxC1Y4zuDm4UheBSOgVfbuGbB
GeeyHm5qiZqpQUmoSYgoeJ7XdUHGL3YghItUiNJQxoQuhuDGFCX0ZSxyKdHDpi5w+dXGd2zot/r9
IAuAJ01bVea+QmN+Qifjs+GwWoc+/OcYXHX/wTj71RXgN7//Tb7+5DnqB3H03Vr6xq8yof9oB6y4
FnhSqvJfvA+A2NanUY1etsTLGbT1bvdSmOAL5U0BT53BD0zRxxVy+jxDfsHLihCTaOME5Uk7fqud
bMrVENKJnAurH0Ugu7dA2KeDsh9nt2MJNGTRYwyYYZ8lV/DJl9sxIZmkVXPsNUlIY4zMmtFV7IgH
oef9CEKhpkvY70kKecNvGq+g46EF5BK6bVFlrxh43g+SDmxUQgzOn+pincaypTVJDq0SiWdfufUf
66XPke1JzWF1zae+4WEY5yTOTIOD5dkrW1kthGrPp0wLFrAD9uVrLSXdvW/bniPsFOq5FmEusZ5W
XuVAHlbrqxn+A7E+KFOzQz02wbhG0QGKF69HfaD0Jmq9fmGGdn4nMpdaHmhut0w2dPBC81yyX8hJ
xz6kMHn3CcXkLOXPtjg9El7wirOKgbqdoUUcUjqhTmAIa29F6wY0Z83lIlsBuAcj9AVcS8HZ1p5E
57rO+OjmTsetTBojTpJ+GrZZ95FnTde9dzksXH4C5dGYSOi+QZNk3WKpV3hD/mX99DVeoItvNBsm
V78yvTqKNyrHvdyp+dh7ptxWkVExI6bP9HpAEvWn0y6Bi6KcUtPedZ/bac+FdiINrWIoad2rHLkE
T9/XMQSyT89ULzIwBj/plBl+tHUgfcO2oro0VcXICtr+h8A31OPZLbYgzPajfOzR+h159p3hiQE6
2TZ3IF7KEzlXU0bN4dqI18qHqUG4A7YMmgmI5AnmnXarIuvZx5voFiQx+h10+iXg0L3l6AeG2Sdu
t0at4EhRpB51gq1oWAxSkOtGST23M7Dth2vf4aCV8lvfxRSYU4YRHmeC23vr72hUkZRlKbeKRxtN
nxlbDikeujkYHEgx1O++i+PgRlaJWEn+ViLGZnCzZ3UdoN9bI3EWt8rsXb6SlAet7xiFV6XRUW8R
tUwKkk1CqRyKlLJwsKGzhYLCP6AaYMuIeN2LVoCsTzJ5JhCR0R/iEo3gitC4B3cNvWzDvN4gGZJm
Rhk8a84b3AjxoNt1Vzl0EnbE5y75WeW6/6tZ5TZhpvyfjUmBxz8Wm1yRnok4UNYECz66RdHwiYXE
hnrm6Ln4rKEcWPe38jvePH8H3MX81nydF7s8sVbqCd/e/kxprWrX2h51wlezDrqbJni64PVBtqvF
s02BfTNcEZJJxziJtEgpYMG63zHNVlx7wx+r6K7uSDUtVLelmmHy0gr6KrPVw2lC8O8xjG00eimx
20HYMaABOap/TEQ0nMt67GI35gTxaCs3coDytnZ3Gp+0gIvrWsh/12ZJ0t0liglMfFzBFEUQFIaV
yIh302EjlVaBlO5q5IFWt4CVwmCfIxtIB1ffIW8obULKkk/UT3KkW3nzuHwJcvuE0VBw2aOXjv/o
tKTbM5TU4Jl4Hqs+jKDv7nS7KRF1+UbVx4NaWYGWDMmI0jLdxpOv2yxmKsZMndTuLiLyoVdf99CN
nuPk5doJaNqPA0fVEawMCvwsST59M95bwNVTPWJ8OgaKUpyqNdVHiKMycS0+3gxnhM7a6fg+uMmC
enfioE23208sF91P7wMGrWdo+qHBVZqBeInEFPKKPSGydrOxVB3+iCx/t91QIKNn944LjoUBnFaf
yOUYk78kM2ktTD0mh3PWMpG3A8VrXUksEdX/KkoHN1+jT8vCKx2OM2pMRsxlYlnwF+/O3kw3udmU
aJyR1niJIBliUVA1f2qUucUPX+y1sA3+tlEs/SnoFixx3qz8etLNaH3XF1wBFujakZRY20aGoRoE
6sDxiQEKQLNya9wITF4KXj8Of2gGn46Qh6RZsHCXfMe30M0YITQY/zZhv3+XT8GWKE6acD6CcgT8
hraXuY7Ki/5ffri+N3wIV+yNtr6vUjVSdLj68WXpZPME2vvQ61zjrPaSzybuDzM3Vcg4V/remY0K
tefakGJiX10Qopr8pGMM/po6WfBSiwJVdQYtW7RBFBdBKINgvQwqdgSMQqGkaz40LSDly5+uobv1
cG7idln3CSgdZQkUanILDvvX0oT7IHTYcsq9XWeSisbvC8z0/NKVkMSPxEvCF02Uop5y0CBdzxnm
tw7sSmAOx48reXxYw6h6hv2BRMwUiM77KVk3/eo3A9AK0doBTE/s3CDI/shFPYdDgIDVWDbkDYi7
6oED9i7UsTs3/wSjvZ0zlCCQUfH1dpFQdT00QjcR8yeSKf/Wo1C0OqYUH5pRUGzt3Vork0t3Xkc9
R3ZqDdkTxR9eu/ZWyqnNq4KVzYKrmjcdyqXbYO05ddSZSFw83hBUNJ27r4Dks7LGCXEo57E0E8IQ
tJBYs5uDh+2vlV1uasGaFB+UTfToaEy0dfNhu4xem99hLre/7N4jOiSg5IdS1bA5B2CSOiBWZzre
AzYLmzo89suUaLUg3Wohz76HF/1J1onCKoh2H7FZEDbwWFNHA5FwuSDKZyVym3PXDQeyp8JBSfe6
U5WX8e/CVZ0DAkmXxvq79j39qdzzpKNRwjp22vcuK638lzh1TDtgplLUVdzHLGl0ej6qMSyct36x
LjaeWcop2AtYuMEGXtXBJL4xiDBgu5b0nwmIAi4m/by/FuSd9mblNPKPgeTcGuWdNOyQRL8t5eX/
TaPgc0bv2KzdD+xscdnlZR4VZ2PRivmyHwdmk7w6Z94lyFXN7BRm/G3Ae/MNZqTG1nihaDqpwN4W
lgbnmgBCOd8mmQ8HLtyrD3fRbNiVaZi3fKj1YOi8FuTyv0qAzhlvu5m/5i53nmmwmFbJriJcpr1M
1UF+aqPorXzl56C/I3hnKhfWdPDCPz3u4Z/DFKMm2jQr0UwIO8Xni1gbnDjWBBCy4HlUZr+q3hWD
xKsgQHMCSwe5yJz/y2Xy0+LvQi6j0cyStv4xIbEk/f3npWFbvZQFiITJ6Afa9yt2xJj0YNi8uThc
+bC804VIJqvg9UYc95nsaO4oPxpPNN2JMWV435+LjvV3j1wClOCH1vA2tPekWmVenT+epGPQI3Xw
c3KjW5r5zfyW5UL6iS7fZbsQm1+DEp67UnBSaER6jTWMOb+rhbl/sxQnqGVOWMhsjk4wwM7RoSke
BKmNCTJoiOGVgni5sx3JawA3uwe55GOOfOxJToNh2OmVmBvFyABsOZVIwxUT1ru6YV2uFuivphRN
PptayR0ucwY8HXdLK29BpPYVHe0jt0X6IcUXW37bEqpv31463GHHiU4cgr/cHP1uML7tArXEuKi5
eEnQ2LSB9gZ+hrlbt+lxz+reoPAuO0DH/zc6GVnw+cUS+NEPqHD/gLEfZ1RJ29VBdCMTiK9fr4Ib
KPNXNjZhHcvcd5FiwE5YM4cP4tJMRntuIXTiUMVjnwsCno/98jtxgVHTjIw1slRKvtWf/EbYwZ3g
GOUGoBmholzSriPN+Bev5GoFlA9tZ650vQRcpHsRbpawx1Uw2nIhLfDoUPkXe19m0SBmszYWDiEy
VshzFNEx5z/MjBbLVg+V88Ak+kNZIvYERM8RFI8mlPQbZG31BDFyCE2+Hwi2dowDIwVmAZQfYAbb
96UExn/mhOFtRw4OViepvTEEmSALdkgsPanLKCHR1Z+HVEVHdnvP+9h21IlIg2qZKQDKaLdzqI0P
XmQTk8XfyqNzs86d8JXHAQBB6rKrmqra5nPcZuOs7kHUbgyxP1FgCROfrRRUgSXcRW9/YMH1MCxr
z5YSrBsAApz3g/BfAsHqugnjz/6AH6ftGiBVx5RLujkaMGgwnBfFaQZAVo2n7PIXQjiORWMA5Nff
B7ybaB1qRvG6cl1vsyIZ6V+Bq23/8PfloLyIyCFLgPDXtd9nRbrHziAfaQJHwbMZ8O057Y58XxyX
2zj1L/c5L2hQBeZs950ay9VDPvYFboomCKpJyvuE2Gmu2Te6dV0UBbFz+LXyvBpr4u4R5jhJ6x8B
kHtBDRw6vL1IrSScG4Iyj4azuiIxrPdpRCFcsbXjs6ySAwil1uRQ2GukgM/XNDbTzS39TuNng020
K2IUwuY5b8/c/MHZio/zzASvn2rSQJnAS5SiLFywqKtjSvCb+ZuYnn2LdQ/yhk/nBc8Gq16mN7wM
NM1E0lqoPAAnsCT3PNpxYP58S3498MiXpdx35M4Z2EP2920ZaVcI+SY4I++h9YFi79a6EJ1T6QVy
zWKW5Jo6YoeIEo2yPdwBSl8se51WLC2u7v9dX3wghiOqduOvN1G7ZzcwcWq7sCwyir2/oEnp7bDV
Y5L0TImEh7KOKIPP3B8zpCqGlhFJqUKIkBwAVc/0YY88Qw/SV9RJQnoDZvzU9JSZSCg8hxxCjo6+
Bsyjky78NaeMAaQNc24Vb0GX+sb3JaBqZ5urAsRLj5tc6C2BC9+MvDqwY89w7nDrbkJaSIQVRfdF
X+GrQaISkbJ/DuVNrg4S2VpJtEcBrxZ+4NfwwqbCENUGJ6+1fmTfRm3hkdMXw8D4JTi8WorxBDJN
4yTrhl/eoL+N2FgYdxO9WttaPZ6QY2dxGcXfB7qy/lZobFs0Wr5Z0jC8B6l5K4bAcoag1/jS1qCg
UNJ8gchLUSxc5DjMEFzwjXMD9NHaLkOnoz0AyqgQek2PhELZn6Qf6jt3R2TPpVFob6GS/AaSVmQE
/4VWRVh2U3oQWaWlXp0BON0AX5yKAU7tBREkPdjCyDZYqJDPEd+QcVGd2IPiX0E2edkaSRmi46ST
7Nd4YONQVKSUfvKDnMlMuEpx4zIteyj1SodiHN1t5Hn7M3C46u4M3sMEVt+u5SxR/czU/2GRmxkB
gnivH4X14tdNZRQwNjdtToe8ITumCLQsj0w1/DkGOcYM8/h/qtlaX2DojQfLg1mQWW1oQlkpmLEA
BaU1hl99peFqIkTY/0Nj9adOFjade2SMwqQsdC8PEOVs8jh3hiY/ct2+mxsSwiF07xp3rq9DEqWm
774TTz0cXjArjecrOIomQJditLgykWxoDsWHkFBpc5yySnk1UhtNC43hR1YquZt7N3txB7Xldxnx
TwN89rJRQJZDqhQ5bwLEOPAlYJdLCKlFOft9gc52+UqPLULgOPK3zos2KJgkxGA19Yc7fx26b8jb
JNO83vPTdy7RkEtaR3PCiw//hdFLqL5qxcobWelwCTHLU4Dlx7/ou4V0f2AhT6sHNcbJSSaIat7O
oO5IPfxeAsDxICg48QHu70KmkuKKsEEV3TzaHTZYaX/6BSlk6aKAuAFcK1OhFiQnYSXde4UIhMHw
yyaBO67IcL4ed47RQPkVzan2TxEkxLeXcf4wSm1Nsah7bpqerpwpoUslbdj+2kTo74hrP+UNjFZI
AqAV8OJ88NrTXjQJCL/7NJ5I8Reb2jgZxjRjLTOboMj83OClHTCeVkW40Qa1XCeb/YQ+A9MeBaxU
4zrHE4KN0/5cKAA9x3SarZxta6DEkY90TdqjCN2R7lV+l5K5F8iR/NVTxbBZQIE/+8n9MilQfN7+
fGCepBNieyzMvYGSj3OhAoGpkF7/wMdcKgPmwmkL+8rBKKYcqGQIzxY0GdxiVwr4e1WXnQzvOGVE
JuHCBXfr9/IXR5twW+47+py21AqU8D4kg6C+P8ArsDm4zqh2KuXJ9bjqBXNaPOrX1JtyCS/Scq9o
YHHsESkUxmeUJELSqcMyszT/naAK2bursTv6mYQM+HWaep4fXAk18XxekqNEM3FdT4yH8eHtQa/O
GByQf3s3iHnKvXFsUvQwma2FFEU1wm5gid+cE64Bpe5+ZmjxZ3XgfygBzNAb9z1M8xj2OZuQABxf
iqO8IhsPDZ3cOa1I/JwXIYBp2gU2iDyKJFtu3zPYvjQeM1v6eDV3JVFh8TW+D6ZNfDmNcE4qvmAN
Rzo/Dv+cD8v0OSxDsYDv3WblTUIezzl1saqNUn6XqwhEZLKdKW9j8M84TDIi9XbByi300L1+KU9x
RjGqNbW/BEeqxa/0hKwoHSBQ4hDDN4k7xV1eGSszgtJzMwMYM7Ep6Arr3OJzMeDJ6autD4DeEmEd
Ngox0llpFaZy8g555eirDL8GFZB2JIgOlbTBLCKHByx2w2LR2Fp4oDlySyJ6Pv//F4ZF1ztS2RGc
D75bITpPRlfkAKIX6WT97mP3zsLHLUzlNnxqRKBdCzH5pGTjF+oIEz2plFkywaCpl6mi61c5Ry0n
LbwGgEEmdidEIivKl3f8E6XFilD82KTzLFRjoABKiEth5bPHJrlQjYQym88lKRElQmqxuCYIYKKc
R4tD/tCKT+rT0ZTQ6r3raISGCcj6KPBMsNntFq408Ou78T02vqwnXpmzOkBIcq2bBlAwCHrI429V
zCkc6C4k0khw9kOBU9yOpGd0oIvJw9HonkUzBm8NCZxBpJANJp4gG6pfQnOJnMSIReIDph8tIr7R
26OgN466pQg0FL4OX/BU7jRzpbgDZS1RbEEp4QFxmfbmvDz1JI2YnGY7Y7TwWK30Z0sMVVWynvDg
oRYxjCMf31dQiksvWByLwDqVcvsnv/LiqgcOot2jRIkdb01Pn5dIiK5DbecJsJyyULvZdbWnFGWE
H31UCQQ5qW8CXoIpYcbkBNRla3guAoraDxE4ZwNYqFPgeqtpoveUqbyhIsdK97gICHDnlsMgccA5
//QbbtmstePHISdVTkHy1mXllJlnM2di+o9ZDkqGCq5Pwj0eJA45z+NPqt8KeNQ2QwFZIXCHIMmN
eUlo5aT/DJ+D+2S9YXQ+yxmYdSpmaJJtzXQzSyw9Kt95TBeqSANfkATPF3eyhlipDdhCoYtVu7B8
g+aS5M+FiZgnUaz3L3ICzLOoqxbcZ6W3dcX3R+oQG49wMoDRkZvSK2Qo8n//f7bkC9aIlU/hPZup
F9lMKJV5mgTSV7CDUxihY31NiQT0+BRXrQJgmHG0lapFNw9vZRm7H07KLQW+KtNFiXpV7kmZI6ln
zBUmvyAOsJGdDtLrNx4YNUV/3uTtBAer6Q5xWqj2z9fdgqRUwgtTJOtnwExCO/MCRuVzVuOewApj
p3Ymuq/4Z6V1CIZ0pK5aTcW+ndCtpFKF67lMsBbWeXoUNSz/shUA5MXySoYNIMKZzkdIBWwB9kyZ
43UoaK2OmjM4An5yHL2xIF8Mf0dPA3feVm9bgO9okOUiptF9EpXQfg1PhqmFWNHEgrZnLl0d8Vu6
jsot9uI4qP+WAH6HYQySzmdosnKFr9Lptyjniere3EdJi/1jbvY422RxXMwc/Q8rIYvLqOYYB4Iy
NbbmXZi1ENE+YUl8d8hxvnmCeatwr3f3K71I4xlT5oJSlCQYOHftdG8hn/TLtCviFp8sfNEuDLWr
TpJD8Cxw/pIw5kymQ4VZBhPudo5gAcDRfsGRy/cZnKIulIcrYWHKT8SqjIsGm8OXAg8iT+2s7vim
QNxCjVRoQZY++gyI9fNb36u94lrtRAvjnmUTbzPf3GFLfSdQOikw97cdYMcd3B7FaBqwiVseiVqI
MSCGyRSBBrhYufg9AUrrWWqBkPCDk7NkvvP5kz1GayOngpGdZOnqyQ90bmogFDTxZqTsjCCISvRc
RKB0UubYHG0CD6PVz072Pi/EdzyDYhX86Z+k0NW+5elX661QebCTD7yKugv70vJYRfvepXJTrulh
ciGs9jkqA0O6oz/3yXSGto+6OIFxM97+s/9GCru8SjoZ7WrdqQiaAvXWUex9N+yvWFvtTWP7W+8N
d3B3xxMpTU14wyu8rBQDLYP4xjsirK1yuQNu5ZL8zDxpbCzOI+z5etJGcgGRvooSC6GCu9J6JR7n
DgsHLyeJIMSP5cdoT9eOZpc+b4J2SD/YMHN5MzANLWmEOOXbfGsqmZjkXpxxh6rJBNEbDWxv7vJV
GRoskCXEZKltC3h/Lm6Ey80Hu6wd6nNnvv4YrMcmyh1tQK3gfmDzwRwH7ZYHvPOdnf2ZzIL6h8lb
vPxiJRyHNTDOrEeC9k2xEFx1O4IQE6uPbkUtZ3Yl9EBgfla5JGudLq5Z/2PSNfcIUIPPv43cFxqR
hRry9+JF8TJi/lngMl9bDCXDWexCX7r4M+sXT2/H3n9m6ZnARJBRD4lOceFFI8JZvLVqiyxeTycH
0DDntXBJM52emKHrkcfq/uZS6SpagZ5t973L1MjjUswZG3j3Z24l16viAiSKu1z3dN0xGryEBdt6
2ixIbF7Hq0tl3M7myAwCRDFqgyzc+oIH4NuzAaaywgLu4S+G7wfsyEtA9nMLVXYnuQswvLAfpiMR
Z6Mq/067UBkkR3JKHNX5Lih8m4MDUO3aQfDgau279nflHDapGTP2DrlyilnFNs2fCFIs5w5dN0KY
8zfbd1gl0p7GOyjXVaklWElL1Ycnul18AJCc3m31R4LIhR8AukhaS6oqZYLlqBTkjUtG24SZJ6In
1ZJoDn9GFalHyZBTFUnfx4kLFCzH9osCZjmFLBE2Xs83P1kR3ZSVlkw7C8xU/8G9yZVl/a1rNZKA
7A3pOCZAQVNjHVx86mPN6LcISNaxAbuDUFjANKK3vI5LnEivmwVVLkm66PTM+Su0ggddmPZxfEp7
qaDvWIHsvyC0Rd9vxjkYYv7r3G/SXpT+NnHsR7WkprIsTP+z+Pp5v8ICXlEKBO1KUwiyDGTccrwb
eJKOiNT12f3epui+uRUa1ZZlzGUJLgspuk9f0AWdkNrVr97kOO162kng8NwUxQPGRtbW3OrOFyHZ
zWG8trNgjt/nhn/irhHfr1CC+NqPjTsOFyLwaz5S9Xzcc1oHppp5V12WGx0DEYT/LUY/ykdYpIx9
w+uKd5HwYn6I1m59dPhuPXfbo479SN9nr5mORqCK28U0Dqm2kMw4dE/oMREtvjg955wG037G55fg
fpfLvlSJ8RLTLg6BKKG/Oj/rWqSwYTaU6b2ltLJOikiXznY99aLZQ8AgILvwUy+y5S7vwiC9Q/ui
gYF7H0AMM6gUlMqze1aTBzKUOfa1osu5Tbtm1rHFo79YZpjZGjpBNZ+miEwfNw229S5qoidt5mF5
ZkSGmVq7jhodCLrf3KItczWHCDPb9nLngLgEx3QvjxMDDXxq7UuiqPLf3h3YfUqOlLBpx+mPyf7Q
fufZHra7pT75rM6jhM4GlGVIObDRU4pvxjQnz2R1wkESAiD/UdGAau4+4Kh4Vm4IslNKnGgM75vT
LcGiE72LHqrxO1S4QtC8SYq7/F9DJ/IF+iIF+SBBn1P59JJSv1R4twL+1/ZdSO9ZcKYhRwtAOly+
ZQU8bnS8dsMg77/vNvIK1zisINet6yHRM/+9S+zpdJxZSlJQz30ECDvhThC5XDge2ppsCOskUmjN
4pnRUCyK1tzn2R12Q6LjFo78hKaFqU3bLlsF+hA4eDSKoqq+kSA6z0+WCwH35srUdtGS6Xka79xa
P0nR9A706uXiXKClqt33V/o5EJcTp0gDrIQhqlAI11OnUk3g4T9ee4o/X8gUO7AWNSKOh2zfLYNN
ajJNqeeYcNlxWDnFsPD5COwEi+RXOcbdNyAX3EiNM7tYWE8WtpYT3sVLbPxWjYvCsRFxvFn1JHh6
KtoEBHSGAcV4dnhYdhbdsviZ2ZTtA50WCC/mmxLyYHMghM0UUGHmZxGPBq507fbGC4tQ2+nSZWab
r9Da6bxHKxOxkCFivKwl2Sz1Jy6GFIjTBq+C8x9viYMdAw7xIx/ySCvQnYKTU4gxAJlXGIp1WZW+
8f16vtqjB8TUPa1bXQT52Zydkp/N7sGlFjquqmAVSF5tExp5mahUA27/JXQMHqMqVv67BW7P5gEp
+eBXHqZxOEecuQFb/iqJdGjur1NHQGLqzMT/RIBaJ0XbNIJ1yGNCHiDBnlfbAd//zTsSKgy0PzJi
6nRa/fWWvcsg7NpFa4KmFcvvSDWg2c1VYEeqTVceimnRHXLKpekCpNn49XThYMws1oCHDqliFZh7
N5HTt7tYVHi9u/4+n01jRAV0z5ivUjYQ0scfq5lrC0Xk/eqz2qxVIpjzYqUzpD73pAvA6d+HEXdY
5ISOzyUMd9AA0SxgnO4+1Col+tMxCMfNbs/yLi360hujfox/3ASrhF4sez2EBBxh5qE3DMp+nqKq
hiPltiEl1d0YFOiKVgsH4BElfFS6+dN8IRsP/hm9JWX0BSAxhd6A13Ljb7CdX7MB9ssnY4MURNbt
oTxfuG7mfWMssV2r7N7Xv4lnxX8Yl/sJydXhNN7WUbHklQhQiAEkPzwdgfnq71M0gPllSscOr41N
aAfxVm8VKWrehNdDKnvcTRbZkEWGLy5HcBBI7DRkDJyoHlx0nOa4KPlpicHuHHbxzYa/bt3CtdpF
fIOWOESxkrtvPx7utc3P0L3bT10lIH0PzZiXUs1IxPK9Rfgmxti1gFStBUCKy61udv861/3e8pYh
hknL3KHviK/PMCZGVXkaaaG90En2J4U3cS8RbhrZl1TgafKv/j5zPNiBxoaoyDLKoKMC8QEdL13A
6HTfvgCZqBIUL9JskAtQhesmXMi/86b+fe2TnoUKyNTLX6ZwLln9Ec/xtvqaEe+JMZ3xg0S7HkxI
LqQA7/D1PzsqNPStKDs/fwu7y1TEiPJDi1ofXZrHH68eMpbM2GeGzfqUUKA+Znd0rihT2EgfXtV8
HzuzcKzPPYZABtDTzaEYVPzWZDilqnVUKs10rwCZeJUJ0kTU1z+sJB6dinx9FY6C2BXRUOX2Wmdd
skFqvWLjCQwR07F11VEEzqx4VqIO/ipmJiC6ZOEcT5Mk1nxB61g+M25jF/yzx9TuNqNz0xP/f8ch
7BhcDBnkLPypJ/duladl910jGZfJTUJpw7EwkaRucCGp+m+g2l7S2QmAqIaD8eP78r43bEyiv9J+
cxLrRnHkOeQvX+zEyxNieKA82wgAMHwGo43Fqlxd2oqu7K/37ReHgBI2fQ9UvvIojXnRSjWKH9mp
e27TVN13BLmG4C1yjl9FRZnIQBsCA8bk77+4wCtElq5yQBcIB2ZPiTlq+i3u9dLULUUtA9mXQXv5
K9MtKoc7FAbjfXF/YxCpcoTQv++mCSdXW5/a9vN3D96D5waglo6CPapi2eIIpwUd0/BDM3k3XES+
ilVQUURchMhmavVlQ3ftNxDzXghIYYFcbLMgWr+jc9wF7Z4s5BYXxM01lcgk9mVcNeJM1dZQlZVn
MkXaRzAGkgf9pafajWBIyOpre6y10sa0sgVBqzibk0N68c7zb918j8jZWUZn/WAspp0T5kWyiAIt
uIGXdlDDwOzhNN250F4ReCmllKCvnFDdoGUhKEiw7pM9IB9mS3XxNsqxO+C/zPbEeWHvD+jMEYHl
T1p60ATH4IOQypqBYRByJcDLCVTzc+xKfHhahxvrVz2L3P2uJdUItSr/VgvBXyjKhahE57MdpYKN
pfV9ozvnWuKyk4jXZ30GLCB9GPQQ+cmo7mJR5Cn709JAxoXAb3IdjsfnPF1BfBxgNzFGHQY5UvXr
jdVYphETN+r0I3+6H5cViImhwMbjKWTu2WV6z8jLjurpm+Fjl77Op9uhs8czmav+BMoBf8OEqRPZ
/QjjvstsuAYZhHLgXiazRxLLgxzllpKSy+zRaTNHVazxqlnXjJu7WsZ4pJWlr9nTsQzvGSoQnwSi
//H/hBvSU2rrhwEMHWWBnl388rtf4sLwAdnFKTCGhF60Pmunt5EOABMTJj5NNiyzINbI57Y+00f4
GnkDxNQcs6LwUtbXivPRN/h4dw/H0SG4VJEeTvCi82OMJg2IH7ecco2bLsd55DS/Svy6TnoqOsj/
ayMZe7t8HUlu1TNOK5Yzx2WXAoWWrJvz7o+4h4J1I+wQgN8prWCmoSmxjjgXlFskBQVcVc/kT5HT
3Lzsxbz8SCtClWT0x61SM80ycg2SH3jCUB3uCme/Sbsk9ulQd127EEncksMyD2p7x9yd0qyYjB7z
6x24p214RBQxuHyjVKtnt/r1V6/Yg1OnPNMMDbh8jQfuxW6weVbYfsV3IjDLHH0Xf3tSFGVIPj5F
JGSK/c5NKmG6lHU6DZqWVgIeoZS1u/yRuuZPsm07WARJrYZe0jiqInuqUP4/Zxihd74Avrqd8q7Y
XQjft1jZtFQfRQzpim8pkJcC80zULh36jgrLAADkM3C/I908zZ7GrgDIh0x5vVxWL/U2xn12BIUy
fX3IF2qlij98YX9CyA1TkSjfZ4XkJss8LYjJMGWbp3S4yEqTUGep2KJ6XxKXTzXebRTj6qwhKi/y
WakljEZIAX3kuIuMIQK2qN03aUAilC1U21epIKN++L9MjNH06+kXHW92JqVnTPx72ySCcoS64+pB
YsQHpWGjVgnd84cywbo8Op8JQF2+Z3nvGH2QSv9iOSs7Vk3/H0ectyDEc6W0qFD41jEf9kX0U5Zh
lM6N3umJ+HrprDDdtorjkrV03VtpPq54FxGCo1wi6aJAG0HmeBILWHEnBwzvG+bb6kJIM3SBEAPJ
CM0qSjk9jj7K0L41JNWGXd712D8d/xEU8+Zul1TumW1u3pdq3GxrufnMwTHKlnYoTu73GItUjOlO
D5IlAlNSvNHl3cW+qRbfiUlj2vR7/wcZ+OQxNs8BH+lF3AL1YeaTEf/KcCeAth55c6yNIq/5FzMe
WwN+zsuGRqLy4Ak92XePGSLkcqbPi5CJQrlLQOECtcWqzpMtsUQ3uHWi99ZQr1CIIS4JMaAz0GSF
7WfFB5kCpj9IXbvroRnI/q9LSbcxx5WSVGznbQbxS5N6EW4upBygDig2dUkcKpq0wVrrmHd5WL1H
87EdKW5A/DS42tBj7/iAfXq24lx4LFatqsFEPsuC+hQmHi66q3gLqY7+kRfv0sfQwdz5Gg25z7zA
EHcy1GTIXVqYNc6R6CwH3KjcgLPQ4JYZxd/hoYNuZUICGRHZ7YNlBj8qiyZz607N4ieRiS7F4dDy
j1gushEdn3RtGhZ9LsrNd/xY6p3oqaBa7Ht3K18N0ySeQ0cKCgLlRrI3T+CMEftySeq4q79qw79G
S5uvKyLUNm6fhsREku9Ma4TCpwHsHoXR0f/rYXgKanWutxGLhEhbb79PRspndB1MoVdB46Y102xr
6yz7mqUnUAq3NZLXZmBr5OMD27RECfqngtf3YuDWHuYXRgGPIItceYCNlyX3iC+NQ4XiDsx8GWY3
JENnQlJPSLTDYXMnZziSpV+Az2aNV/Iys4gaIMVy9yffpo+ibGb/AgiG5nplWYjLSEqEi4b/iVb1
E1NkJ1YWgKGp7hXxB4jl49lx8wDdz28mClopPvaPD82JUysyXJS07vYvf0il2soPeOj17FnBlKrq
1/HiQ7dDS43PAzehkAlCjL92cH2BlIpTj5ooG0oYA3xa0nI3+AYNBZg/U6FIVcDXXW6zQDffMS6K
t8QNpV2fSJ0nIax1h+6NTNWl07XGxTS4vi7V6Wv3h0lk6FJcANJw/hvQ5d9YQK6RHxw3gBkhD0YJ
lQEu+kxNMpKJMBhHuvumWiz9k+IGhB9SvG6rWs+GiDF1UslOtoIy/fsQrroXPKmw67eCy4bbjcXO
ApxpZljw6j+U5a3mwdmKFXt1a64ClvqOkb4ieMytDO4wwuMLsSvxL6F1qe2e0D6CMac6WD+aguYB
UD7yhCbXLpSsBvBzEtcE4IBv2N9TxDw7X6ExkK7YD0qoep5wXd6Sb8X2PwqmPH3eSyDI4w/TFD1W
E/ur2ZLGo2ZaKguGE8O3TfzLlN9Yoe/HOUAfck7L31/dOiBPi734rnWmR7E3NTdIBNHv58vFYuJC
65KbA4cB35tpuPGi7HVCquN8j/Qqr8SYPt/A9jozTy/cWwJvyh24qoANZ3//4vAmf18tSYOGyuld
Y/DfqpOBViYLDLVQsO1YSEGIyCWd0PFCP/Nz6FhTYRSaOvrc805TllSrL9xZkJm8v0jtJbhDGUWj
OgG5tZzUPAPO+I3KV7a8mNY8h23h7huyRh5g6CI5Ql+P3QnokNk++ZLi8uOQA8xFWfxMeSbMKsOA
1lejfdFvLDXw5+8grIABcL4HOxq3YhOHyfS+S89HyjWhAQ9SMjMOaxrZ8n8f9OARhEtPt/RUAwjL
LXoRUGwVeY04vKq7Qn/NSkDSSHZQzM8oFtvlK21b5cHK7bOVvtfMS7w+vUinvmCqJES9mHyJA+l/
cNqi0GFDTbfaJmPf0jOsT87rNR9wMIxC6I0nulKphUrVewFG0UEjS3ZN5WdGdOvsnqWYWlkJeMMc
VQoaIoY/plKvq6CXA7RNpzn1DYws4ZbEaNLRvHjx/OHKJRluuOcEsUvl4xHEOQTwDNtdz6dKWDFp
I+for+QNo1ibKmlVmGWc40R5pT+bxeWi1Y3ph5XOGvmdrzgsX6Wz3wLvDqo0mrc2Q7bWtqZYs7Dq
Rh4jvL5CKMadHjDGA4r6Dl3Q2Rj5CMkGtg/QaO7zsRjw7FRJNk88MFouBZGzEeYny7HSfJ2pszXb
oXELMd2HJqwI5ylJY5fk7zgnejPE3o/VTJIvksuM32rTCGouzo2MVGXS8jpUaI4t+84BcsH9f2O0
wNUxDVLY/jhIbBv45GpGGucAxXQP6d1JYKBfBk1UR4ZbkmA1MzD4pPxWcx9Mo50AcaJJsrgw2o8A
+tHWRnnBGHArPX1UsGs3yH7xK5LjnmP3waqWia8Mcq4UtMaptAbjyCung2YwDn5+EWWQr9fuDt86
dse1jOKG0uISAVssqQKp1iwr/Js06xQlj29jeKnN7eMQNDBMHCq5LZpoMCRazD+jATRAOrlnKc00
sclPhhMxIFfbgafCXKOFIv0gNmkXzYx9EMJyZrd9X7N3ZT8CZSNK7DXbjAlHgaBzE8iZdlC7VD2V
0MgpHIk2umGyrQe1e18P3EB8pwGXVYHdUVmZgqMHjh2tRQYHmhCKN2gWcUkeSs/5339IvXtDCBq+
ZjDKN5+XCazHuhCjBE0Z6uoBv8Qib4QhiiizLMYCLMN+FvGmVWauuyAMOxG7btmlc54cPpBPLGaT
ERgCra7GsIyCgLM/iWwTdeic8gwjpaOLJecK0krnGlzYk5Smxb2k2vsBYkFoWUaejkboT1EiL1Y8
f7q7vfbsb+/B85cp74XIOfX7ateNsuBmPtSRaxqKlT5P5V2cpul9LMa8Xz4bYNJia0KHKxEvj9rx
S/WM7k47Te+e0FdJMdp/K/rTP/WvxKkcQER1dbmvxsdigL/ngLlQA9y5jFrDYN3iWtIJyqUi/CsM
STXF/wxwbBcYU/6v6nJQ7gLmwuy6lo01mwYR8AWnjrZWNzKH8bqpQKINp9cfOEPiaYK6NtvyXAYe
QnmsW8gnM1X8aWaBs3L3T/TkbBrSiyQAw08EQKo1wb1WANuwCuCn1iLD2JZP/HSOHtzeugJ8QzvD
71ycfkIUnRlXeLM5LEYYQPqUdSK0jmkFo4/ORu75XJNalHS91RO/emJsIZUGSZK3fkOft98ZiZyt
fg4EAydcZoD29QIlSW3HkE0mheEC47nS8yn9lNTy7xfhG0OPRiz58rtoQ186NguWJwcZWNSQ/G4z
ddryT+WsUc3nMZztZ4JZ7VsAkuMHQMTuTpLLKeSX0+B3hPcaUMEyeAbdeX91uCzM0AhLLcfcFQph
0Og1g1iw+flsYCvFDvy7I6EJniwRIP0raAL9Y4+S3TaOi+/jM7EolmtAD9Y8wD6HEiUYsVmieWow
8ezjV6DAsWCS7HwOs7XyaiYzUHJ5Bb2Vrzeymu4V8iw2nEz3QjNXCljnmKM5l9hImg2WZcyGC3JP
zXSrjgAxC7wrSVm18xT309aZEnG4SC0+oMdmsrrFKsUaJeK8dC1oCnnBh+PgCtU7mFSDC1YiBXiu
9YTln9g8w63KqbLqfdiRZTsW7SJquDKIhB0KDU/A3TjzTpCFfHS8N8f2L0PywZC2f7C9ps+uQuwL
yRLxXUtoivEZsIucR/Lr3SMn1uicakkxqxy7lgJnwOdJz9dSvb2fNV1RvC4HL8edQBw2S8SbRGaM
Vh1/Lv3E4hxFvC9+2soUPHA0TKHeQ2esvOn3os1osz9zw8rYgKHoTTvkFtnnpi+9PCtWITt0JM8M
vIZJTVQymBK4oniajM8mJaD/7WkkcaxtGH/JpmdDO7Fp/h93wd1UMPiBnru7t2yS0XKswdRAhrBF
2Mj/t7QydY7qzh7lcCs4qr/4kZYvEtHZiWcn6b80uRovfKsdcmSORio4sxW6qfvOGK+nkJq4UEVt
fofnn4fBsaQiDu7+xRUaiTGm1Azl/QF95BPMDT4GAuJTUnNZuTIwUKISUWYlJgy+Wnlt59IFtsKN
ixNc5LRJw8XT8h37khkAiHxw7NAmG9kdpFrw+thcgLEImHB7Gr1OdZNCqoaXRaTGH4P53nXQCJqH
R5JHCmyV4dtbuN8uSdMcnIzgyVqsIlvq0LkMcKJhk442FYJd2ZvFbcIewFxTibIFgvGHabiwZ2jq
t3OCIEqjcumVh1ByRNpHsE90oFRZUbr11HhDlPw4TfuNhVvwK3sahj8gWn4939ZX8Oxqm/UoblIv
G7zSxUmvtd3UEqfTenvRM2oBeEkdgNuqfk4hwxRy896uRguXDVlJGgIqhq0X7FuVKEAWQSozR9OJ
Mf9hsxMyMlPRigxATL7KvTWkTAz6lkohTut/KRVHCHSSjaGFVequi5s9KRJOLlSY2KCofDR1fsf5
loZ9eYgOqygqt2qrhuFDuvRd+HSgOHI2AMKoDwrB1ZgKEylIqRsSYlOod9cQNqbRsisEStzlnJ7U
YUZyq0rFJEIy7hqdy1434axp4tQ/SWIfM/ZKchy3IUv73F2yKRzsmwYuDlJj1xfwtp4vuHoII4Qu
GZe+bntqsj0ME60CDltnAo/qFabl9x6JczeSempj9wlS0vS5rH6rXZ6wBf6Mrbo9WQSF10uGxqqA
J15y/sx8fcAii9zZHubzn3EhpGggy+TmyLrguRGYhq6LGRQfh1W8Gt1JcaH8rIoAEdPtOXNrDOHD
6BRF89QpLmxHJJDoRV0g555aMA9cdgNxdjiFYd0pE3S1xZJrAXc1nc5SrF7kyfOrf+nFFmRVolH8
c6p6Aj8bpS7yMH0eWGGvU45qqurws0bWbFDET+pUtwlRD1aJyei8IojyGI/09yNa3l52wKF/ILFK
ONsvJSgLE9gGoFIJsd8BKlTXsk8S2ASHUtQzx5jFL9uUTBInuvoGZ6Ov0fKiqrPV56wcnpic3Y9e
m3aTBZwsqrQxGM0OoGnTws5BseBoWKSL7F5y5xM2T0Ld/GjzFiuDv+HLAw3W4RO9vQ+yfwXlSgz3
0qkXF57tEZmIMhN0UhWjBN3CLbBxHNB5TiKEYrU6maVg44SfUslk1o8lkJGIWcnEZ+zt1MUZ66vU
jpbMDXTppr4qc4VdrOIFXLkxmwjdOelL49GnJn4fHMhXOK2adfRdXYa+LvoreFivt7XIOOGhz2iJ
v+B2qQD/lCYIMlFNVWWhUdplzZuu0oJo0X4BtQeqrNAEhaqR1SuGH+Rr00GHsvfzSiHBbTfMpBVP
BZsma0D4Vi4nsJpRUWmf4FldM9wlLn7HxYUYOYCcEy6F94vNC1Ar76Daqze6BatqsL/MdM8hvEtu
Q4SoGJ4Uy1YjXFSy5eyosx4eLHXSww520t1fAZ0Dg4HtI7PS/rKiqay0E9CN6gXcdxoaLfzNZzol
gJTYWP5JwCf5ZsPoIJxVfcNGW/w9jIPnCBuD7MTtw+uBVgYcTe/EA1zMtgwT8yDWDxoMeImdY2bs
R7jxeLSvrauMdvqpYAz4KnJYklD1r3qOgIg2M3YD83b2uBTY+KDlVxHjoVYGDzC9AuCWXA+z9Gwo
D76vRs62r+FArXurVOIIncEbSV2ArDa915w9uoYg0aBc7wkQK1SkaFM0KBrdEGx5NC8s3lW2v+tm
2rBCxgxFcO4q6EKWewmxay/voSdhhUZYwvbaw8r5g+uspdER+bxDREiCm9ey0A/uFB4XrjgbeEAl
8NbeO/U2APdQlxsCpaJ28Ojo5QFn5stmP7u/27WoHWx6vl/5sZfiqokm4n5yU8oUls81T67eBt+F
qlDalSKAqXM3C2c9Ln8/xpIE7zBGJ1KnhTJ/ZmGcpCH53V7qNNvYoPcsi3e+vyscmP71JsX9BYfg
0IL3QLrx+6/OVK4vaKwLfgcSO8439jxaEZ5b7Mn7lY3U5SuzTizZaNFlWBS3INPY5XS9kx98/N7D
LhwNZuFW4IwJGAsuc3Fwt1M86NO6UG7i05W5kNopEFyn5eFmn8iy5t2+MNycyiCa6EjvHrpj6DOz
Mc8RZ733TQdZ4QFYg0lSbbDmxqGEkVusViRC6kPfKKdpMlNOsKpBKDyR9AxXnfEcTIGPt1NAFNt+
ahzfLGhM7E+Y4CPEv1hl5PPKbKKEyrGHLzyyYAgvNoZ3mo479xSZDC3mqBBl1MBqtYjkEcsDXc4t
u6h445FSQAvggNTrH4dQb2yAeFyGJQ0r32N/v4lhx9M4tubFYEhnsJqXF1Jwm/IPolTWDDfsdEAs
VamrnHIhjea4geVQmOhS2qGbQcfE58zK+GR99a+YbLaJInHHpGFaSbV7GiBx2Tq5kTQ737TJMcjW
pkisTVnjEezxjTTR3HwUYHSvQhDZRVukOVDmo8i2maI2vD3el0FJpgFu/DZpB6vh6aeqc4MpeX4t
qsP8SD0dPTLb2uX5nkX6XU7MgDnh2W65lA7a6JAyyzBrJT5OuqAavAbTCuK2lO8P3vMjAz9jBidT
dU8wM3BZfbKLV5FRm5lFr4yORaRIFJ3csSo88xdD832o0CZoG2gF2vCIgh+Uio4ytS4F8nu45C+Z
g9xtAFHejfGRR7OlNJkTk3qSF6p3Si+Z4p+mw/9qLbUYhYXaJLnMoS8a3YviQ2+r0G1Wj+KL7EbV
PECcEleIX12regVme7maCJoCzZvmnNllsO3VtAYfXBxCUNri6wzA/3SAo3IyYQuCKwSL3YHrJnJy
ZmyL9hRAHYPfDc8hUqXQsDH4EIopArQOf5MkpgGjtR3M0fueKrRb+wtx35JIGKUFcTONo2k0+04D
BHen+XDJVQ5If5ZD5idiOlCqUinxoQ0xqjChyYhYHU4ucst6SR9ZShUQ9iSQLa0NcxFcTkhzReDo
5lIqfGKW0VdxrcRO8nzL1wDOWQnVvUo/FALlE2mSQ5woM7G+CxrwVsqWMagzsAw4wRjQ+XVvVbkr
YeTFAh7EzKm3L1z3kny6OQZsCGm3MoEE8OibWPMouqf2W+E5BiiRshmt1XUlBfqysYRnA1g4uMOj
M08IWbEFHzmYQ5CGA9rSpfAZ7FVvQiFbPr9dG3geU0KLY6bf7VD2wot26+Vd4/D2jbLHksScCVdM
krH/sPOJ3SNQVd/HkvpkkjQFo9NO2lmMDq/o81iks3XeEdi5CRUVzfXCveaQshQtLaXnlD2RAjyf
3xfV+NWhwHCy9S5vDPtgm8LBkzrbh0iYNzMA4zMWiXU/u6fNsA/YUmVcsgzJxuk/RCidJPNGf4UN
oiPt14HVAN0WM4/NUSvwwnbXe0+Nehu0UcQxOEMZpHq1+R8YIDUXbTXjxdOrlt4hKvwW6cBu5V25
SdQicfegBfiaAX4lkMw28LyG3Y5dBNqXHDAtLrVMR0gvvFrFc6CLC8Z5YvgLg5oSiuAgckKFHD0R
46vnGwnEAOi/DpqBVoepOvuLFHfwoQeFTdegWBJEj6CEbJO/KxjeXalyNqZ73Z2cSGmAwVhqqpQ6
1yrSi5duA7APpWhp5oPitdCYL63wrlDMXzPIZdeKykD9VB0zl1+zyPYZBSX2SLjTDfQOXBVPa5iY
3mQ0Vw6881GbF2jQqeYU7p4yslQdnhJtg+n5ZS2j05tLNM8XpE8w1Nm80b9phJSFuA7xIToTfK+H
Kq7Gn68C3MGOfDJjRdB4bQgzlwZF51T+iF3IKQ/xtNUXloKmfz+7ufDMXAbbvl1YEwBbW/vWiD48
c5aoqLwS6yGJoOzeVqMExg6kOOUdjfsZL02BWhhbkZPr6sUWF5ORzxM4L13tRsKmrpULvK77sISd
2fRrtILJO9MCXOojL6wTsfJ5Q7W+JVLkDiBDFAlYM3SiwDdRUcZjV1HDC9nbqzUxN0MukTaEpLlf
SRaEqLOEfQM4zApO6kzwyJ7zwF52aviDo04JbdHwPUwDpkVBjMAJRRs4dvFV10xvy5K1enZOOHzA
5dMDbGQSi9tsu6UA0SxC8jsqrfeiw5TYgjO5nI5vrHn+tAEU8qSuBJPIGedIF7kLlLaiOR4jyqJN
eNnAtoG7KgVKi0akHnd+k2hjK/xeTh+DGhaMamJa8nTl+SKWrnFTU2T0/RF9aChJ4jD8Oglw/KiM
UUGNX/uH4fFGgXo+purBNCGiuc/BPfZQqu+rWoY5TToCmsmZREm/vWd2xcdyvasnUa3mMLt1Gngz
A9aVbQWNW+cl+djBRhEFDB21WxcqEFgHFpr0LHLlrjUYbTntGH9o6E3VsUbCuaF2FtavBxWua0Cb
W+5BfFLuXCI8CSunLeGky2VhqKDrBc/rchbWMX3EHbbGYUDibxGtMHEJ60Bgkmg/kBBcJbALxTgA
3AFg4nNPaodAE03LQxfEdPUATqgnRioMYPch7j0y77OlGKWBzOB0nIiPlHlTqPhr3mZi76oA6TcJ
UAYCh4Ae7uvIX/R+m4wTHaWE1OERB4NsIF6TACstolhzuO0YfEgBA1ZK9o1nCkDii2Eu20Bn1Xyj
c0XwIfkYY5Lp0S6Zvsxn1BCxhjmAX0AmENpoTvmvhWRc7lDM2qvP/op+cyKukPQzztGO7Nor2AhQ
c/XeOcyn9CdwGDezwsblZ6aAGEyvV1l+YXa9swTMXfj2Fk2AekgH5VLF3obwE/0wzzwQLhyKAZWZ
RtrAn1YrZWDJcIj55o3R38GxDVEQulpkWIazzn+LReYUa/eDilKJDwnYor98oEiRZ9WRjY5vQXc1
kUWvNIN4soZzTFaCuCRsyXsDyVVAp1ngBbb6JBEoVrUi8NuaMr83q7Uxr+Z7TfKiyzdr01hfR3XR
GkQkE1nvHsnKp/IseJxMI+yrT+yAEU2i9Qj94piIrYOcV+CG56fwhvQ1J5IbLFCiJV9+iAO2Kiuu
EPRgmqc7cy1BCT2aIf9Dy4f6h9uPOQ7pxRL0apBF627POc2eR7N+lBd2rCTdrlowuSdEish6Sjdb
yCY3L5Qg2hJYNFjAX78iYXAg6Ysaw1rrm5d8q3iBOh8P5KO28nwVmMfqRSJ1/XqVsXMoPXelwcIU
4yd6i0yjfFbKEcYRtamLMCiPIonJZaIHVXQcf8jTA5xN40gqS7DZVQc+aVyD8bcMQGmiFMtNOG4k
a/LnFM25kcGGaDiBozu4UiCVSji3H5qy7+38iZMA22LnR4fD4tT6g1bR2opjOJuc/oc/0TZdwTVI
AWZHsMm1jNmMpY5Czy0urFLvIUTQTnga+ngl80kwvr95xvhGLgcraFozjvourOys44boWc4IjT78
HabcUzf3xxIW0BfSeVoYHotoOVYmTdxXRgaDao4s9E0X81p9STFuTXLbbgcEMJJAYJ3Wb92F2WHg
7q96s+ubXN0RhhYFnkkXyVADH33wd94Wu084skKO9Z+fBx0JBQY+lnk+Ee5xoqA0OORX1aISfSbJ
jeLv+1++n4tn7pCOcm1s6J/F60gUj7bcV8nU4nzdRP/EGIGreL5mPNXP14lHFYt8T9MajfnDBVRx
bYPOmyHmUStAU8pepe4iENZU32dBr8aPVhh+59U5+v6k9umJh7LakOVOiPCOUafYIMzzV2YGWirJ
NP7+wLN6ZXVvE5q6jbQtIqIclV5lCt+xNqg0zyULMM3lVSNiuj2DKsq9wFx3TvKniZoAcLbyf0K9
2IAqNutthAd/jaZeF6XVGNIUz9BMNddrEoI91v0kk7mmJFN7JpkGH3pRmnpOK1oukr4qREyZGYru
PGNmTNEtPniviyLH87mbvO3XANE3fSvfZBgbwrfL2vO0kGyoXA+l2/MSIC4XrU5qhewJygYwetKw
WI7VeVqQhKdHP4IRKHlRp/C+nQ5r2fw2JRKZcvDLglSPbyc8kNUoUetOhsJ5UYNu1/IC3JLK03+r
pAvR3V5g5HKC55hJ0PbhKffyhOjyAKKJF5qVX/8q3cvIy7twC9XVtbUH+5JXHPa4civ2WiFS0rbL
2H2a6mLy1q0ZoLuMIh5EysZpFZFBprQkQJDS5hV81RDSriTIIO0OSEeOGsaiJuIfbDQMDxdvU+Jq
N0hGnSqNQsKxpWtcKy0PLZzVj53y5HGXz1Cg/hYt9CFbu93TTZdslh/kix0nMgsQsndtq6Q5wGeW
1U+5YgVL9FB3jw0reqEnm/IZhJ2no/ECVQ28F+I0On0MrwQMnaYG1bwYbmwFDBq/gf3hRpsBYnoa
DmriIsRl63ICRL5BpMQA0AuepmwPeXy/fR3cuXrvLjcOQzsZrQUBWGzI9kcTyrzqVB2u4TsuTdJU
7MO5pHI1ao/EnoXt+spXoKGWGjHnYUf3GOYuDk19B8cJDn0tgS7rBHRo4Krugy33Edu8GFtZoiHl
1xssgvdDIfJSi8/4/EYot93ytae7+QVo7+2X9iv+mqw9Y9cX5FFDIyZTptwcXjryqaxgmDDiHoZx
6OCsF6rUTgQqZs5JWghNcpfmo4CaL/uKp5FEu1drVscGjSCYaivbw7Zy3Yti33oS+DcHt1Q4tZDA
jaIXyOJQBjrZNajTMnS1MFdKDtkiBJq8rw2rCLvt+N5wfzjQmW2owSGTd8Y/NuvcIxKSLxDiqrZh
pYG5tOjveNP0uPYJpXR7Wj6DevGp/A4IebthvCH1nytxI7gUZjNBUEw8VRBDiF8CY+kRD/AL34Ic
ZDEaW9CA5dqsxM+31WilMVNRzNn8QPyELZzgqfCqNA0EOiME6ttwdYcMaPxH5YKjapMxu7VgLO81
an02Lk10vIeAh5E/QLziMxMkTMLMk7bvIN5DTw4Q2DWLOEkAIshm/XZUmCm6HeNuORyA+lfTX7Fm
lnsoytNhx1TpWEQlnIGVERmU8eak/kvoN+xxaEj4ws6+CtJnSS/LouTnp6szQ+XO4l+CMkUrxnWZ
z/RIgVTeI4Xyv2LbHzbo7R6DDkT1lcIboHrp2ihI7W4jyzfCJBBbmwoG1jlc7+I99tij0xjuurMY
LHO4xmR38EwuTbFGawcwe/alOfBrYOtBh3EUwRGuXXJKC2XdnzvWZBFWMSfYLJRl25lfFlt21OIr
GcSfph3VfSYbApYCb21/Glfr3F0FykrK+yEKG7mEU7ZUwMCYZUv4BKk+P5XPTybd06/odwLtvznG
LiTNbumu5JyMVG7Z1l5oOI6M9xECCZvguTJ1y/HzLfvUoq3BFbSJLqbrvai25s3+1dfztJuExQW4
zlTgXLed3PQ5PNfX+DYh7WO71dotIc35Cc486+UqRYQj2XSqzh2nBeFbvP/qcLi/35uuntyD9gxY
hohi6T0q0Xv8/38VY8YQdlhlVq1JpygciCMsxIlIuVN8iaL42RY+kkvzYGphtwxaWxdVRke7CzqP
VFA+dV9gD5rJTePaF4hm5N8CrWBqeofS4PIaGiPKEu5356kxHNTq8bFq2K5t2jFQdEcumuEa5mvC
3g5+7mVL5caiNp7gY+FhTETPod1jI6Wu4Ox0TTE413vb2neM4Kp8JE5K8KLG+OQN0B7gsio2s6w9
6eyJf5NRIULwfrI6XqfMcS7J4O0VwIpIX9x3JWCcBA/nPyDbGjcJpWmF/7SzTgFeORhQSVSM6I2E
0qeQXKLd9s9vQ5kKI9RK4li8IYY5okqSHpegfF3+LgwEdNyoKvpSlDyLGBl0eRzq1C7ypoOVCZHR
xNFo/WplWNVC6eUrgTsQSzNo4WfdfNhvB2AawQZRAjDfwTp0pZa7axa/VN6tLjWPX16FfS4v9GRZ
L6XtAYCyRrXlkT5twks9gGKeSRebU2bdl3kbpewANAF2d+Ka7OFVl3E4Fk6e7P+4jwPhOFPxSl24
+fLdiErLP+dHuSgY+S+drjp+6vlO357Cuek6oqHy5DFTgatVEbHOb/imZe0RjkOkshUOM+Ej+tLP
U320dFfgX0QEq7zi/k9fhi59Rev82aFgTSvZZzgnJsvyjKCCavEPH65pvLQv9bDUiPB9VhogIp53
lWZ79IZRL7AwRdcKXYuz1pffA/Bt61cWdmzusUb1/t0VCRCCzrw7OWRY8j2GvUHFaidHxzAnn2S+
TktTdTxTxQuHTEb+ToDVWRT6Ld+4PoCFOHZGmMbnu7H6U9QeWzwcoA9bX3d+P/to8i8EiulQS4az
zwXajzwxzc8ZXpFXC1HQlFBlYiu4MhOpGwDblxAZ+LmI2AHYV83kwdXqHPFMASvmnOxZJi1gvmLZ
9K1WK9olCq/Ng3gRevOTJ+GgD9F9FiTqDLbEDKAf9qWn5mKZN9+yVcjMZTleJ/tPDFXa/aT5LUA2
1pRrcc1lekxMFcn2YGYK1umTfufjjQVrynvVJl+BbwZC+OfXqzwzAHmleCmVGhPlkO8Khar/mCT+
MqpubedJG9SY2OhH10/8SIbU9w0xmQk3JlGemHyGT508FkVvHM/9gKsJOp0MHpJSral/3Shvw9Zb
L6Cy0Ife+I/iIQn9cmv7fgZ7rOCnbHupZ/GGuv0mASL4AR6ZsSdN3HhczbXLkxPut0CX8jnS6GaI
PHdkq7v+Ng96i8h+P6BuC5uEzF8725uIRCXCpRASfaNKChoiXdQA49Hs8CfKPKlrgbmYvlWFhkrd
C36xboinneRXvgwpOozJ91ljzY/pvVdjQKDykG5WHOtE0RqW5vrnhcmKLvdPltLkE0s8zIuhY6lp
3qApbx7byXrgcBsp29y3h6FxVxUQaQy2biyCLRb7QRbbBjpxiI22L+sQBiUxfZt/R2Td0xWqn0II
OCcJpJN+kUTrG0mGF8Y6C2i0NodakCEfn8jJHb2pHr3CLA69gJbA/3RQWf+spXPMx+k8hJq51Iha
z9pd0Xzw0XYtBn/V/puJk89/b8YI85+UUZv/1S8ZkHEx9rIISdrxn6XisAbdCGcHrI7oCQzws2ZM
Uhc/bMPW/57nskB/X2ugR0JjvbEd4Q5mGpftRZi+51aXIV7384FECisicyx43cICCVEHBd9qZTlI
l9oodwSZa+uIGXf/ncjbOoEQyPnc3NvTZ5qkF5QUpS9BSbGfetU+D6nsdsd+hbj37mYVT0yIcV8P
tJjC8fh3+D3RnsGl3kGzZePPP54UxuS49mthvIQAEutLAjIRkmfGJguINLWmbVqWhi/OyJ6J7MH0
ZW0CwB/FMtNxTJsNqsRuIRbfEp7e7HaKI6wvyLTHjWolOK4d1rYDgfP+vMP71Z7XhyvhJNBrx1jb
AORlf4a5D33ounOp4UQPpRGWWqkuf7sqQdiT3mmFuR1aph679gNkYkcCePEguhpaIXLWPMkIfGjT
c/2iKhHOWQRUwMiCmGW1X8oM1fQFOW9NC5w8k1aB06oKbzIzS+OP05b9KjlB5JThh4bWTzM33JxJ
5RBT8f30DLHz1HQdOfZFEqhnOJt2qKfhCoCZHsVsRn2PCn2ZrK6FGc8r47cinshSxD+68YaLsipa
qy1EK7duCc04BZzc7HwEQ4N/IX491X+rbovOJbZm8uDmuUhFOlzpWNWnZpfP1qRlii+efSAdmQOs
BkCpibXsSpZEZznEuV9VzsST4SDvVBDSK/tYyRAaXInavj8ybT8/os+Jy8qOUnulEjzK/Dvfrc8T
IyFc7UEy6kmZxa/PX9ZdmODlX/rGi/3iUIhLpLlmiJk0TSx2l/hYfDzgzBbIDlMwbvq81RFt3fC6
ZnU6WB6neHkXhSk7NJKnpqaLKHBiwAjB29MV9L/DVS1L1ZIokIWThy6fuDCFdD+U/EAHSpJeqkKj
b6biiPm33XYV4F2BYdMacQyA5qBR6C9svn+dxg350dxbkxgPwmowtZ6ZNuV8r1GoeKadfnAC/ukf
VdrAk6M3xOf7XFOEPT4jtEG78nxXFTswUIFfGsGPf5NelmJL0hn0gMRgqF5y9Ws7CsOfjrxgIS53
Fvt8eKIxB+zLx49yM+QwPqvv/skCirJtq2dxBRRN1TpKqescabPv8cHqGftaHJZIg80IqsVmmwcK
4KS5CFTVqqDixWLYreSeppZH3/zt5mHWT9u1iPdRndafResQhw/xBYkJS8vfrJiqP5zAcTWCHYep
2IryDn2HOUgzRY8DNbDDszn9Y/Ah3QHjRVbEUWzsjaokk8el30aFP2howXBLKFmSnCHOhu7JsD9y
kjY6IVR96Uo03TSC2WNHJHwTCYI2E/aY/2ohOdqg21G6EOyRZpIgIFw17edQr9uzU6PAJf7Q/bYO
S87tdHr96q5pK9/4m2wgdyftBSDFh445lyj4uhVkAhqbCAz0hTX8EnEg0SPv+1Qzui9LBHFR+kN1
R3udJbpl0GemTIpS89uqowjFjLnScA885Er+XSGXAqwY5NmEnzJGwVLBL8Y8R5PjmWT9njfbPY1x
JEqiJ6SvBVeJ/YUzBuZ6cvj572cfwufaE+jsnafJQ5PFsT0xzLc4Kpbou0I0gyPRiWTazMqS4+D9
OdvIn2eSwD1np9gTfBZGDRBYYaIaWZgRJp3XAJtmKDYNpqqtlryCLkbwzZpNlTdJNhJHDPPahLUv
tfFIyTiSX1ufaHohu7eyAAASwo0lxe1Ddo0Z4uJw5LnydBiuods3tnscTXs19pfRU1IiWNkOnKEt
OmiH6vzpUsDA0567rA94ZkyYqgNyxlligBInj/bGl0C7j25L/WB/9oELuJnmt7oMyXEGxQiz53gH
mFUsFFmPVS3xwx6xm0vXziyx2cribb844lLTUIWn7kC1EWhNONk5rA62ehmlDjqckn53U4P5QyyF
A6rdJ5BhpJ0XTXN/oA/iFithbidP0GpbVSwvAFhTsUgSwPYwZq8fe6TOva2wralyU5Mgm03ZQKMR
jludALpGS2OBITfM56SaWqhvmAyTZLRPSCf7aTMnDGqgwyaDWep1VF8S1JG1VakmA9TTIveVoAcG
pJgSHJIiGLH7xUEswRK6O+WXxhc4xmM9hvAXAgos9UAP439x/0Uxaz4Ix+QiyOBrP0qABJnB/D87
O1lEn30ik2Gv+2pDx1QrQtkSxsgWPzCFu6qfaqV5WmWH1vKLG34M9KfWgl27y/R/bzbWFiRlobHh
5S2TWfn2QA1NX+aRcsNLAvFvwm4re4vEIfXrRcUOS6Ef+TpEn8W9y2s6ouaoa8UzeJsv9HP+tX9w
LL6Zbcu/NRoNakxhaTNIk83vyfUk3eLXZDgWNiewGxe6Q7G63OPzU3DVDCuEzWUstX8g0RYjDhGj
CHI6Yq28Ef4IWs567++bpnYSMQy5aKiQDzEptqwShGNPq80GDDi929zSMhhqrVxsiD+cXX4RCdcv
nzEdZ8qeat3DVajSQfse6hXjC7tr4YlU8u7dxHNB0guvhFbDDAxCUCiuT5HULHTHDxlbU926SMwY
BhgLYqHJ9BCN9EvCtpZMqQJ1vlN8qNvKcbngWVFYT2wUwSqfUP53hdthu3iCcRMGLkemnTTqA5WY
IoS59wUioSRjLxOn4U8AJNlx8asMtCkOQ2SmhVoVANeAIGVgDF3pfUwacpt1UePQtX7rbFCa3Odj
R5uxbzRVTTSl6zMLZ9TgGQLIV9UTJHOBETyMV6LjP15vJTYkyWQmpT1jkPai8znMHyKRAvPQukgS
NM2xYZCr1uR0QSpUVI/S5JtvZ/bfitAAPe2KG3XVen8oNzRSehIUF0HVdXMSSZDRsHbbsVy39E00
F63OEBf/s87xQArIn46OcLouOkVNLmtgkcXkUg4uhJssXBLOOJM+7NeAb93bt3IZsEjCIqH5x3vT
nEL8NXyMhmEvBngLJKVbhpnr1n8DTvzrHSeW/DfRKwt5pJKSCzuzJD5moBq3M5JIXMSCEoX7KZWd
eL0t7i1KyOW6PNaE+uO4Rc0Jq0G55KD7FtiG0hO7JvdfFeFRrB82iw+dFaYcw4BjUeik7XuH3yfr
1zJECbXJYxctY9X7juC0Z8QG9yvZ501wSW8zdmMBUOyLmN385z/C7xJIZNRcId6fPFcN6P9n7OYm
Jw454DxihDOHnAYVinQI0VAjd7fVNqQ6/8ekHvLJbr986mZXCk1FfgPeSyQnewQtj4MggBWPlfoU
XeFhfPXyvjqIKwBlg2HDDGRmuQF29QIfLfkYO5k/XddZeZYl4iZ7rYPhSSKzHcEYBRd3EF9MVIwV
XUqGHNe7C6KPsm7JF+lmeRjh4wgchSqaV6HukWU7T2xO8k6sV/8SIgyLaQlGiU3gxYdqYlkmzou4
J5TXSsQG0SuexqrsoORDOqmuwUc2ZtGWpxY16k0AlwvYXZxvyB/WySh4SxNwLgsZnbH457zjFAx9
ZUqkAuWncaQin+x4HVAP/Yq4rSKlJpvUg0PfmZWpYwYPkCxIB19edzBGgionqBuA+WGyQjkPyrqF
VUANQZrEZ3SP5PgqivuCx64w+juNG64alSxrDmVfcMmgsRgUfxTwMfXR47Fa+Waawy0PF/CTym1a
BJ9G+62WkRBtEXhwJJaLFZcpSIDEHynDOe9WBlbhr5QFaq0RCPe7SWMu+ftVgEQ/Pl5eclrkqZNi
QgDpexub6bC3SKrNZ3MmnLhxu3nKKBrLKtQDwKklqggfqF1IadcheQhdIFqp6hZy9GR45/jU9jjR
gooHJbgj6+nKJV0CGbF5ZZzXJPPAeK/r9CsDmLWGThieASnu2FaRz/krs8QJBbj690nEDnsv72Fl
pwJTm75JsylI+gqNoCgkZVm+XK415JHesXoOQAKRH7o6+yOwj5A2GJ7U5Nl41YM11PCoFiD0FwTa
ry+jHH6gDNdoieaDfZTqq/K8zPL61yCnWSKXeUbdFiLhJKpq1qex4IC5NKRFvFW30kcl1yUdlnvC
Xy6niztq7VggOvx4XfuhLVUrqxbc/hN/R9Qx7nbTId47pWtq1i/c6hzcJtbHK1hO4fV0GKuHdmZG
DGlGlcJdvJev14AnKvFoC+AbxCWVrHAAZQ8hyJoDqsTcHQ5CIbknDmSYJcndEDFGwViW8D2tEnvK
2fKcLXnjMNIpHYPrXwe2wHRxQ9+uWhH8c4h7PI1vcaVmI9Gev12Q6tCuBtiI8MMp28Aq71ZM7qF7
vJs6nmPZm2o2nxRZu8NuFg0CRAk9JFKT1jCou71lxo1ACmv5EnwuW6QuaJP4TkBiDc9msiUss7xl
fqIQMC1OPBKh6YH/sqECIF9+1b66/Db4mbrOHSNWL52JjrrZugInnTt3W8BWm/6m5DMfEqFZ9Ua4
py0C9L8raqYp70gvjOdPsb/MtDT2b3fSuW32wZ5VgMVFvnRoA+u8CsVcloMpa+22xPnIHcJvZj5Z
A1Famzo2CMGh6QXyntm31mxAJFANX/7YDbSXRLc35L+3nnTupEmLo80UxO5t1icBjIRJz3dU7YzF
2fJZRXMwnZfNZVZWFLG5rPR5epXoEBaHZ/7YV0l2TLKyxjp3t5ml6isqyjybf0PbGxWrnZhI4+X8
cmJdjn91yquHcA87l3pifyNS2ZnSSYL8VCRVLxmCr/ArK3UmM5EfakcEBxOv/qKsSSLuD9r9Mbvy
2h159nAJVPnPY0SGQbClIZz5aeweKol3xui78XfX54sul+TjN6tq+vBJe4DimySuqd2Bz92EHoz9
JtS/aFpQE4zb696vcLjPvY6YaNddVY0ZlhUW2m0yhcSpYdRraOpyZ2ln+VZD0s8sJen284Syd9BO
pnu0p+lRyTPQ/a0dcLnHW0lo67zB/yRme67sQOdD4++/iyFYgh4rVIcRpAa7Wxjx22MNgROXELIr
x1ALN1SHGLj6bQI0naYiCJMCh1S38DTqCaL234IuJUEUK24mrTXrzW2TlWGyAvk9dAcJnMKGDYPl
vaOF4w0ofrlK/uC7xMdbxii3aYQBv/35+uKGg4bc+gWVsbnf8xSjJyuHzMbHtcKua546+PNom9zR
S2gwlXjN7yzwLz65xYo8ODaOP6TX6GS+wYqPL6POOPc/fWUu1bidUMwQI0oojNAdj+weKdbJq/N0
XGGy+9036GDB4RcP9kikjKoFGccYQSH5K+VJ9RVmYfSTFuqImN8ERoygsbD1qdNd8c6Qnixiec3/
gdXMTui4Ekyue4g1qwJh6atAx2N5mns2kWqSQZy59QJH8v9/Ng194Ow94Yj0nDOcFtBNymFgt6sX
wtnOcShzHGEtV/1PDxMPNM+xbzgwDazlaN/TdaMMeRUDvMMYfpyGtbv5t4Xb7Iww/Un41Wp7QWK4
76pHPJxPlGWRcEkjv2H2+/eEqlZUKgoZnZIjZ+JzscUnDDmH8zKivoPMzN/OmlNkiAEvnNiVzHZw
6XcAZ4ni5kPpMsZRKOCdOn04826iD7GwBTx0cUyCgdT2J/Jnqgyy6lVciHSzSUPQ4AR/6hRHSzoX
DS25SNlKi9u141VzhqLp1acGe7XNNkMSjmdSkdUaESOcQit9JsE6aaT0JthWkcYbAAUdlkF1QVpZ
51FAjyWxyj5Bv4gYxli0kGhSfeAcccphG2BTOtIvrfhmHVqJuxl4uu7Xps9EEEFAPodQN0N0uc/y
NGYosRjeE5lIp8D3x9ZjUd3/qcTRmZR30qfaYqEqV97gtVdPlb7iU6u8Hse/VFSuzA0uSB4xmJJf
Rv9/q0q3DoWiyCeXxk8e1Xwd1k1WONlgh7oKvcpK7LeYKbvUraY9TDhy99fm1s8dH7/VjNc204/A
1hRwruigFUgEaLwRJ7uvRcS6XLP5VeBkJVIYjqi/ldi7VU2gkpzU+q12sBpnlNf1Pf4XerGZH3DE
ycyitA6VEIBDKGHvxi7kUTl2DK6DtgrHCWXA/m3gxNch6m3Dmzhr2dPU2lvPd4ood4QkHE/bL1Fz
AzIpMRLH3XbIMSQhxPcSY+XtMLiZ4Y1olMNMUwTI6D/wDUKHrGk5+RITr/pHN/rmJuEa56xZw3Vu
GVUe8mj6b2eH2KTXm9lY5yIy4GiMKluDlhnQ4Cmc9Sk7+py+to1nmtJ7Xg58Hlj4w111oxHxBBT3
2raEbG0P7O6oNmtXK1FVPQGpu3xiwsmisQTdOhFxxVnqbL4IzOQPkLrPM359ci8oetLw7BQvQKjK
qVcMv5+wE5cUj62RvDx9FOvK++BRigjJuJ4I5leaNFBhm4iASyakAgrC8264iYNMc+1tlGkOFpVb
8wx1GHLIS9MvjYc63omnEk8yMWTdsfL/06F/xqT0ag//N9LidPiTvXwm5IhCeuUIVRcYw4oQi4cP
4ftwGJmNe8WyVZHP6i6hjRwnCWn7VHJWCRt5wP/iVf0RWb0CeqomPTnp3NCFr3hifZMtPDqDFBSi
myddsU8vvfAkO+/wZ9r8fA3DrgZZtGTVNbjyoxpfpMiQKCaBW6KKq4xxZAx8auq9EB6mHffzf+aZ
1FXP5/MFjNTPbOgNntlLxi3pdRgaISJJYgJOIsQmMpltMZ0e38HYacbX3JWhj30AZ4bXszYX7Eha
lccTWY26ODqaMSxKpJT9/1YeQclL4GN7iiO5pyY7qP06JtVNp7m7ReXj/Q17OMFAXUbxYJGkDkeX
ibKdeZ13z8OEAu2+EvF1MYCYRNlqIbMp4ipzEVTmxzy5nnVYUgeHdEBtTSkmbuKXjDxUyOFrjtFy
iodgHJhJIFyDpVhV/gG1D3a/V6HVr6T9/Ach+7A7b37TdD8/Zx6yGp4+WWONcqJtkVm33fvHlmAA
BOKy45l/PY6r5ITIV5PblLcf5hk4x8c3yrHKorT3KQ+LzH0MTLQ/k5E5GGp5YVJQ8T8X16QnGpGO
BRmoJ02jOoDtyEoVyjwGYzcqcZKSug6j2OIc4Fbn9qOf0818eitz4fler2f9gwILenkx10ekFGmm
4q2yYfWCuTfpO3jDT6MXiTHkqNRqXOSnjc7PxTSScpjgdVimYRCrDRegomZ51qv27OhMyL7xbrf6
ZW9Y57f9DeaYiqEHgzzEuuhhLsRxsPXLfP79DsHtEnatKG0Z72WFfxV/M5B5IajrFnnc7HrEyeNa
q5G4oc8CpXH6JkXIlmeW1FVA2CxK2teuEG5Q5zRXhcFUAfM8Z3U8znhp+eLhUVtV7vfxNUQ0J/Py
ySKOEtFIf9MA6X1AlNYYQ25zh6xTt/hQxMBQGpS5bPuQ/Aw01KWI9EcBanmKdami+g028IJwFtQ2
rm5cvNUavp8v6N2IKzwCFoDXM0GEb4bZGc5d856HSIqT+9Zz3NR7MrE7JL/7mesgPwZc1liHSnQA
dLFzWwx/WXRhbDkZKs8xTTO7jlZjwPum/n/OMEFKHh2mXnWwAkYmNiJbAqjjMwUUjPWQID/OXrR8
U3Ad8rYmJqtSQTHWQqud9/NhSZL86goLXTbXHnIp4sVhvNCSTxqtpN4enTCpcvnWG0Hux7gcpF3T
z04VGjqy47S6EAfqufZ/vkNJuthHHoVRI/MR2orAPbi8uMXxTCSWk1XB13tJ59YdjOiVrBemfg6c
L2MxsXICepQzkogmXRukr3MDxB3LDSF7s2RQ/7e+h9LNRakIpQWKBx2WFws6C5S3PsaONU2EHLZK
CAatbLSoYOiC6yfFt02JANUl3kMIhLtz6CuL8rBsOISCHDz14v//8N2x3Afq1Pm2k9YYeeTh8Sj0
fAIIeil94YCIreC0qoBljRzOBdPan2wx7VPEulhMPeoWvhR3Kg1Ha4bCuCTD5C6J0rBb8Q4+XFe6
ix5krQwpDoOF/QezgKquwuGKk3fCkSPR4iNdN/BcMahZsNnVu/P+9lRQNQK+Cxa8pFNk7ixxfGgn
vkSwcRAX75KibapaQ2QiD5/EUB6K3ZraGDyd1t8GrmX7flWI8aZ74jtegpxIE26AOmHDejMz/bPM
K5/IGpXSA5KbaN/tJ8cgBShYmlR8iiU7f7xaP9jEWDYCyjxJeYMvbuPxE+zc+Q8N9k6jqCny/dSw
NpOmsGWV244ImFG8D3VzWrOht0a38yRtmjVAMYRc7QShUQnX9Ul/6CSIiiOupojEdYjunNji8enB
Q18aR/PKfxE3Ybdnd+nlrkwisRbGKnTrHDYOuAqjpb5jlasb/Ig6GmGK2PfjUKzJ2baBCpGIMfsd
gtbC3zBj+89gepOGjtHxsuxe66aE5TqRug3RWgBriCnp9ZYyByNwSHs2/KA/LIwUer3ayehwCwsX
m8JUA2uRFQUGYLdAat87F8h9CY8g/HlCTAoDnzlMiqbKYU7upuy7L1XlNeNP2jAyYZWrGThYxrQg
HRKC5xHKjajaPwrt4FSoAdUfmSqsPDxfyjNHw0FLF24viHx6NY41M0pTX1Oyp8XMxhtE0tjbxWD4
v5Lke9fUuKcUbUNytBe92COTEr4pKMbJVRVsQGRsFcdeYL3BLU1JOh6wyWYfnUeWyTORLx7dkQZ9
VNsnCsuC0IGiA/t1+gja1eEhf42qc/x2hs5oU5or99dZZNqG1FKsnXp+x0eegfODAHRbZGPlQbCw
5xrcNL46nAaZYA5Y1XZqsS/1RRDJ5fQ5Au4WaqyBrAR3SEa0+oOny7CD8awuZin2RwxpZw2O0yYO
3IAFA3XrVrfIvhNu5kJVGlunQI20cTWSmzjvfR9LHEiXn+COTjE9GzgSpDKS7anlCSH8UQv5jsb/
Ar2iLlCsaGBPThUicY5DRHTmUAOzy9whKk7Gk5g2OqRZgU6XmaN5cWw+ZN9XpkEMGxFOuMiT9Oxj
ZjMGcUaH32TcCWVnXnqCCI8UDYMnrdJVqFLKC8zKVbGrsjJnmQzcmxx6aEOeSmULvspE1djyQ7ln
AmdLpDUBPPUoi+9HZmCYFbntOAR6yHbdyFOCvN+Meu/6/biZYEP9eKgD8iz3EV67UchJkVAwbrEe
DdC3aCecp3MKyMZdXBDEIejgt1FrVCCwKq3g7nHRtw30MdHCPaJFq2IAMLe8dsywdwr9Cb0USnxw
bFAvJZrAOmzdIPkQd52gOpacr2GIAALrIorSJlp5ar0sObKeZur+plhmGxr92euiKJ5EgvlebRX6
m/9p4GEVcOZ/RSHZBQdufmWsnDY7KRuxWCZ2ivm9CSNZrjPr8u86Y8eUbuLJ7ZC/cqw5K1tJGD6q
SOC+zYZfVjWfw35N5wJtnYonWSk5dq2ja0LaUbinRZYYWXX8HuD4+nmiX3Tn/XsQtgEk917HsfJO
uG94tZBX3BbsHWP9HA/IeIqDcBA1tlhHvMvUa8mKMWBqlSv7NI0LIMJcghwbHHVu1A371a5EvSTn
07Da0bjiftha1th6xEx5Dsrga71hDzXW6/swEYyEcLvLkW7yVW1UD4Fgr2rjL6hil49PrwPQ7xZn
H3VtWoSToQrUADNIl7TLgrjeLk0/uVm1gesZOagGJjIi4+qn2VHTg1XglRnsUn+bCXc6JDebgoh7
hJnlt2YWC1ecylQeR4nY0en1Av7jqnxGFwq2QVAHuwnrJ3Ld70L+g/HCT72BZj2hf7fXm5PJgJy1
16ZvfxIrZ9fh32zlbCORpMjSVg+327jj2+nm6I4HG6rqHpn8ULmtXVuBYzHN7eLHNVfY4R2eKimp
L0DOAo0Qc3AyB1kq/RruUu3cOipwuPdbafZg8CZlef/7fDcVPPlTLnO9ZA4uvPCd3d6ksleraxiq
2UzUGzRlmrC4S0jzqsUyXzUiW7+TdfcIyWOOAMrvUFif3QaO/CF0vKRq2uXh/oPgScJ8HArAoL++
Vmb60o2N6bGYaAo4RuSVeLWM/vCUDwGnbIK9K9kZ8h2u/3iRuxN/OJRYfZf+4CSNSsAzMDZumGZG
HazaWi1AfXAbu1wQ01rQ6gNlydEIHQKXj9RREkGBIzOsi4AVlHBBmO/TqukCoDWHD8jYeY8Nc+yZ
YbZtIM9wlncBDN3ovzf+RX7yN2J/sRpfLA92NqURK+Q5ULQt60BrZ+DOEVP419jtVPdITNbJAJ+T
63rDHNtJpjMLjJllFyYXn2IrtyV8HPI2sXlSlPXvS23O2oc0TRE8TJeZv5D5DDvHd5YM+NgvRftZ
Zrfv7baveHGpsRzguJ5qiIWCb9e4nBp9WUE2kDoZy5mWU9/tivImMc1XyTj/wmM4S/Y8v1+Pe7WD
131iJoSqxAQgM/ubdcK+kWuF2Ybub5jpfGDAyCATZYdEnLfMpT5znKQdsGmBBDO8aB8UOsopgzeP
mqtzX1LAMd8i/6zb2d8ptM50zyyXFIFPcddqo552dFiGcx4VtOXJmNhAxAUiy3SC6UkyrrT095Q2
pbjt1a9vnu046q6QAhen5oU4LSwnxyBglV9OOx9ILTNn5V5BwyQYWZRfAiCoQGrNCP0VsnF6D4+X
C8nikIcTr95dPVIKSDe2HkFrf+ZuLtxUEGZEkZWgj5EJZqtoVAlaUVGZbjlFOsPAewrlvmkGQ4mN
80Qp0645qiCrN+f6RwcPFhXdAtzDnerMCh7wXKwbVBt9Pfcams5my3oQq92U7+iB+PNWd1sBUPOD
kT5l2jC3Fja4+83ALDUeLxJ5coVBBP4bl270zUuIwOjDqdRXprerU6Uo2Dwg5l5gP/O6uOrsa/nz
Rj5sujkIU68ZH832mKbXLCpY7J5YWUtdIp6X/boCY1zTzZMBpoGPv8A9fBI0TZRsky9LJeLUnID2
opVBs58bD+0NijB1jCKTYnTBWU748d1r4vaP672NKL2CFR1IqX2n8470KdfoHgdftdoPfElpKnBg
shrqSHb+A4cbkxyqMrO+GWlVU29VzJ6veCpipJx34jA0uaGSrH7YjNSHsGA3nm3g+xNnj4hF+Pb/
AP9G270aDdHQ8nov5P9CVxTv0WHFlz6kmHGEYmT0ej6QlyzINPWuzRbVelbCn5iKntixK8KJh5cf
jBVlLRhnMaOIrUsQgvvj6jAPD25rmB7kj4rK7GKYKnXRX/XbGLCEVgqW6mtvtWO8ysPo3xF/mIQJ
+wNPSEH/6Y2tjeohgr94oyLpSCFrpSYH0nZC0Cu5A8F6nXzYHT1fDYyt7l736WJ3pmMtsR4HGEWt
fsrctpQvb9i8v6Qz3ISeShcYajXI3WWI0IEhVF37Qix4PrttD6YTTHZ0Z4aQ0OrJRTW8MQgdWico
prOrymOWuQpN+/rahADy9wyW3kWYCAJO+66XUO7gke1wp2scQY6Uw7rt0aE9s0q6kzwT5pzZ2EbD
Rw4ycI8kQRZ6OWFviK+P5wcKLQ48I4RinQ8B0tZ0gBvn46c5mjBGfEmw+6zhjzXOAMJXNT5UOmuh
BZWVrH0EbAcqpau3TPHV+JmzXIk8VnRA9g2KizGbOJIFB1Sk6qAotS87Qb6I0SXrkLNDgMp8kGYW
HjQNoeQRELGgITVrurVWAmCbjncgX+qu0U3DY4gZfj4OV/DlOsd08LJZZakJ7xfUwqIZEUHLrABz
S9fhKhxKHDnbxFl/mTAsBRYrnn0MiL3JVBEYloMWkF4mVGE6xcdKxGb+KUlJkiBGCensotCsrEv3
5ltfIE4yVPOPEeXFyg9s9NIOfcRYa3EnZ2j69qUmo4mNbh63oJWSdmO9txiQkzWOyNrPbk8xPMmY
Tves4uTyAPM9YxEmuItpqg2j9jN5RJGLRa7mbBs4zWi/75hxhQZFWNvTGxa6qWhTjbK2ePlxMXxG
bfgxFr9AQZKytuBkH5JYx5zA1LtCwVla+06laMjI4hrqpYf+084Vbxdo8gSHpIkB0Q9/GWl0jIEc
on07eujPiOXNVrmwMPtEXnTH5MpyXKNXZgZfoeMVhL3yQyYbjZZuMf0zJx3G5IBii0FqvTIx4Pzw
EdH7kblTuw0iucOBFPPQrp9WdsOVIGIOwHbFDm/hMoSUqwr5PRyjROwQxFzrrYnLcd0F9/MFHiRl
a5wTL9IZHYYUl3g0pDWxL5RlJx+mzVsvSS7v+ehv/jMQ8iL6ACTdzx6+7UY565rqVm5PNDE5EUAL
eUMfnOwtulksCsnHzW5A2JKidO7MruoFeQXgF3gDx3jk+e2tJWEp8Fx3xJzJfpKnS/KKYAGtxkPW
1nmZCZrmEWZud1qOfvMQ/hOgNqUvBRtjgUN4/uISBnT0cPacRFCkgqITK1H2LT+rwCT2WEDl2hKo
/SuSJkbQbeODPNBYdjTfg/8WAdxLb4f09t6zjoARE46ELe7iWzEdim7lAvbXJurO9tsR6AAll4tT
3fmqvQc7slTs+FoP0qq9O4M99jnaIk7tX16j+PTZP3I50MzdZQgJzDhY4szyitWX/BacNTPSkq75
Vnw8CR+hra3HFQ43PZ/hIsnLdUBHnlvXjgW61CTVuucbcne/iafphlFHhPiBI5rvknBaWcVgt1Gv
N0WyTkknLejtcLh9LPaCh5HSZu8hd0rl79DGQA+9CtCZofKEX9peFO16Qd4sQrkO66Ze2IEpzEDa
PcemjOezb/6arHhqEfN154VrqZ9P1TRmbkUWDn+c+qGBtl4Tru5HVGD+n/D/PcGFFuOG7SAHXjnf
u0gUPZaqUJR3A2sQejSIP0cTNvDpVuEVn3J0WKk4/3JAG8fR+Bd8O7h/KdqBQ2rg8O4KS5qhLFIk
GqzJpwy311jcbYT1z9HxVXlIk+NkuWBGToIY284+A58+DF/VAkJ4jqKazceOMUR8PopDKrRo1X+C
G2xI8V9t0LnGL6B55IsSJSQepGOTM0Ij31mqeGmDEb/MrmcBCETlsT9hNde5pegFXh9UuUnk+w5G
rTTPgudzz6x3vL1IRA6gCmBp35e23t6+Qo/aGqr/cT8rwnAo86SbBthiZ7O7MoHSSCJKF7YlvyrZ
mfBXRtBdO7+gqEdUDh3v8dED9K7l2OOCwKnbNC9Pqgr1N+VzAP3A/guWMoXMs6qTFeZumWBXAVOw
awxhnL4DqDcvmfos7gu7lW5vREnX9Apr+TEGD8McXY5y6blHKXq/NORqOrRyrPH9WCDh9Dalds7g
oqVnMB5mV3haNCb6IYIiC2Z4XlVKXKcVflGmlgEUoC6HnpnSEDWrc/d9KZjsETVNYGBkN9WRkrNT
AeGNLAcX7o+HUKngB2ALHUCQwYuCxkTOeYoqrWD3C/fT3FJQxUV0dfWvTZs5ZXphsqQN/p/ZjJv2
9ZFn1wRLEV34la96FpzlcjKE1/SxlA+8BKUZGug3dMt8izFHk+a0+Vuc0ogpVz3lavW2cow4Gmle
3khvEEk2I9XNlxcZDY3+7qg2VshpaEQjZgu1z0D35FxAh3MRWRph/nSwdTm4GHnfTUNUvPPlG+aH
US1QONMZAb9xHTfdJwJN0Cs0/P+F7g27wINC7DI2GZ2qDAar5bEIoaswNVN6c3ucwbWmuBCaCKwV
Fa8p4r2BA7bcr/qysYnK1EH6/y2PvNVfN9gIYlvgGg53PH1cycHfbDr6H0BPEl704h5SJu5KYTPg
klXczoWPHQPcDd44hrJ/cwHlwzT7vP2h1KWrFujiXYD08Qa2EZUCEHllF+m0BKIzeeUbLMqWfCtE
5rvFzmwqvLS9T+PPOJPRSVyhV+FRrWCDWR+ny4/c9m33BhmyeraAR22wohTZQLvkYkmSihL5yH+i
CxnzFSCovNM4q0fFnxnBPvKuouR2BTNZW8fWTUoXHi+EHyIKHBkjZSznYXpf4QVQwTvS5GGQFgGY
gQr8eoi7SgCBJlWJWCdEb09Emx8NTYJmM21qNZdMl3VO4RCO7CKP76tTEm5aauwdBXRjGTdFAeRL
MotPfM4j1TkjEFLf/XNrbjBL9SFmBYkPYiGye7bZSGRj75W57LWRmTiPNnqZpSH+2RoIKxBdQ7V5
owxjQSQuNuD4tL97lzFa5De18Oxr0dKbivAU/Z5qMViAToYcRfxcaFWeOsuxcweR5+cryPQz65xw
85ijOdezFUhiuOrSmmd4tjuQnTODim2tQ63dalNuYz6HkBfKKGCEGNcn2M8J0vgQqZkW496MKH54
jumZNxPvf04S6f8YGZOP+guBBJDVQAutZNO78MSlOTnxhDVsyC2Hrp9aNukSe3MLOO1Fbd+9N9j8
5/7eE5csG+WnHAVgFVhZPO/Am5WfbHsu2JeCJBs2lNA6VyPZEus23CnjPW8nA7I28lSeTpWPBrtt
FKaJS9VSAKPFbOeDk/R2BzssfQyCIc9F/CxLBqERne2Ma4CFBOV/yJ3O2JZ6pJmNdTFanvpho3Ic
wSAr5kBG5LL6O7/As4pDOhwUgU7KFDMUuIgjbI2Ke474k+V8G2UecvSwKZfiNZGMw//JAdZjav99
4XOEF8g3irACPWQRaE0vheJefp3iI0LVExVOvE1am83fQ4A78M5sLJpv8YvACAY/V66mhMg8JoAx
MDxvwfUWmZXZvy60MXD+axDNwLd6CxIwsjllrX1m9lVU3Bj73prSHTN3NZ4hsRr17ABFeLKOQUdx
6uqfBcGsjOUs4EMU9IBBowYSs9ZBK1eU5cq+KLKhjlGSuzWBvr1t0LOMDpFxY/ZasR28f45pj/xO
EAUOjkF2BPSf1sVAi4VustsKTII9ZivWWCQ9Tysfx0WCdOxX4tBjSCMKHmK8mvLyKWqIYn7CuYXZ
r41k5ttmYeIsGx6/8d0Sv5J9u0HzttMAcFcJKpguZJ1CKieDqkgNRR6lVDHsFhBE3n0SedYXuOdW
3sn7Ppyn1s4BOvYXBT/ALvowTX0fQtBQT9cv/z02dLXDnTQc5siBk1mY3DehKdP4fSNvw+6b11nP
MVUWrw/avkeIcJPFHd4ajO0MdpaQ0h8JjfhFKWmqMi0zrbrPcVjsWL31B1opblYYgX5cZ84IWqx4
RaPOQDmXYjwRY+9kZ2J87Tq2aH+s1fuUbxOWf7jq++Z73Yhp59cE1MP7tSoJsJj/E6YRAp1Y/e4S
aDO0s4JLHa8jYFxQUjlmVCZXzWHJpE7A4w2boaTDemX13tLODGGMFyQGalDZylNNzcOM1nxJMVWC
2qLokxHsQrLrzXYholSWLebQNW5SVXVXapEJoFNxjr5eI9q/ploTVLKcKMeo/OSce+takYyhn7+m
tfjR4j8TNY71No77mQjh7bTn8lDbnXkqefL6QNsWv1+85zG5CuviR4twKO7gCDQK6w8NjP45z2+N
IrHApdxOjpiLPZLblSZmxF7jO+wiqUbBirF9R2K5pxpyc/jYAg2lB/5/jj1z2lI5Gm+RDnUDHHkQ
6BBfL1Puju9mwZx8vyONHnOtesm6vFR7FF0RBRKewJBQwArdbEzkVK0//+rfcNGsKMYYjkUB04JP
Rh0canpc2tkbPP6aG+oZWxVTicCrXO6cm++VuGmkfRkSR8Lo/SpQnuS6m/rOErOJbXIJ0il1rwrd
pGZmuJgvvij1ARKuIrT4Qn85uV76ThEJTFYivUG+BzOpPt29bWsazJHR24fZJKwgHVsCzqgBNdpy
AN/VSJEYUnFsRx1EEHQTNCgNLHxmV7HPoZQD8/Oc5sCWezeShTwWSUK2zAuMjnpuZEYIaSOKc8cQ
shJRzotxtOWT6jzAuaQfaPpxytUy5vGYDfj8dSnlFPk+oxq6EFJN2BxDlWfw/0hTIRJawpPc0eWT
cPU3QNK5a2aZaORt12Ei/rTy2el8Vfobm81WzQUPXUZhmva5VmQazeKhPGx6aWbw2oWgatl3KRdz
jESocIwDok0poysutCXZX6KsBGgA3yko99JvJ7oJedqpoUsRlf/gmt3n8YuRr6FAlm2Rn+STwUS/
F44sWKcw7ylwTClaq4/TfQkaODFlz92kZIWm9U+wMO1PLChNVHj118ocZVBktEIQrWagFuZdFoV6
gYYKGFTF1trs4wSga6sbfSf0VQkA/dU3jpxJQu7kFsANcpK5/xNYLElkQA93Wo+vBbT8n+LcijlV
uQpowmYcHeQ1A2uYmzYJ1xzgrLlr1NSFJlNs9oerImhWLOimBcsegSv6PynTtyc+Xox1NuZp/k/f
S5/le7OUJqcvooHwgAbZ+02N2VF4PlxYPo1qrNct5b51IU0aVeq5FKIQRXzQoH4PJfEGYfImoaJV
gsg37Jb1XiDy94RMKSOmRkj3WKhe4LZz5djNhZkT7/To00H03jerOLaHaogTy2ZemT/Rt2Or9vIA
/1Dq3YY3Y6bB2XeOcg6aM2cjWOhssrKIxFmoPOhy8V2tiA82O3T525VKVr40uUVr7oSc+ZuTAikW
kvygbdFzyo8sGaW9KiNXsPGOPPsJOblwRocU9fIYeOCIE23WVPEDCK2Vulep8GfGrlPAho6DcEPh
xUaBmMpcB9ErfgCnXJku+t+ntTl1+hSQL+u+A0HxYd7GEUAnt6OZPnHQRPAccarj3P1MOnJy6Ofw
hXXuqI/W1cH0BO3jaFKT2rdHVru53rjOv2ND3nW8HlAJAUdeIm7VBiWuSm1xMufBIuBu/K1h1Zy/
kC5yy/psiZnlbHjVc9DuwualQoUmYMV7LD72vr4joj7421nZQ9A/rHbO3TKUOYQ/qDsfpWCECV2I
NNG/vh1YVuyqphlKc94gQhzWS3ENKvyB3pUyKJ35jAYV/L62aJNRp19OMcmj9NEoS1cBt6RzfY/G
btrnf9EvUn9xGLk0W/XW1o/KPlWkFDz0t5+aIQamPqwWZgWtrYwDJqgrXO68YoXVvOEh9KrX4rif
P/LeV/jJUmT87zsMkCtnJ8Q90yjr8gqf/OrDWVxo5lECgAZyrU5PgD/Of6/T3vIBIhiTLBP2vm2w
LOeJphnD5V+2MEqAfM2nfMGysBGyNE5lB0NuGXa6BLE3RUk+ObMJ7gIwocqZwhu1oytkq1kLvQw0
yHg9Q/t4o9kSgPoOOML00NC8F66Qf5emyeLv+A4cW4OzfrPb5k6XlQVNSFAXuewVc41WsYRsYdTg
W9e7478h7dQ0/Ac23DSNALwERXmEj6lNwEM4LUWoyU/J+uCLWoSFcjGnu0fUfIznukrAIJMaeL3N
f91qTAVwuGhC3/afDQ6sWBw8xfjqgJSV5yFgG7wCJ+Q6FitFXJPPphiqxZqOx7IthB7dSE+oeoiQ
MCSMrMtnJOmXi/rwzjdEom8vgYDDhink9GEqb4YERv4KRo/0bjJOBAQJjF1ByE1Gv3OphYzq2PHE
fosB1GlYArpvTmdYCosAAQ8AZyjBiFsCywHHIKkGuiSwU38abJiKYSM26B6mpUw56uNpZRe5Bcbt
sIAS4BSN2GtPsxYMMLXLvTsrueYbKPfjm8MgeQsSljDYVhJCcDh6ZnceAhw9C5CGejLqwFmXDtde
KeiIBXW2097YkgIqZ/txscrYQ79oIYp2xWNnlxx8JF2XYqp+WtYdznXxriWsn9dVasMES097vEjL
zKczrw1FQ6b3glFIm1WdYpDlDyhLYJwyb4/60dRKFrr3y5UqYmmkGFRLx01j/ql3oX0tnztKzvqx
tG/jdmLlRofN4YxsOS48Nr/Cx8l0ozmwBFh3SbhvxuKQzIi4XubF/5yKHS2B5K1tViJpFNTLjESr
CmB4YuX4GTXJaqncemrucNkr38nXTygpmugDTo9tT0mz4i00/QsTl+XQzeuZlOqUiP8TkWBFwVIy
rjuB5qG3ivZCNeciNjGnDYU7Lyy17/fxBdip4xKDYE3owJBt6YVLBINeAyKoG0FebgQFeU/Td0IQ
g5NFYTS0YHJceH84POx28Jse67aIhR823XdgwTrY/m/nkL8OR4TKHynumPysSbhrFjlLd8GAs+53
WYKjWCXtR603KMJgPiyqR4mikCRXd2bq/S6j1gTQay/h9q7fXVzFB2W6QGCH8yGJ9i6TOoa9MhbS
7ZLlYX0kxPpA3eCL4wm+bDqxYHx+30aJ0nUChPGeTZCxp6DOFU+za/Bj7tP3itGRue+FFo44kcmC
kVO8o8ePKL2YUeveuxbHzDiDbSjeYTjQTdFprURVfHiwRQEsVbMmCtG5VbLnAV/b5FfdzL/gii0v
UaqvGJCzUhU/qgly5PUHOvgVhr/yekw5EhYeR681vj3DPWFjZ6X4b6ZWRKkho4M/v8Pj7b/qu12i
YfAPK28OrOFXSAGDxTOxq+SWz3phlePlqFQkOo+RsWNak2GM+lMaUIF8z/D1Qa2GRv0K9NmN4nyx
6k4R2+xrov/q6mDYBBtdW+5s3tiVxGv1v5EscFZPKq+oOJ7ttF29HOhZ8dXs4eZxU/Qw5k3i680q
d5pfMwz7B8CzmgLioh79MayavbciYgQeE86ImssVq8nw+sGT3IFQjVnUvCjDfC4clkgS0/dHImnE
oTumqwxHqGWRUm5i6gUx6n8CWZElQZM0W457hk1LSX6MQKd/AJQFnH4gkIb9FVvXzm8sFaL8iLV7
1ooRjPPjMTtLZAVPkPwqgJvVtMesAXvs5g0P3ZMGrSIL2xuBBOV7eeP6yw/7yvQnLulRhuVQtWqn
d2jqFR8K3ce88hyvbPWqPRgfl2O87q5IPkFTOU5A8hDBqWVlP2yNDdjr4pXl/7EDmuE+/+EPYlqn
Xu11eO2752qCdRaZmili9GjLxObHueJJay9aXvjmx3eGpdDnF3b+snjQZtQ2yuKALzE2fd1Z2qF1
IyF0PMr9W8l2vxq/opWW/R7c6ZUNuOgAvAvtGpLxJ9vWQI69M/W+zsC72vsbrmWq/BUU5W/M+nMb
UjR4Oa8/xVE6Agd0JSzUlg8sLzmAnA7guUVNK0ugVc8Z3RSHCxuey47upylnHTl3TKvV/5AQTmkO
CjG0UFHz2Aac7+tdnzbzbtluH8Q/1nnxCKzjXYK4o5xbB1/JMPKjwQc8WMyyOpxZ8N9zgQ3CdYCZ
uJozD1lH+AwIPi7wD1c2nSoPxGyFJx/gpinfTztRRApryTBiVYJYGvNmd6F52TD1LCaf+r5F4gg1
baSkddHzSipXnYR9FvvdAVicUjVFrortzJdNs30xo9umM3d1RCUb8rukwIpOptyk/i0BfE2IXYJa
4/OqYrCGFvcg7MMjHnLu9Jxe7rHAgPX8CLxFyTvKaPsUUrcg/Hf2ZwtJZEIl8QugUb06TQSuoZIp
SwDccu84WQI+3reLlq3rCyIiFIBW1WWx2rIhlkwUj28LNOMtC7or5GZDhsFZo9gI2oFi5NiLTL5z
iPFmZBoBevai2nBZX9bcan64C/BHpf1RDNePQfgl4ed2pLfvp7OuRIkbVMEEqWj+FlORXxJFl8jF
goNVGTN3w6RBCTAPz7/ZfSWn5Rjk3vEDACgq3Iwvb1L7KXLX8eS15gmxUUmmvSUjDjkBnpDhAF7Z
nrPuCHAXaheRX2h1HhYTR0hkVC+lCqjJ3kox49BGGsMXNJqO5mW4lKjKLvBifbe53zcKHFICZuEM
xDT8lWyjKLJjq08Tgdw81TURacYjLX8jTN87hqvHktkt8FJhtrY+eWyVh4HGFyKvgoAbYjtQmSW1
A/iEivsireYT8SILs9avl12NGXScDxLFxgYvCjJHPooEU5TQ/cKJ9MVO5U+ZhHfaY9PPnUBvq+h7
5OMvDBQkc3I5ZMGKlg+PnnQJE5BP2bxKUuaTwI1Pk5wbvfKn6JYIjGu193NWSXLRll3j7e0ypH1m
0RgAlEZy7kf4yutiQ39zV03TBo+EkMJ51VqtbiT8zCGUGP5I/i1OKrKl7y2g0OiN+EAyjjNUZUF8
gL0WyVBWgaws7iKdhoZAG0C8OdHd/IvVQNOPdXkwNIEyLLe9se0iGjCnBkxMw2DeHLvaSyMxXsjV
TTAKeLDa55/XTGJWBXVHKcRRJL17rrOjLU6CX1v/rh3vx9d4l1L42YAOtCOPCJaLnfleM2LCd6OM
BnNuWxBNBtnvsVZTrg36cPKHwx7WD4mbxph+X1jcplRKLFr5NA6EGkE4Bdwoutog3kFRb7xagXOk
bvYKONkR7YNMaClr+2X9WO/JgYjKHYNQ79C384p4cR3vosbbtlUZOue/S4y4GVUF4l1lz2IHCv5V
8ZvtmuVzvGp29BZb5v8lerpYBsO/PiEaJfGpwOGwfzdFI9Vz3sn9myIsAX+8MFbdKZtdVWvDeUq4
mKakcOzaY1YJ7zclz11oZXDssDqnuLN6HMyEd7+9GRiixk3uM9Vvq/NToKbPNwa++BARr48qy8C1
f9To5If0qTdx2BynZS2ve8qcTDlBU8PJYHdk9alMSql2T+tMj/oYdeICLqWKhCUl0tbtQFr9NhNp
/XN7WzIFGvv8hOC7X+2kW6u9PbiGrAibHQW1UFCAz7+Rvpxpo5CaZ0qzfTYfUfFJCu1kH++bCaKc
+D478U8h0bajbPL9MInH91L0cSCh7rnuq3z421qYPj0dCNMaR+YGLxm9hj6eoqRsW4kGUCe6WEMo
YqVSFzSWyanDL6YT7gSXWXtnSjGE4COmhqFbK5mFT0seikWreJTxGiJm1iQgd48SddnQjk9A3nsa
E6pORddGlGqYPcSkkX9BsFTr/fn7e5f4sjR4OcywrP/c2/zQl/75xeJ8xvXubRYRGe6U9feu8iS3
iPYVj3c51xc4VUCOtn6eS0iVwKdU3P/A7n62Tua+rOMleM4yQHWGLWdhc2kzgZML/0nKbkBjc8NW
Y05TonPKLG37IRtytEwvCRaizDi7Mi5G9YEUecfPYxx50FuH+TvF9WHvv6k1TSRmcjZg5OPixP1O
4uYoUI1pQ53Zggs/UvRgEQR6I7Gxj1CQqXCBxO7ulU6cUR1wbFpPrxz4y8lWUWiDUoNe4E7O8eQ4
0+e1EJPa2OYLm175e1vrvSBSnqQBH8hbjL1J/ZSehXa9+G7mwOnFHu9+O6zGXRpEe01+wbnSi2Or
/443UlxXGgjnpe9YyXZr/Uyjvvpa9QJmzJ1dEyK8yiMeEbz9n9mg6bPhJ8E41rlNkgc4VRysFKOJ
pmPlKhuVQ5P86kxvaUPXvPYVkEUW6sT6zEGzNbXP+rmVC98PSHaHof6ZfdzbeAQGtvZOWztQG/dh
LEBJ7Ltcu7A9CnRHIL0V3IHx4QuH6f28m1315/crn5+hk8JspqbfFntUZeN9u+Sz/MYdVl63W0OL
Z/rSVbASmjldo59suibCYXx3wPXMpLOktg+W+pOmTb4B4NgPJ5vfznOY3K0fGxWaFtmuGGQvEhVj
O8tbGQ/Rdcn4Asbuqt6fIRb6PoDLpaIUCp+f2Ivjs2g6szBqUX/wKAj7ja7OO1CYCtWzRyzH3Gt9
pP9CitVXwJbdp7wXTkcH5NLsILxN14pP05OZ5og78OuTqGQa9qhSA4+KOzHGs3OATIZhkB5V6zQC
4DHtpwSNv0ByYGbwBRH+zet7SiTd+wpPoZe77qmz8QNtVH8RbW3fDvFJ+ojJC8nkXXSjwCq08rwN
6CtAp7CDXcEnZUKQSjiMl/SRJTJ594N4BLuQulLK58HFmtEQ8+vKJiAGyCvgB1amqCWw3X67m/6/
+HVj53heLT2YE7l+2rBItsjom32mXIoT2CoQQtuslZfv4b4ZwcJCIP21m4FLdlbsLuJtXXBj+3sG
aIYMkQnx0mUb8dz5rpiL1TzPEschCyQQr2MKW2DfLhUqQfksxZJQk7b+0V0Fe4s9si7Fm4PCEy/E
ot80emBeYUMbALmWu0ycDPaPChNSNzeBNJWGY3L9lvr1JGoO8lG3wg35D8bSRfYu3oD6L03lh2rB
9cZlL0seyP5B6pa4Uw5Vbs8XnSu9UpuQpnHFOaibNGXvLa7D+lqqwxYqwRBUa6d5CGHusaLPz+XK
yK5tSAUSFBw9YJmOMUFDBDLZkXj5H4nIe+Om59XWUq2OJhxBsOMHN502qL2p8P58W1q20JBh/tL6
IK9ddsNBCc9kmt6F3maOFW1ix6U4ux5fmyykWnHxVLy7MQXHphoJqpuJ3jghKdJoq8RHm5h87tya
Xadun+FlXco9MZQmeuwFlupi44lN/CYdBUunvxuIdLIh+QOu4rYTptXHKovQldXmvCBt/SslNH8G
7H0xfWhv/6O32DnjXb7g2SHyHIf6W+qX+y8a4TPT57LScQgftotGrqD9HgxNu/DXS4veojSDoXK8
ec4m0klbGKSACYuf4gYiVQhjYfFRjhDBfs/5z6jrbciai8KRhbXijDuxzEYlXOuLToy0F1wp5W9Z
jKiHDQtwo2r1DoI2bOVek9Ckg0xDIurHCbtOu3EoUV0ojE/6inm1L9zaClMQIM3zjBthXHXDB+eN
8w/++g2YZkjItqk/aMR2bLkhmdW8mvmIhJmpoSk7udwhW2Zrf05ZjWcBGPPvHaz1+bOjfOMidOfC
SxkIRYxsAdml6Rwz2CxemDxTvKiDTbb/fRECwroyWL2Ii8iDr2DC0UiNUBQfiaXs1yNgB4dSZumv
uU6tuq0I7V+gcUVT96UOFCidKN7oXM2WjOi6v6qYtRTWAYC5t4QpgVrODH3DlEnxh6WyMj3V1JIi
TqjAejGSVXHQf/D0DBjBAk3T4trljvU0hqXA6aAt/juxtzlNz0dJNR9CTv2uAB3/UE+KzifHK6lD
gGAA3BGl8CHX68UZqehNwXv2IZMUpN2GfG4uGHcUuBNW/cVpEdAFaQmyuPWLD3Xh3YB12+ytH3F2
KlK2Wf8k4QTgmengqcxJhbeBQAMbVwR/z6Qy/LqEhDqoiC3/405CV+XEOTt+A60wFncs/rqGnBYs
vWTZwWv9o2QeTGroV2rtjNXi+c3iY2AELtgPiC0tkKDNePY/o23fH94ijjuUapQqYkY86PDZVbbL
mOoZFtesxNpNyDla0QB0ypH1D6+WXnXnZ3FOge1BXfb0XK2rnoyKu9PTHRlC+3faK8nWZvD2rmxP
/Trw1XHgSGfZ/d8h+WWe3uLLmeM6C5TMNFTsjK5Yv0mCa6Lxf6sJN/epaprFhRRh9LTEU44M36Tu
943Mni2COZa4729OeEQ3PJaSBy3j3LXwD9fZ2kZjM4bgUMceXiiWzwMbgTK07zlL4zlO2HT6Jg1n
GgZGZvF86oR56bPkLk4T0ryKS2JxB01dxsTbIO7ugv8cR/aT54KwkaoP6+d+MRwFNsl9LCh7nLQh
28CNei0qafyfxiSXpj7K0uVc3pcbD4RX/qkHXQ13m+Yp4fA34XunuX74yZCdnvZm8LsBRzjjnB1V
gI4UAJH7ZectPrfz6R0fQasaMibxtmUlPpjHDPvCvsbXAqx6tL3K1N/kNWSnuOQujG3nGqveDAp9
nLbw8AjaiJSQKPDTd1qUNmjpt8u217a+n6krCjyJQgglhceAerpjoCLgGwYA+sAefkjSdjC9ENzl
ZlbbeHOooE8FrXgopymfjBYQUSO53CpCjDZgmtCACPWnwIwxPZY6IbwHC/TFn11gtKuacuksNLYa
0lK2+R60z+Uc7ExHLiJ8BGCSw6Pm6dp8bRjkT0IQtNF7kpKs1Aki4D1o3s9GTl3DWzHvsMJhG5Jv
W7hOXMDh0G2aMRBEqMUjWRrmNsWHTRuHmM4SJNM9e8wJLEeBHtdNyXA5DcZMAksIR/rNCmFrTDA1
BPw3GK8YRP2tnXHAHw7RYxVUgnXOe1bSa4aXUnTRU3sMm0bH+LEQa0qX1GPwDmYPY4ayMEYLk36J
yX+t5e1r5uznh11WniOzBtRuMSkdWcIqKhfvzYuEgPYgV9V/G9RVNbukyRQfubXMf+Gp8EgQUASu
EhAbZG4eS4NLTUbzCpJN9SYMHlPKnkGsCcxnJeBCNrYIcFNsN2/4Bu4ERjH/BEi2y5tvamsFJeQH
UnC7jwCsIXFHEWE5g/P7CfiGEx9NL7jHA51/mVuA5Z/qWCtoai4EcGM621c089lwP0lOM/2sNoDi
QOEZsgV2h5pndxtZHFbGu9pPXh+83WBGwY5t9xoHTXne0+TKUEgEDApxKpQnX2dnWP1tVibj0CMh
fSY2Y2FQt1h0+gKp1LQ/p7vsssF2ZSvJxHWQ+MoBQ+O5CH51utA9bOh8Aptj8wi71EZKWoExvK/t
vuN68Wn6j71jjByB/GwK4+tTsal50ZOqJ7MqYuLidXjBVc6MDzYDuO9dNmliEXk5a9jHmhgrAu/Y
FAC7HVWpzthWB540cZeQvSZEp58R5v0MYL1fADOrPAGQqLe34Ym/bsA6CLM4bYw+JfJtFeg5EwTT
h8bNcOLcvLTtlZmIiuhVNZC4EFdyrUrYfCvT56JnPxpp5lDhcKmhdm8iAb+tuW0RvHXXzyhgQlX8
vAhXTdZC4/gjpOZCgF9kCeyP9Piov0M1VpRBF0prdnJtze/JMD8E2UY/8bMqFdQOpJtm6JOalnfz
YhRdq438Qywr0KxT37qF0zt02wmSDpxdtnyXEnUoD0p6RfFHsF8v2SmwkxWXfzGt1eHFy0pr7s81
9IA+IxuJdXDGv3PdoP7JrW9eDaSeyjQDqsyYEZjWFzjWRb56hzNYPPYgII2t4ouVdZOD3+gxvUUg
GpqGuQQ0wHV8fnl06Z7nAX2ndSbZN2XgXqy/azlbqFV6s9GX7hEFHi1QXP8oeYSCd2NKLyI3Ztjb
6OD2Nh1dDytDG/U9x2zT0DF0OhovSodOeVKh1hCHwgBov9l/Ftp7i3BBk2aY9FdkTQaHhfV11eTq
wAAzZ8SOAZCpMylBl7rs/3QKQZ41zfUc//uHzQ69KnUadhXfrCiJauY+6iHrVnLLik9jQjJ+LS8P
0hWgcBTlczi6u8GkTr2VfKuvw3aPKn/orT1jVGPIkosScJR/CKcpdEyAfwEBVhr4R/LqeMnPo5eV
EktCvdug4DTIgzT7qRtaLX3VrN+JUNpu9C6emIejoXjnX2AQYmjXNptIvuObEk1bHWNBoCY2ZdiG
rDeUSqZEukNvZptH0jcSR0Lq9niTYDc+gFUbj24p1Fq4cf5/fb7JofBQF70mjBCG7v1aSoTywxXd
lhNFnPQKYDWql6XB39WwJWgdQuI3ZOgW7mzkpt3omCLsHrL8fZpiLIKqdAkpGlJthIcNwJYpNFUy
cPr2jTb9+rnqkOYSbQXxXdrR6xYMkiKBjl6Yl4Ta+5AfqxQIXVrhHN07XAm8CvJpGXg99k1DZW0K
Ds6gDAL9fXV2eBBaWKjhtRPw8VQ2/ouQ8QV+wm1ofU1pcmEKFNzbTXIxjlnulLJrDDXCOWDGwspC
nFJh7atacn/ifdJfoA/Ih3AI4N2xWFnjvHK4bbXc6fWKUlleBiKlYU7OtSDcdgo30wQQi/5bF3hO
tG77q8j8HpbkhNkYCkdcNli0LSbctA6WgHwdKdSyFskyPbGHbx9/DwAwGheIareBOr+9MusTxc0i
1MoIgZwx81xKRIsTpfZkw1oaajFY7X2Is2jrFVRzkKTBj98njo8b0N0vNDEC5GsVqSNva4IKKA+c
7+cQj2ggwl7ov/PMOBL+XPn49JWvYF9981GdpnF+FrpqkikdLNu0OMmyqwft3fuT9lPZCN989xBL
n2vKnbH8j0vSwVXJWN6YcyUBFhB1Il4BpGrQXL5yhkDb7DXMJAUUuzt6M92/1aVOopKtTfGKaltp
4Y0Dy8pCN6UMjDhYKyELTvKDIeLsbbm9Qzv5r5mbNklpJIkPIukuafTguzIaLVQ2O42f82gIXx9L
IAfxiU3IdukwQj1sAxXPbFzacp5yCafz9DaUD+ztpxhCICLhEdpI4/QcetIV233sl+Zm+zD0ShEj
RSIBeoODSqU0Pm+HsXnFTRmbwupxFJqQWQyOaKIFfEG5tyLhTsq/l1Ew6HxcR29e9Dob2lZzHZLg
zTTrBgarCkuujHX0pvdL7K6tbRsYr9+RXHWEe5XKgAOQYOaGwl+Rg/NXDGk4tGkPCvirBiZbAooX
bUe/fGVQVEEt0s00Y/PdK8maXl3+7e5XYIc7D8o7fvzH14oenE6QAkVPr7Z5Uvj1nZF+gI40h813
+EiiY4D6WSynHIa5UiFOyvdn7udEjH/qxBMO98IQB88s4uGO0VKVGdfeGKYOfCAdqvGmG1eYG1YF
xUqUml1EPXzAR66XZGj9m2Ozti8UCiyH34H5z7G5lRZ15ramRH7krKY6zHl7a4vZbuYoQCfVfwpH
2OHKIPBeimMWM33hjsmUt3kmj9Bx4wSHrSfJC9dCBJq+XPrNqFO+O/r98Lmib1bCYTB3Xc4l9w3t
XMBBudoc9YbXkO1339onR3h+VDNYIRTYTgrRv4JZptyqUNTMA9mbh4qqhWbGx3ZQR8c5TlvbzwJ0
c0Wq2l7zAPLMvrX7FV6ssGh+yhRXKF72pwnrApvfkxKv18B5RCppXhMqsdcLH+KWFKPRivZcHyvi
fgvSMu3znmRFrOjx85BN/R3g0MlCXb4bMI84vVeJQQbVsqe1DQZlHvT3ombxY5yVkRGfQTuc/kDO
ekyiI8LLSNXYgyvrMuuEjAFCHfgdgjtt6oxig+7Ow7zFkcn+c6d3OMps80BWQrj2mGdxUmlR2BlC
6iMuSeKSfbtlIS4XF360j1UyY5438rTJIhYJ/g8Uv2WMkZgVLKqBl0FSW1TZUccqEsymnk025S3Z
sRVsOFcDWCmoc5y7Aj2mswm7Mb/fi+yFjjg4eltJmIVXGQVwk+pYgIit5DYdgaShYX6XgD+/zYDm
U4RYNIDmJv4xqyaNIbmsu69qanbQEsXuJ1XczdfnI3ZIB/trgJtJqH+9xOfitUU/BJ5yXZK0GrwN
sQo0dXkpZqcqDlHbijxJUalGUl1D4TIUu5O6UcdMyNMe0YfNC2ar8FFBCZNEho8MGCycT4CtcNpr
A8/ookx5ahJM5G98dYsAFrnFTN+ZLuVF0ruup9tpWwklPOMVbKoiyxBNdUE2cJoWTNfvmUrrs8td
ZeIru0s5fpgg9/i7n5cG4h2ugk4HWvP2ClZm236POBmIfCbi0qKFH69/zGOqj7sq5CGxL+S3cpsk
MDbFXNN0nErXdAJgoQhgVhXusm28LqEj2gWOAOycL8Bh6Ih+C3isn6nSYXcAmZGJBLnd3mrSiGFc
6ZCzJKfxxDP12uBk2/8TXDaRxYatvA0IATA2t3ECoswDYXyCOj3gYGeOz/XG4yGKVXvU+MAUjrCt
V6f4DeuMEDpaeiO1SuNZBWFjzqR9vOA2fb1BB5pztqkxfXPodWQTCDfiyunJnzBeNZunNk0w6ETX
N/jUtd3LIrvU9WmdDtExY80f1h9WDzAq4Is6lVr/F1Guqznz6EQIXgaqDR/h+6NQU+tYF7Bw39QR
1sS1CwGIItzKF1J8cJI2kfU6Dt6LdZumkUohKTb2XAHfqZPJzAMZ5wOoHR4hlYsOR/R0z7Ojos1s
TtvCzJs1ia3DPZ8TDfD+vT3u4NcF9eRiqiztj8/24j+2DR/D2v3w6pdE/mMv/cKW5gdQPCqWaAgd
QtezFzBfxrMbIVCB3V4T9pp7hdiGvJBWaEn8iwH4jEvBnGf37xzQCCsOdcigVdTObyb3tdOjVh/p
SFZKVUdgPk9Sz7I/OM5cvneaydNs8Xb2nUn816Paf7GtGf2LWSkL59Z620nxVRH+OV6OAJo0VkyF
6JJHn9O3Zvi//LT4GxcJNunV4OLwfu0vdfLnIxdm4rzldD69VE/afMaqNbdxU+ZGTs8NBqFAsOCo
9Gj0DvGOyoymEJpLbjIjzhXzG8h+9kg2ROcDlaMqUWIaBFSF8GqEtaiP+20NkZ4En6cDAP+9foH0
kh+veGJ9acpK+TSVlfykgDUOWmB2nfnqsqlgkNyK3rHUUTvDMtsid68QRrbjlGkZnseJsogs4JUb
2VEKHuRNodFBcc/0lQgWQk1ZYCpFxxeG8cs0H70xmYMDDrQvlZZczuScTyWffU49q9b4ss+nBp8x
GDa5S33N9N1OUpddZv/aHYbvuisSVFk+2313LzSbuVDLcgJjjqpd3zXI/MAU/nbNOR2HHzMn3Eka
v6NXnAQgYGtm8WbUui66hmb1FGGxMD/VDr6cddvimU9ipU+8xartWVrVEOnHWL28mJOaKPd1wNjZ
tgzoBelIL1h3KihvuHFC9K9wCTcN6etcp2CgFRIfvHUATJMTz3baqmHFYH6sHzf3VCwd3OTQrMK4
tOLp7O/4iGA7I12uI+0UxP/atc+bAxueoIplUGQ5OHha
`protect end_protected

