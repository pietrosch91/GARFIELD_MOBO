

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EsXeRsPajYX/YxoQaWaSSiCwfBR719VMFy+WbPGh2UU7Kp1+dfK2zv2NuQUxEGnYh2IsgOHOYx/7
4D14E6T+Iw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fwNmTuDBeFQhprdSkaRvfqp+4JN2uTi2veIKP9lTdMi6V3vFfJL2e26ZwNopnqXVxORqcIxB7j4G
1obXJPT2WSCL/0R7vCUMg/xfDg6ZfHRQ4HvE6Q1qt2f3x2eHE9gwy6LqEJ8d1O5yddIUz0vAxT3E
MCeNfnm0nCRZRRRR1XE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kL9kQOh4E6UtbQ/npzD9A5qvkaHmW4Q5TOqEPVqfbEiuDvKyIkPxWrP2j08vuQIG/7EyOqE/kj5s
ywoJMmW22K+cqgqvRYX4CWXFmZSBkvNI1XANVHol7+tm1Q6zcn4x8jo3f8GnUuBouEp969uv5TVb
C6W8kRmH5VAQXDtD7qgbVeYKswRn/GOr03sH8N9Ixf3ujy/rBmCmzDHZAfpgrSzHpSBDLuEk/POo
Xr9RNXhKMiY0o/UKBWTOczhocmLcg0NMSjuIOOn231vhyhTbXXcQqDAcqV0PuqZO7OgMM9AUBcta
f5wQBZ3NAv31WeWX668oqKgjV5YgAh+FAy4XhA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RtCEHK8hoBVXzxMIwgNIEMWUxUkR5Pqab6pK2iAMH+eKzf39R1Vn3oDa1Ljhrvx1X7iUngAsgX/3
LcmaDU9gqDte6ddNPkmbNLHvLhT9m5FvOkIIYEvIwBd4IBifYnydM1owSggUGKGtS8XQry6CERrW
2IwC+w9nzwdB76vItXdw1s4IymWgY5uwNq4//tpnCTkR/OMjCa2f6M9qEfWJYNlBJ+GXDAJmYmUS
wk9As7MfL7ue/D71kahi5ZCHlR1I+tDM5txkG5hGeVCdvwQTXth7HwqgDY5sYW26p5uvO2ZqvlfD
UgWjG10wynX2xKhSh6d+19vsIic1nRD2zh5zJw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R3wbUw2LtZKD3E3fbP2KygA45tQjKS5V6VfkBIYGo7BlcceQkKo0rH9dIS4uarIFJdlyweFapK4J
ePxAwMW5ynwhut3dqSMsEu3D/QC2USMsVE09S32y+GwiJIOKc4yR4T3A+F+DpWiAENZtryn6RnBV
jZ6etPI/ggwkkZm9cLyFuFK1/x6BNvCtmDYBz+NvlP64/yJ4zISqL2xL7EkNUjtPoWrn0H6hwsMN
LWmwS1HAvRjP69CtcKcn/ZrOsenLSCoE2qMOpIL4p9JrIN+PO8HJDrOUWtQU8AFS+CmCXdRF4XvA
aw3d/kbIocHUShnTob8znWjsVn39/MpEWEx/5Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NPgqApUBvoFW73rFSKf04YnhBIrA8CIHSiW0X2nssipI98eewlp5fI3AW8Y627oAGytBSN0EzSw6
6mWHpipQLQVJA6VeUIO+8/hOLRzTb+XgsgFpVaE2fLeCPOj0g3idUo0VTbgU5/uqesDE0Vbbrta7
T5odN3Lm9NJkl26/v5c=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ejAJ2cG07D83mzglv1+hg2mXZeeRNlGMZpMWRYKoOLgMgbw7dHfDf5ZV1yQve7ZbrKv4ydzeaMEx
8KfLuTCue4KY6+jlpd+KL0RPlmYfM6m/B1rwwR5ILj4xN3GdnDEXXsiMW/kLFu6ZLoD4Gg0fG+Vt
XWxnZfKM0dgbJWSRVoxq2KanJ2PlZ7qdlRIn3DOrtTjcJYuKzzGfxtNYdsTieTfk3SVn5bI2qSkC
3ck6p3do36oxO4wtfit92yihFVrV0gxzgLHMK4c2SX5FGVkm5jB2zgUjTl0KTI72iktv+yeDkEkh
cO+wtpTtK7QSUkTWzCgR8DX8WFsIX5CNO6bleg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
9Yak2e0l34P9sd0cbGGiabFkn89lRBt3aKXaD4Akwp0KVKKx0kc1uEGQaznoAFs6eiTTMMzbWRat
Y5Z7w5+aLNkw3QympkQEsHaSIrtRoZQ/bUjYmoODQb8rExi8MeyR5e+djZvAOPfZbQpLr/mKvIgL
I1/lQgzkJdNA5tVH9ez3l2LVEZTLXhHd2Hc9SzGIpkJ/XbCAAS2bncp0YCSsZex1hsEtDZ702Zyo
oxMbSGE8KoUWh3e+DEu6RbuoPGWMzhbVS5RyUCpae1vpQ1xYoRkqXZdHX5qe+eowhx5XwbyGbDwT
MB5KxnUXU0bIoRBC8S5SKIzrnhQfVergHmc1Pn4znDNn9fV0G3Pn9+T8FO0hsrm0NSQ60zE/+/8j
AGXLryEd/U4NCSv/nQGHKv84uqwFEDYPH3IPMHDv93vnch/tYXMSSrE4tg3s0CW/evnNRcT8EJm8
vOU/amYYwxOZTaPxL+WJSGAqCOJznfD48YfypxhRhhjqRv+GyR07Meudg2qxBOp6JzCu+5HttliG
wgyQqKN3b5jFDxbFAaXO/Tq/Mn3oWO3iPcYBVtQmUoQqKyv4LwzTLOtFkpFneLzGHMTF/prDTbgu
KCfrKFGnptV9p9t5fWv61NuKSUvh0QY+DOkZpUswH3ypMz+VIT5omVXqxZgAIurMSES2/e0uRHEG
6pAaPtem+/tsjGqicNVlAP5EqW1GIZRJDXMHKYg8fQ/YsLr6Qg7Ge0peoMFvbUVDqb0FA1dOgoLO
8SFiyLqrFLPNMa6TYLFbXykQ3FHbaJgegGhXesX26ZiBLdJB1Bp+GGCjYLWX4szbmz8u7WX38jTB
IprIx9SDZ/Yd1t/zvnJii4OgpmkoyuqoukhsY74MxkwD/Q5VKSnKVQG5xIfo+1jC3HFwij/rVxrA
VlScyALKNwMjB1+2E10BjMu65EWf3Ay60e//VokqK9Yi1WzAkrR4hKVwd2/ytCriVrqz5MEtgmmo
jtnAL09CEJlUlQXgHd4SBSxhQ/GZUnp7+08/l7+MpP3Dj8sVS8J4gQdY8wskDQ47v3UCvQ3yO5tU
MNeLzVwuKPlTW8/6TV2TS/evs1TH1TKjj+QvNgg7Xn3Mf4/Dc6WOSr/zLy9qGd+EYCJwPiu+B66O
9im2OqbOwfLsaPQSnvSaN1J91tLDkTc+johkApnG+bqymr/ypGeQFlJrPQhjMnECM0rrO/pcewo/
o0R3apj78eucEDRIJK2aqw8wVqQeOs53X8VvbfrBLJsiNMGTOwDUUWkBSFayuiVg2DfOdnKyR0kM
LcRMXXASv4si7IXRTN5qGQPbxW9Be+0AJUkxo2Laq5YMuNvCM2JHNtt7syMudC8yOgnyGzoMHyyI
nrY1dO1y/N1KFzvs+E+xyTVJcgf+6pGKN+VvqZZg7c7d4RyrNbPAtQSbpO2Xctwq4KqknM6+Lo9r
Xf5DQc2yeRZ5KBY7m9IJyTa2HNBseUfMLtbP403KigMfsVdsN5OZYFZ6w0F3Pimg0Az88AKds6hN
imav9WOSc5nb+yqC2IRK0SSvwi+in1nHoFPj8NWg8woCMfUhw9HWazSZMjYtPsOuNGwuBwbER7pL
PCg3Lu609K3FB8A/jSbHGBSlqrzsCOP/i85jYzKaURPVBqFn1wU7zRK3Q84fnVdnbwi0SheGh3Zs
ExykKoXRsX2gbx8v5nq7LvuvJVH8zFbm2TNb/nPa3rwKnV6z3K+T6aTVf42F3Gj1qMaMQ9PzO/Lh
f4qLzMr76lOSNOu7Scu5/YXfx1cSmbPhQRLvoATpBoUWlS2n+y78DzOAQH8B1uRXmF0X0W97bNSZ
RH7FQaKEF9UC96hn3o66EcoK3hv9qxvNojFTOKquqbjgCcjIFdJM0Qw76D3bHbNOsu4KGL+sOBKs
hBxslPrgfCYkrIbbIW5uYahP1GDnQ7v0fTBi9hd36vntzdT3Bf0B6VAGznaMV112oHAUCGCbvWey
RmsWHZv6UfE/jMsyobLZSvMGMLR8SADc44dQ9rrt5kgdBNPYcL+PcvptJNGZ1fYGpbIPq4c1NKmc
uraMTAljMFZ3k8C+Nyxu6Q3NQXTTDK3cN1SKmmAVoXcWL86QwRzcBqZ+f5+SUhMIuDer1Pho+IqL
pmbL7c9U3kiwa4XSPJIsprb5qTD/XfnXo2XD4Fhd+AUShNbCT3XGHnH/fwFymUK1mf+X8lBuMrbm
82UICrGkvqf1gtDDu9dh2zkGgLWptrWAK4Y9FTrqI41rOazuvpDIFJuRABtf+nhubTGhYpL53ja8
7jsZrmPvJXqSjwXKPR7gKDq9DFUIB6XIW2ND6rqSRvNM0oSr9pxNwNk9AlmQ1SOqteKtwfThLLd6
ALzQs1E1Q9x1HFpbu+FIpLQS4WVoNRlX561EEV/2jeD45gMU/gW5Q+cLpfkoF4qikM7T/eD+hjkm
urt0okXSj5GLwc+5GZ/9dOqM1bTYWgKSnfdDINQKAg8gqOKGwSay7/0qsHte9flDFKKTcvILmxwK
nqba+R/ANfgu1/6p+2/WzSzokVS2m3JAh1xijei0N/TjmainzneLOKm5d3M6t58a4AQVD/VkZQOy
gbeXMm5F8Tp/aKnwxqOj6pFh/BdPvKPu42cCmAImmyEKE35wolT2xdkyZJ1lNjrXnK1B4nL6eoYm
7/fwP30qFXKlnWy8nN9LUorVeWF0ASHenqdm4mqqhCOzC5up6q/RXGC9X840AxsBsDT7JtE2KJ5g
KwTzsgdmkd5mjIhPYlzWFoKqB0Iy7xN+ZEW4DJUmNaRUantESYS9Cp19CY9CjK7uS+syY27d06s2
RoXgbuOm7DGjCthMDXJSsdS9rWFBnsnxa8OKZVkGIWcACOzwrn+VXCFO/S7CxKUGHpLJfB7I086I
olifbfNdDrccl0RFgLQp5tylPQI7pd2SMcZZpAqNVLv7ZNrnqA7sTXSGLMGySIOU12Z9yn+MVPWi
xwla+cZ0AtV64HI03jlgLqJ2G3kmFslr+2twxx6tYzXLcrTPb1/JJ08+MDKn6X3Adp4PXErqx19v
BcAwni8uj3NqeUUVTyUnn8wJVHMQYdL6JDrjTqWV4SX+zm8v1hoJsxR+QTjFe2Mh5n4qrIEZbs4v
ylcrpdQAxov44Xu6kH3hzXD+0/TMA8aOi7cur/ZnMzcIYqNOaGqcpyrRQPLLrO19fdAAGPKjXaSu
aWScmMmnW+8JNsHSgvcTfxG2Fw2GeO2ETdtEQ1aF/QYQL0Jyc9AirXG0DIII5GsdudlUkvuvUNW1
30dyjHFAKBm0MIFrKETb1LFv+x/H7kxeONKNtAKerrr/lccgY8wlDIGEvHuTaDBHArPWye8K6Lpf
otT8JFCbV5LClrw+Yf/ul7b6xetWjslZKAnxEEn6pSp2W89pw/iCYY5TdwPfSFy6rgiwzzrf4qf+
UkR6pZwzoOYvIGa/e/Q20ZAKxWhCR3kbHa9b5MPsnpaZvSZYeTVfxPpPj+XCLIjwOvR4h5CLgWAy
k7V+UhoafURhb3C7Y/bKROo+AYjtuqk735SMckVLQggNycmmULe8FCdckO1xqsPo+jSSxr1gc/xl
lZ4kbrcJ0s0YgEfG3gdkd36HNg/aDGI7BRazWNgBAhS2RNdB5Nyyrvo3cvb0YPb0bBCOKOypPgOq
1yiDvAL/+w2c8GGl7FW/PBKS0ifKW2fZG3mcXxzKQK6NfCxF5AKs1e6cvxdsKAYaeOPEdfl6qeFD
6K3k+a1zFRpuaOX7f0gwhkNWdQgGbaX2XHYytCP2QZrSKMI3zjQ/GFZz+AAR5FUqDW/22bGb4qSi
CbG5EsaLJ8EpNMjn/PT/N17UUg48EmEzU6yIZWdSnJbw9nHZOxcrix9gki3sKCdeicKH8bfGhRoW
BRMnuEVIpbMcflkdaZ1hmo3+a5ph6cYm/HG6rI88cx/qCasq+7jd6+mvmVjlMRLJeBZLfx0JuCWC
RZ19jHc7G21YLjEW2j3MuoJ7zT9/UMTUbunOQ5541y62qH9pdhIsSBxQbshGqYyUWlnIieNJ2K2B
fU8Ab56g1fW+/Bfnmf1QcBZVU72s7i2JH9HuZueikB2u21w0bWrFoiPCkCIpwcbeNQFS92iJxiwY
NJLrSVQxeyLpa17JCBxlLRBPCVtCLFCG8X4U5lr0b24BrNNLlEYV0vOKMhuouRmd/FbcGckvg5ZH
13Rq9g+gOctnQ7ElvXECuOGJtjMF3e+QrA8nAMgRWbq5/wno4JKSD7/x10wp/MoE9X2Xky4juRfe
9mqKUvwLEuVinjltnd6iqTj1RRO7gj07/S0UQw0M+y+cGOSz2+anBQb7KdRRekHF9j7L3d9aEX2g
1wwiPmrzdmtmSe9cq+7QU59uewt4d4iZDIBstssveVOY2OLIz2NzQxfaSH1QeB/5GbuzAyGe7A4W
9biIFGkmK46EfPHBgS9v1lJvQ3QIKTVjDGzc4Tc0sQYTFRg/t8jjOOWs+vE9cWgxjdLyVG/WJOl5
mV78aoF8dOGJ8XanPtNuzxkBXv5oSH2B+4qg53fYYBvw49ENzjrgn+Giofq1sESxv8hGaBtooDVn
jSBsajAptHl9eH4cTgT0RO2nEFsixNIN/rth7SPvAHIhvA7KNFvwQJJm7GwiFDEK4nda59aXMYeU
diuOBZZnY8r7LEl+7y8aF+JsAtbaZcGzkl5k/rGxD/5aMyi/9K/NgOZ++yjWFbqM3g/cnKwqBYwH
XbuUysorDVGclfJLaHcRLv9szVs8PZNWqf0OhGbF2t7LrYy2X4etgoJvK71jjnMooDLmP16hY/j3
t089ifSZKNXs8hEYLge33TM+PC/AiEOZGNbE4qzTr3Ygv7+EoetCqp0ViXFb926Hu4LXn2IBv7TR
sj2nODSLScgeaRSDK9+U8XZ2xnv4qpYSCrHbDquZ0HS58TK3WycnzdrWk0nTVVuflJhn21T+ZygW
AbdarrFfQiS+6SyzxZXHUasiv9WJWRQY9xtzoWmlkHcFklToBNdzinKzlPdryGeR+Z7kyr0/3JNt
0dIk49x0hzX0NbLTmqwYpUabdjtzTx+IVOInH8Zb2sTJa+HdH6UqOw9h/LE9LhabDPkjdN4JRJbh
HmTsG0pz4gxrb/5IGHNp5dnuCoeH5yzs+66tDaciOGeiGTKyXhgFoAdm8TiNJTlsrqc/Y+zIt1Fy
xYp2A6c3d+m88s/bmjhz5hBQ1aqX73bfbcvN9WjWfBQx+Rghg9W8dCGpJilTmVRq0IRmDzy4C6cT
t8VpYqDZx1xSnb/EKJ7StSxfsJryY60TO6KWdK6hbdGxV58kYoMwwnLUOJluodqyvwgyndlOZA2W
VxYCzztioJr6/uRBdMQi2OYDecU1QmK9YzgZqg/ksOxfFZ54YBtN/MbUCLNnSRCNRj+kuW6Ete6I
QT+SRzzPx+GFlh54sfchAoe7uqPRfnxfRcDSMz9qif7MkDYR0t9nssiTBnR0CtMZMYKfPLKag78N
+8GM6eQ7ySPUcSq0Hw5HK5xp8toQak6qiwL7xwEycagYvVKkhfO8eB0wA5m+iiTxy6d2MH/W5roN
FOijfrpA5tP8IA6v12gQuVwCTZ+rC+Hh8ZvvBHkI6fki3MJhh+dgs3RrviRA/shTSC043dxjlhq1
GmVIHe0hRqKswOJSqM4pHO9s9GkRo3UUANhB0nv/KZcEGQeX9GUI7wnWDUDnjRv5OBHEOSRbVGi1
WllPfb3cArS+k/IiP3cpxpuSU0zcjEr66QaNI19AdhQJdRmRXzgiPMw8et+Wv7+2oXkI9AMFWspk
/QTr4RchpNkfM+G4ST2ODq9cnmvulckxzb4dS4rSzVKByObJZ8SCReMSdQ7V9ZXQg4jW/i5Hq9Dr
9iJoypuWgmxatoO8lpWRFz7laCzPr2YIwynkDtil5xZJk6v7mSSTPwhj+uPbb2YqCwP9LdAmPHGq
nu5ZgS2NYHKae7N7wj+e65SzhYe2EV/pI3xyFR9geoeJuHSaxu8sE5lEFFB53vCqZQb0pq3qOvHb
fE15LD4EW6Is5z2G2KogvpmdIYiBWyR/q5rn6p3ZLWwXk1pBsduh7Jt1g63Yj44PvwScwMDEziU7
K8UfjBqNRPbDvqmOkdQqtkR/c9HG5WqHKPu6lFYw6p/SLkcgKXdYS06RIcRIOAWYqbAFNBLB800T
xLsS2V2iaoCLWzP4tzrpOTFHq7TIGHHOVTG45UYQqE+a8gpP0oi7yR3mtH1QH7c4SuwmhBjjaw0N
dzo1MSGXx8y3oxJ8AIY9rX4BRWRA8Ws9fZwL6jUIxtm8r5EH7DkZhO5Cr46OMyjZ/P3UXoildxns
kpGHPhxHskXuj/+8mpGGXDMOQQXg4VG4EJg1Wqk8Et23ZEmIMpalukvoa6XGfE+XJOVqyFAcUthq
sSRcBSFqXd2cWMVk1+idMf0V80bDRKWom6H0me39uEnWAfEkK+GiSVIuCy6IKnuWYoHaZRCU633m
yEpJFhzxj/GsRyZs0YjLHkgJwDxZClf/91TVHvy4t5dy5W1IHksCckFysl0V0OXlhFy1DybgNy3u
TuaGwMaEypVREl9AZAucDmNDfIewT9xYZKkfENQiosVA83Sv1Vq/UrQ9kKtRlbNEb0XF+4PYcNaU
hcVT6eNS/jtwINaydwAjga/EnAJV4q6dP55sM8aJ9B8W+ttx/3AYjpm+aPAFLCSuqLVVSn2X/i6F
84LQZVPcu+xJs9+bL7+2SK2LhVSXcOKy7azjNyZOJN+JBnbjbxIEnsBFVhXFilPj9XQnVpzs0IZs
tz6ju+g5jdK6i73clAnDyAB9u300PNDB0R4VXbLLsZyNuqssspc5ClsBxa0vChTbs4x0r+b3i4Lh
pw/HbEPacX7Md8NtJgeGK5Cm9+rdDTAieoIq2zXpsnX/jV+eBifHAV0/SHpC5vYdlFdiWPuIy1W7
InaKlkmNlqhO9ufoWRPDq9NUvwFhTU4PN+tQo/PCZ3X4PuNbHACwW6Xf0qXCfwoNURS7D5nFluOu
9EZR62Nq52rC/OhZVWgA1Ijr5XHGqgNGTxoZnxmLwytNvopkth2M9ibV091HBrAc753RwZd+2WVG
4l6RsrJgSNFLIBfsnVq/JBsSOMmEmY5ODvsVNh5eafX0OLvSwL7sQvYRZtRpHDHZ5uMSO9tevuYy
SPJCAhchDh/mJjuwmPcivDYav+eScZLjaz/4iM2ZreBJj8e39PcmbcWh0qWV67Mh4HLNqhsJxyqk
aM7AfV+am+YPbPOWBgf/Owcp87HK7zbPNeDI0a2PVsPUya9S1HiXwTqypAaR6O6AFGdSAkoGsu/Y
BF+BM36hvVy7hqVvnd0+SveXBeNwhd2wqk6NBMZHDqwDYwqaHxZEuXIWRLF3FKbaauxCO5wTB/5X
8m2Y6QEp851KugkAIKFYG2/FFAt6v7uX317qJVem3meZ73Ed70oaqLFXHxzQujk7JT2e/DzwctCb
ykIDDi2kGLCByFyRULlKvTMZggvmiTlSgj4jj3KTc0UR0Y/axmcAwCh0ooIgPg0L4fD4/tTKSrPM
8euAUpDY8kHVRokVsCd19C7eT4e/l7gtUfBB0acNZfEhtuvWAePgGF7FBH221kBzPw+YkbqV5ASB
BlqQhpH2tsbDfYkr1TwLpxjuP4zXkvQYIwlId202wSxqP8FBrK7Yoc6pKjMUi8Qpz3ybe2y6dBZx
CEyiCVL3BfG9axYRTORuafe0VH7j7fnq7/Vd87BEoGfljCV/Dj7aftcDIGjlaWzDF/RpbRuzwz7e
juWPecsrL/1Nff3AYNWCxCjf0ygw1MwZFSva+jzjxG3XKFrAxFBABaCZGkxWtEh37Crs1AsuXILV
anQC4QPFknXdnMY2YZCen1Uw7jDXwxstlWUaIdoqIUiP1JhrGKC8emD7nPvQRzuyMiCdeUT4FFCp
/ZsOWv5inAjh1iDqI5TkAYlmNrHPjMfAm9oDjptGTL4IeOxBq27iIfWKorGuWqO5u5noD5S843+1
zN7KJwy+ZXygO+fgnLmgmsAs8oK15OsvGIOy00bz7iQcfF+SQmg7SbzqRA69tUfAKjNro2itprk2
d7z8gpAqMxKiz5ekDLe37yk7bwK046XFZFRbKXJt8BcI6RSpZqO0r5X1eLK8MQhmweFEATAyEsVf
6SdliF+17in/3gJGSm7+XCILSeQpvJayluzKR6vAyFBc3y9YqPZEaBXbc0Een8mdcAszWio/wcAc
tNhqOgD9uwHgcC/3CqF6W41M2PC6ylJJXhUQwL2ky5Eg77kx+xU0b9Crs9HOnOXUxtcJ3k5UgtQY
1Zeyfj/6SnVdiUEHDGkUgkKWs99+qatKmgiWnr+sxOK8NqK2KGYOcw4luLkT1XK7SzkZ4AlBbyNb
54D44G8oJiuHkQ+hMh2MSL3pqrfwsKOSKOj7TdzmtxbllHMlaozVvejOW7mPyACp0ItP651PrdOP
1NPeqDUDwkFtPo13XEZGNMevrKjvfycxneGgxX9CLiG+tu6VaeaNAFtAksJ5uWvsZJRUEHZ+lFsP
Hhej+QSIo2yHmXx/MVAcVzEOaMXG0EMGQSeEqNv37xna62jbgrfemFvZsyGHxJsMXb9SDHpsezjF
S1n3xFxAUzksCYo7MPMVA+sNhpDNEVcI4RqwDz7wRgMOQ91XfRgog3dvoEKe0wHHP7zzgy+0D3iA
87Owr1tDvRo00ScO0rnJqwpWVDcFmicnY/mvh1+rOeOFmIF9mua6ponv6Sp0ILJiRaB/Q2buQlHd
kQzn6hqs4y2ldjbuTGS9ApPB49817DBvAYxbvQ/1d7qIro3pNbOgHTUTWhdEiYjnOtSILaNhQoyy
YTBaML+IYsmKgmFO9mu1ReAiySiW5FzibtMci5tSgOQ1qn0UxzUwqeNvAjLK/TsFmbHI2ZfKwm3a
Wcg1JmjXKNWQGc8Vq6A03G8vza4UjFsophT8GtCBZ8SUU61RQXhEnMR2+uDTOehXzzw0qmIb6l49
fjtAVn09bxct300+9m071KzGnnVnb8stEEJ+vK6pHiwqNm4EifPyl/Zk4tpuZoHB7C5XxqtnJ+Pv
LS92SDV+p4zhOVodKvEYibCFe9p1+f0a5hJ2YktbjHt51YTnsjPk9cwIgxqSpGCLBO+8AY0GElo2
ZblqNzeYD5frivqEhd3DB9HLVZ8sBeMdX9L6NJYmLH357W3w8Bn3B9vIypiMZ3faNSIuhQ373+DT
SnJv50/XupbrDFiJVGa1NlIiz7RbPeW5+8Z+Efe0+AMejDbVdN02CbdcWmMy7JNyZMp7uuy5FMMm
0VFNpIXpxkLh+WBVLSVIf2MSbd92c/4R1ZyPbzX25o/fT/Os1nRa61fNsa2B/cn56w41Mh4zNN3p
E8lEMlhqrklK4Hkmqqki1rNHhgB/T6tx0Gy+qcQnRP/FfovSwFUcDr29T+upmf+bXJTSpvgiDaD5
v24MpdrYnZeWAfBKdKxbuBSCjYPUmYdCVmo8JtK0YhdJUkBoKYtopapqPq6ExSRYzyz4QM6bhMNm
atVpvziqby6K6a05r6acvM/7KyiDfYaJfXLKQFX9aATHAgqdSn30I35pawF7kiAWL/3rWMj8EvMg
64uzXykFebUn19sWFvagKtzgKNXGqRO5MyT93JxjoueoJKhhDIdxN8wekfQpirt60VRcBJ4SEEzs
3xOHq77YffcW8o4WTWDBYQW046Dy6uxuabILWMxUwLmbNIpsCPSs8dRuUO65m32mJTJmGSkzqZ4C
Vs38QpNlxlT/MzyppKbj0oW0f47IyUYEtR2lA4Tum1EXoAW/xcvacnG/1yGl57HrNGaxYQPnvpfM
+yThp/pCFxTRIzP2NPOBoz2KL5bQOLZOI6hjrDdwMjEFYU2cj48rSwT+nIDzizUscQUldHWJ/jRX
oed8+UdppUiUkeuuKbcVfmhP0udLVpj16CXrVEycne4oKp4I2jmw+mM83L4MYxssIzFsYOxznXE7
9MdfiA/19Aa34///oK3Fro1C1SNv92pw1BosLxEf4IQndmj2v/pYLHJ+9h+C4T3Lss0FgR3enHFT
VBvVJTLlJVDNUl4cC4GN8koqaKv7tzr0weln4FnajNl26FMBtcIRyQ2AvQZJmjM2Qilq9GEboKP9
nfmtmaH3mljlo/YSAEoRsL4bB+xK/XyGb8wmbeR1LIYcaofIKphHUmBwzFTHsSxyyt+bO9zDA5aO
xl/1rzTScNQCQiIE9/ObDXgDYz4VHFK4yLnS/krLQUIhUQ2Ajl0PkabgLoCSb47R60cdmyqJd/rk
BrqAkMKnWNiG8m8u3u9kmzUgo2p95yghoKljIht4yJmspJgDiwcKl8awHR3jB7TWHK6cWQ6SLV5U
yq3rJ+cHku/RHLyUF7kICF//d4j3H192IN2oM1g84XHPoBFmPxs4RQuLPE4033OBbeKLwnFawt1T
x0qqrbd5ypOgZUGIazFCyIc5SG3Iop//cG4pEJD0P4Xyk1gyAuOyv1TzIhwAZKo6NNhbeFpwdw5t
XUz0DEzfThi01CDVAWP6tbz1EK2kGaGZDWWjFC6MUxuppyilEYP1awaakXxoLB+VZePuwXeMEv+s
xJA7pF5a+FRDiywYVdJR0FUpNmi4ACcfyFV/U7Xp5HwQ7qs/Afuui+K6dCPKENAK5RKG3dyLfaBm
pitM8l2RTer3XFfnwi/hoUbTFKbAQK0JC//0Y0lGyI+d6b//Jyu3NAkFp8bKvr2BjEbvF//Zt1ic
cZBu6KrqwrjnCrAu1TP6B0hHaCm+55f/CId2/7OyrOj59cPJjpnMu1O9zeBEIcHrSt4ZYyeRS91x
Ms9y1Fz9SjfB4USPkRJia90grQ2GeFfQ3Vsu3o/92Pt+Ic7v+ABcyk9IGro65Pnh7RIerMU8lyIa
C2qLAE9ggxYB9IYrHjUOed08LcSZU/9rMcdvQn+6grzr8MgzegST7F0f5rw6RcadZLFakX+lv6Uj
xMr2Q09HHR1SYOkAGA5xvD8AXb5va+erH4Z8CbO0iQtaKaEZuhaAuPYPGHo4LlLmNN5a2qIG/7cN
0MiTWTQNF7wFPNgHZ7OSXhJfTuqZzCFgteUwWktLo1cWe+Drpb8TUm/HH2POoEnWtyYUFMqzTQio
W457AvQ3OhXGzbKFRbvDIE5QGgp8X1c4wNzdG/e9ZUHCMDbR1hy4bxIS0RPbO3NFVbGK5+QjSSw8
1RbcPOeLt9Qd0YVhpfKe3gMqFarHgIVLS+RvxggYPMPYlW8XCylsflruiv3FYKHA70jeNrGXyGVk
YlqrL3cgcMpI+PIf3FuMusjqgC7KKzGvMnC4QPYa7eiJdLNLYPp/KSRvCUsDVIvaPX96XBKunWSy
Ym8RDvKqs7McgEztREQPbMVQH+D89YKiebZ2WxFNLtjju8Kpo0C9fgNEGzNnuIlfnhm6xIdO9cjM
G9Auuu4MPdwZBRLIak6Z8F3De6lTLDP/7dy3SI+vw868rxAgN/gGRJni4wCF3wkfTyNA6zY35Mmt
uznF/eP78B73AsPKzq+4M/VOLuSFnCm11IuJg7z62zxVvQXLdK28kvGdR1MQx/KYVWiMZAPPOpyg
5JGPagjAriRX35+YDIv867pQKZ7okmY0UiBIE52d8SqFnssbmDNDf8fcx5Lp/XB4Od/NffoSGnsx
euZSQ4hFQ5z/BGZhw1WZhQ0jFqvIcowojJpEXadcl32sQPTMdAfHN5j6UttEFD/k7stcvlUDGpY6
ZjnRai7uMUfoB5GZ69HHJPb05AnkxgIp2Sb9XCCHMseaerWVFRz1PMDIEW/eZQgB5rPd1H5FJzxp
fCtnQl+MmymLCaPpNRyjdDLtrJ1KsMG/1apxd1hOHJORlbWlVfGcr37FaB4O/zhw4rWap7JNZrTM
kgZrmjfE6hpZ29ZCYZbld1rf4N21cJZSYBlQB9WVN7x24chr7kLIbqC8YlHlJ6Atrw/sCppGIib+
TGJji39KvydTqZem8LrJWuVfHkTAGfPUnVVMtpjtE4Q71FamNiY2yJT2in4ae4lZHw2F1bNaM1ve
nj90CYVJ84NN2HW6luQeI0nfLaCT6V4ejoNprOSAGcETPOU9UNL0f9C0Gl/jG+Atf0nEgzmlHxZT
I5iheQl9jxRgGG2aTAnRxf40Wt9/vTL23Y6YhjImFQ3f5KghC/ku4v7eGSD8c1Iy3nsrck+mBmTW
42kWHQiQPd6i4RYxV36upbraaBoStBD0a/Xdq684z+gKtHXAnYCpc5doLZVdwU/PqVF7dqg9nBcT
/UWEZKvvbPZcQx8aAVmAprMoSSPzpBJquxD3gBbXYYvG3dvhJjUkSyLutnXGWUcUKGSOxsrKN8F1
rrSC3jTEEL6huol9Py+ptrtlIXKgTkDyOLZ3lZ6SN+RNeZgbySd8zyOipEOCD6BjWTUyWEs6f8Ee
gcd/Dwc4R3YXHA0Ozzeu/gplkznSaurIWGVKjmYLf53Vgy7pXDOG99aCKRkJ1kbG4jHc2dHEAfhW
/+kydTgR1GT9lgvo5WWTjlNuXoRXRWdJVhUD+/ibTbZEQGCA3wobhG4zSK6QUEzxbBBs5JBuL9kY
iweS9JJBZKDCGOrGsqktZdTu4UHxieh+eKDmkwpBm59wCfOdlKp1oPEYgi8f5KIikR7SzcKxgvzb
GopyXamuFnKEuVaB4qBH7rco1IdSUVWOz/hLPhCsZP9Y9yJ8lom072q6zmWaJF+fAJyPzNtr3VUa
2uRXAUSSWEJgFp7wjo9i007e/y659zeoALX4E35w3tSSIiWkUFfXtw835Lyg8MR79rZk3T3TN34c
jmqs8mfxOt3qHERJwDuJ+T3Cz14hlqRdYlToQQYtASxQZkCDlnQhGDL5fKJhwNG3cm14xMd2C8/a
roUZvc+5lqUxsQOeSaB+hHAFuFeSMOX9hG+3fCJ/VsNUBUCToSJcBNo+RAufNd/Jxdjq5AVhi7MD
47P5U+NwUL+fVzdFOAb/0xodi6A0Z2y7YcDAdgX2lX3ILVyMxADOCWPZ0OVEgTS4HtQhyDfQR5R9
8zMuFcOQejnvZxw2fhaSisQcbM9Z5Ovwb/ah8rMacs8s9OpISeKl7IODVaBtL50gedwc9lV5weyl
VZL4dOCwwxFtapnmMh4ypTRRIuHJbBMIowwQc/LcWruauGDRnW093W9E98TuKv2Pf9ev56809Hma
CvF6hAng4HJ85fZ5jhIuG0EhVECN6wCENYj9Ds94w6yuLfMhoFbkinL4KRC5/PUiwfilzRR1Y/fg
e3usW2hZevsT57EYcW0reOm0mSD5zrurI1bf1H3umvVuPTza8pAslwZI1hYHYU7RGJiYqjJr6RUv
YFREE0MdwQhjgRvsqV05SZkF7ref67Z4RU8ukPQWf+g8M2Qzb2o8PsWuHVqPVxTLVIV+f7RnfMcg
JYgwBfcge1dnut+lcWskpKrKpKk0zS/3zDvbnrG7AIy7a7IZ8hpucqX2lXtj7YWR+dSXMApYo9vc
5DSn07kNoZ14iZIpFWC9bwm0A/KIolbE5K9qRSEqWi3fgGAap46e/NQ7YIPzn6MccNOD7trisbDd
UYZWZoeZJCbUfRog+mdBVXSlqjfrlYWIw7KdR2ZUgcISYisUldU7RjUEwHtTt8GSzaOTo4EI+xji
xaICXeIYWPSU3Q/sGvvV7sANP5XAhtKFGFQoyJhS64fPRPatvbDFu1WRxsogpeMIpFH3NWC/amcU
e1JkUGGKrgdI7SdC10DzRoqCHuLMolBJ9XTOzgcJKmpW3VQph0n8FpcYj/Lu2BhCrz6XJtUaGRT+
VEzzGQB6zalg5Y2jS5AbmKhYInGCZUepLZMGK+rYKPZcBM5V9+AJ2WUMS2oec6arHs1hTxhbXxfL
OBp2l/yTXQse1sEy65JYM3REQIv9XZZ2JIaJJlqGoQecdkrULifNDauDDcyH1CzxG48nmUIAc56G
EVb34a3OjmvfjxLKNqU9YYiCzSwf+twaB1WNP3TzrDbCFn4Ua7JVEj1/EARrVrFPfiIyGSZj2WBg
zskhzenH0vKgHa2pVBIKmsQC/o7PoIdvJYs6T800w45GJK7+5PZ5n5rgkmK8+M/I62tJ71KYnkW9
szqRG9cPSreyEttKw87FY4bSRFMj0kMT1iql+z4BRRfvjWVe9fLXNQiK7Z0xaNWXV2x8ZPrK6KBB
xnUHRgsqQzVYXs2zuQB2OWEumNt7qN+AA0mjmIMH7r5RUfGA1vSsfWw0nAtEQulPaI0PNxwlg9SK
+Likkb9GoWdWJUsqhLfJ1MJBLpMQnf0K3ZUw79sCC/5K4WCtooiUFeFkNXXWHQ11rHN3KYdjql+g
Y/JhxxCK/2kzIEU7U4EBJlL9XWkHis6iMNGlLNCrmCBo3C090Z+zSMPIlwCVjKgfebAiJ2eV+wqH
Dl21fOLorcxYhzu8K0KCsmuSBmwXkdHWLnYmbxdd+2X1Dou1z8iOxIdzt/cb1aSY4/cXYdSM2BIi
kfEYOAG8nXoUDZXCO4lQCpOV7scEP0bcTYj+D9iV2jIhTDMI4H0ATggPaH2+81n+34ZujFZdXAwE
ClKdtOa+lMyJ2xB3kpwh88Pyke6s9Z1aORJMToQoZ0VGEjS+i0oAwpigxySY0dE93pXGqlb0GKsr
09OZvSWxSVtO+6uTm3KSakLJWN0SoBk2q+ZO5UAVVbzdz8hdeJqCZazT5JUouD8OyKRN6zqkpzVn
24tXBuPHEDOLJNXn6HvRr4W7WeErGSPGjmC7X0BM5Tz2r3CUSXGZWElsjenZLEAaHdk1LPMJTbFV
ss176NPo9fHA4f0szzkPzEvKQkakhqUO6ytvSvOaBdl3GAf4AH5EPDUvvhdLSSapHJrr+FsW+FwI
Slv1Zb20eVUAnXP3bVdTASkvloaTl9Q6N+aht3r2FXtQYI1FS/HGME0ZD+J1nQ2a929zMhE6bSwy
DTelD26AbbUKbQ9NVKZgI3eNOojnUDGFbQeW0VmenIFhHUMMPosT2JH/MFemdJdodUK4hFc0F0Ew
tQ9ba182YBq+0UdmQ0qiHWfdrWQolRvQ63Dme//v3CbbYefJpVjjcqormjLh59djqdoou5d+Lgta
7/WPa7Yia94bYNGg7N8/IDGPDVuH4Mg5se81cLgF9bbrt164+vfEXERbcU390fhBZKExIwxOBTl8
OJt3ILkAdShpKv4GC27z+aNpeZwLN3mV1UovHSXTgskQsdA1kGIQsQKG+FCRKfF9E0aCbda2HkFD
CBP1zNh829qck9p98UJshee8d+6dH01KLDiSZ33cgo2p+FHDOqkzHG/0BORy3V9EEni93DXpSLif
ryIHYQq9lUAaLBQSm6JmsFYBTgqT2mfRvW2iRDN3CKZD058LaK9tolqldfI5r1fGzIWCYeEpTD8y
Ks0iWprKqW0c74TaWHqcLzasC7cFLpRDbA3n7DL8C2vABJt+HKCS86DSxSYqzpR+jBvEig6P3sCF
TEdHK3E9093WEeXKOMbp72FOARmc3NmGvfMBpUGR9HC1XFWcSzAfMs2ubY70qGZTGrAKr/XQdv56
GkZRMHZ0BgxSq1VETF/bVYkr71I+wJ9wNUnrp80ec726CFWx2NyiQR4zEjqD4N5M7GTqk770icgL
mDk2Y2+S8L9HuKqMJncM5gCe3EKEV4cnTR0khjVEXhMNH760rExBW/GQjvOqZm1blLpNJTyOq2xP
Zt44/accL579yd2Udw0wramr2ZRCJ7gmepeh9zxtoLQD568GCeJ2cG5QK7GkGgHygqYMg5piv+Or
m6sshv21BhkgH3SYCYjtKfdYrhBwnxV+g7PthTMm5URuxY5bLniKjqgmblHkz6QHkYtZQo6ieYUw
hrdeWSVgzIw1h6q4vKan5M8neRgHJ0Y6qHhM5kTZd9KPSf8062g/h43V3/bY5uZoktHETovQrkvw
4j+J6WywMynL/z3+uMSjveG0fPRgshyTK87nL5g0Kt+rjsXt9ZuxnemCf4ZCbEgmwlXYPoy5XFq1
XnxXmmYop6Avk/OuWGXwvvTlFsUn02OgtMqtl6es2PdVOga+q/LUfqDxn+zdYm58hGEmr+dwcAIr
UIaDDt3qozDOeGQ+dBaAUTQf8kK/8fKzsmL3QJypmhFq35OpYQlD6pXVOmnHIXrySaqHwT8cl0Hl
bNTy80ZzaTS/GjWS9xZfXGPYu6DHexd2tYX7Y0VNCweV7aWRKoiFy3rlANYUZ4S31Jv41sZiTxuj
XkOdQI30ET+z+5A60wJHjc3StBbf6aOsl76hmc1h/Am5DugM1weUvnlUN/oPRoHzwyQx0GT9zvI7
VuT9CMp7+TaXu1UPw1+rqNhRK6hP+wrHMubS8eqgZ3ZrZtOMOOVUKy/yoV69hhUGPDf14Ie3zcwW
uGJUXfR06H0/i6VcLwVqNHOX2geMBSAb9kamA9DlKc0XAdYKFw5Qfy4jUkA7idyUsUqArtpoh4aG
KnPr9hdvx9AueCSm3ZTEpsYLTKwbi1SxpJRrXwPMwq0dDsmLLHMcqs2vLa3puCTOOu0H8LLLx3PN
jO9aGOmxxsBSeL5o1vV2MVEqyN6jv6hbHbcL+Uoqj6ZfPgG6by7H0axccrrxf/bx5I4HlFXOU3hV
0zKDRYWMrykWIJqsPouuS2vnc1KOsy1ATWiu7xCfox4wML8EZlXe7+p7dmlcOv82iQbLOxXX4jSt
7YHjaPqrHYFSLI7T6UnMbgVY5GawN6slIFLtmDpSa3OPsyWxqi2tK57cddqu46V63PO7TXLaSXq/
AoOYbNmme12abWCj9rbQuXBLhFnxmD4WEKExwGIa0zZDnxMGKJI6Rb6c/EmIP3nCSml9+j+gdKin
cjBUVsmzPDuKRzHtMbvQO4FKKkPiK9+K1EEfOyqqnLIoZ0p8tf7VHgrrBtGDmX9z7xnsaBgFvCms
0+4neXwmyzQ43Yqf39HFmiReH+9yRTH+Cd3y6o9J00Zrz1Y+tVpayj1aOyI35gnYe1WS+HiwCXkw
XE6xcb7Gyt8JzQr6Bo7gV3jjLPpYklw4DwGcCRORDjoxfKzIkjrTGo9w3rIDFFSpT6u718ubWztA
zDynahP2MA5oleJoFEcVb6Se9zzTMfNXnhZz7TMMfygt0tihLq1IRzXye61cGuo+eYh9uMesX4tY
izKx5v5noVrhAA1ytuMFLOXRJ9pS6VWZQU1dV3IIjiTmwZFPv5O47ySjcXoNmE74XleqAjWRJVV+
6DQey6uO3a1K/WMFwKx3AfBWIlyj+AOyHNOJUXjyJYbH0NAGzEZ7rDJREk6MXOqYHyBLGXm3TDl/
S1IgRiaspN7t08iPM+Gh8/22j6Nm3DfKP1hoHDWx4qro/otzJVcjBwPFfVohL2EFp8mdFOujRWf7
ygjcoxa3o7V2D/ap8PwPKtm21Brh0PBClCRvOfBAEEieT9EjFRYxa2UJOV3pptE/Xcfzvt3ifJrg
Dpd/RQV7XlMgI7VxsB3eggJRsr6srqMCrC3r20ioAGjUNLkrX9mP6kHh+bmu7mM4pxw2LhhLyLWc
Pf7vBkZtd8R397dFMEy4+7VSgPXLUfqr43bivQ1BS2OPCK6/3rR17C1XlVRrQQ2UJXRjDFH/5v6b
2RkjQ+yJiPXOMvq/7FDPy4tVzVPLSvYdQSpDN/qyhiphRc5teUNoOhm7BaM0pYF+jK+F5uOG4oBE
fHOw47Sfqc8JWtzllVi8AHjVosf+qixCBYMu0k0vptJ834R75Veswrqnc4MiBb7xOnEMsjPdAu51
CyqeDqKS3ASYai+9W2Ya7k8hLGFBJrFM/Apr9IwBzt81fUSzmwrreNACrS4v4pDfYkZQ1/9HgOmj
eg90YSTplY3aKkRmTzqnaxrDrWANoVxWImis4F5sxOxrjMrfYCZAB/4bypG+7E/2l5ZRLW/TvxlO
TIpjzR7BC1XM2TCdoofz9ixLLYIhtTxjb0A0GeBHy9Ai/38g1jx8cb8pLU6WB+cZ0U+0o14WuLFm
RRWR7wEQArPEjlbm7Y4QNX/2Mjel8JTYxXgWLIeYRE7Y2uCHW2svV4uXuxUbVsxZDqsz6UGQkBzH
P6lV6XSVdc/NTEPbO9JDA708Cr/oiLzkkbD4eSaKL4XnUs9NSfwMeoPzpG8skWcU1oprrfU3A6U4
GF2v9PHpy/zfD+5JW1eHOgxBkhWfkxhy/W8e1h/G5LPYW2XY5fBL67HwZCRsZOJf6F5//SS/91+g
DCE4nlNWnvciwJRINiywCAdIP+Yu1Y+5BvOMfOCgE/QVGlusXDO089IyJsXTBebzSKmLBCd69fkr
KP3VtOLtEdRRojGuKDd1DKFa9FQIDkgy+jAcCZ+LmfXrVuby72waNSuUXq2Q4AGPW1gkQqmDTKeU
pO2tuAgVsyVR6suSRkTGYSfJ8pDITYI2HhPPmTOsjidEmNKsU1EHf8mOpjmpe+iuiB0HSLuHgtv6
dcsZ6dOunke291v04ffMz4bFkxISwi1rTP067PC1De8n2S4wVyqgUIUipamfiWa1pDT7Q5J5B0Jj
fFFV4458eZZIrPRxoxmwQxsVrgqK31yq84L2uVb96/WTq16Bj4RHq8U9kNw9JfCbGOpApdT0TSGH
5Wg6I6HbjtK6hkHiNhTYfkohwtQbRdXldOE9L5e/7PDM2pHvagaCHM77TNImSSocdNzHLRUp7x1M
YoCHAAC8LEdIQpuhj52JV5LDcHXqsiyYwEyrJzyXSsf3hXZVoSfpoHCS9UGuSjgaIppL1s6cBh4P
MWwRcYScFW1UHkpAXDrQy/XFybr3LxQIW2iMI1ByJR6937YUy+8UqCdZ5EWbetLWIunsqa+92bCn
XyUh0M9GXBoZz0rjx9t88RqxTsoUySK2mA4g9xLSsyrilommycaL8ZPKrNUmmEm6aEEX5WJTU0H9
IeeZOfjZUZpRgBCmxxBoqQ4aV0cd8R5r4DpMEG4RUd2ayQ639EfgYJ3tj9v7H6Wet9sBKiKYATyA
dO1TFVivF/IVO5TUdo/holhnSeqJG4s3JCsMgnWSnvu59LhzmvXGdGnQuR15Ybpm3t6knpRnJ8Om
6l0azfOqQhHAIO7OGNjSMCLKmaiq6FYtx2VSPKwGqHMyYKglGxCFSaRsai6K/lr93WXhqWOWZFBb
RWB5cJUSvOuXtqUJ/GKViZTQy/4Qq3HpGc8SILPknMFX+Eo2eREoJgwf/4Yl76whNzKVzsai6N6F
YRVF+/mp7SPtLkWdvW+JQTw9rTiIznx3lPMmazzw/gK5E4o1v1ew2zQNccmbC3187NbY0WpHSmaA
XvlpxPEmLOZWsfjtCId6PqetpPMjUzDTTClzvTcDnHj+dKYKqazzEro7d2i3DVEte/vSvjRmehFN
6eBwHnOyyUSjJso0YFMR71DkYCkh2vco8ShVyn3FpfxesC1xZZbPbbkPsfaop2cGx8sjSfm9bg8l
41m+vdkm64xqeLBRuHjlsOb96/4tkZo3VgYPeuymtk3Py/9nnBrYfdhhWtosNJFW/p8w52YV3Gb+
FkG9ktFzCESHJbA71thoY0uDvldlCGKGt0qELayOXyBssMX1Ynz9pKkfJ60tLpfsvuCosweFfhhN
dZhIZd0Ecdpi7CcTMendGoFvO4DguzIz2bzursy0mwZ6HuhD9hwppSDwCWyYKzsbac46PHE6j6Dw
7grZ9wcly9uFv6Rpy/5DDkcypaGxh5aRnrvNDD1yvAPCMxxrKcES+v2wPfsKEr7RwPA0/XjgilLN
/NscNR1EwwxHJwJIUh5DOg4fFaoKP1JuqKi/lzzYEJ+87j9BDpjLmTSoDjeI92UYHxXJFgBdivRU
753lCXQCW5KSGJH9zrtXlpuAz6jwtFQadRTSUgAtuaRcF/HtYOJ2gXbrdvZ2YxzHrmU60e9Z0hH8
CFAXvcgcBaq/bnO7IzF47g9Yv2IhtvGevYiP85/BJcJx2xSudqoZbv+QsAVAUZb9+wZtMRNCt9lQ
zlDODdiGGjtbjhIMdJ5SEfDTYJm1HW5orjFhuQad5grlB5mYbOr8hheDExCzblG6RpZrE00aQGBW
OMkk5a6z4Zs6huf5+iBjikk9igP7RjpNFzZm5WvjxCw6EcUQyx2QUujuH9Z6uou17wG9ep/jQ7WD
S62CXlVV2CzE7lxsW0etuYttQGbkzKaaj+NYjHRHoTvCbReWe+ux+BjYEaev/ZT0GIoCgsY4n6uF
99Ksb6WHVEIFKdoTOp3IVXxbc3EtCN8jHVf2UeHb1Py++LtA51HDZNZh6GjjhQ1GHpuXG2NlXxYK
8YYhQjGeGnsoRoCT42miGBmU4TsK20yUqBDJPmzbyLVEeuDQiF3HFnZBCgAJZtI4xgnkF8ExbWtB
8YQuMtK1wD/kBPRRH7yVYBxDoM5E41ssBW4m59SnQkvrMLcXnz54CqDpR9qV/29aRPkoBGbcUHkC
QBxd8y6C6Jlhdk89eC4VI1mr5ffvkbdQssqHm8BQZlj9pMI9j9FNX06tGrgwDFUhTFgn4OSwlFoH
nwSZ98893t0Y7iKNEjcMdAmJSjqfQhnUj0YKKRzCtw69ahlopLd0TbTWW6xQKGyzQVwcNq57vXLt
wrLJ/K61QK7pMOJB9WLgF8KKFvkAng2+6Ln+WWAvEdgGkCdcR9fVaEdo/d5kgthV8bVUZbBnZNet
/rpJvZ1+9TmyEDLNG1BLfnPPIHhR0b5k2feMQe/dv6+sSleH4pvvJjLnjwBuz9hVu0FN/uzUT2xi
nJuHv18ydrx1fOtWPscFvwq/xMsCdaSLGNfgmLwRd/whllK1h7BzWBjLoDM9mHlt0KfhRBaCupa4
TsLI6TBHM/I5KqGIZ76a3+xluxNy7ZLhhwnZy3PPlJPfX+yGD6hWgshwI/z4i7fVk8ezlNWC9O5c
i52lMZ5VIlV9q1AnfzNxoRnHGPuR6vRx3bST4sSnOJB7O8dOBOhmZuoEmOQPC6bWB5DS5A015u4r
ICQjoBO8EcDnnBn98EwPbDzWZ3mLk9P+siFZocce4nci9DfECQYZ0I9QnoIwHENeEuw6RwMr7jKT
x+drd60ROLXOFcfOdfSFb0dgGlj6eBZZX2IbwUQK5vQBgU4M8YfqAep9vY4Ae8i6XgUt3KvNItjD
kmLS0A0FJvA2T4X4oXA9igobQprLzziXdBau/iRBUxDl0ICu+p6SxLB5XBpiieifTtPdkLiuO0oj
wRhRlRd9usGqwSCBnpPQYMg8IBLi+3lxCFs5FVECMddhHlqX5EPnYM5ClGBLxanIJH2ZG5sPttKI
XLTrhx15piMeTaXmLLP0U/836VECXQoF7xk3EZqma7/7s9EApOKjaHF4OwnXdl1lQ8EXSefWjHiP
ytdMN3voOpAlQV1Eo9JGsrN/KaBd9iknwZluk2dz5HMSXxWIeHtAO6lKNawwh5yXk+h7GrrdZbc7
L991ZO6VonwGSdfe8pFPERhoF2dCM3HSfJAPTaF4/th5TMZo1ClXG3GvSFGQQ4iKmqO0NhWYvq9y
iCQOSdQt2QDm9brqOp0GBCikr3C/ktPE4bnqRqGc2Nrqt/4btjuMLPx2Nu+IfA1ibwUTF249dvfu
/8/5z3bTda1ISdmVBxPDL+LAV1XYwq28BDQXzR45MRm9gilXW3bVr+J32RhSr/9TT3rcAareKe2g
bu3kUzr+4W2Wfu4/CYH/PFuEVUQOqF12Ksz7jKTJawYQO3YfBqWi+YnarCH3WAd/Q2gKS1j4ZBYV
PUmurZs+foT8ErblobNp/cCH9WDTX2xoLaq11AnaMv4xFHG5hkMnRhhzJq2jaUFacT2f8YHfzCUE
Zx/6YpjWTkaoHO95HItd7biiLUPv4GJYiLmQAyumOoN48caOVbbCKY/Ymp5Qklui79zv1sJOXHRp
bN3i6dC0KLENnTGfvhEdvZC5u/yV7FqKOAHu+/Rm8Gd2/QewcV1UChPmuL6K8UN4Hzg2LXIdIu49
kD2/YWMrEib7h3qwqVkO5MXBv6ljOnVdJ6PX+94LHxO5TpqWAPiIxTnsxOYq/iPvjryCADkq81ip
XwmwfuWiZ12DKhjJ3xMq1eU9kZvIQsoESjdmz5C5xyfwW22W55mLHvigrMR0S7B/vYYC2asRBFJw
E65K2qthnYgM9r8hasFLHnsbowBuHXY3lIpUYTH/LF5w0bI/aSON2duEWXXT6mRglE3OiS2yAC1Z
mcKV6/IWML1h19KJ37TJveNNMcI39JqGhbLzi1PsIfU2VtyVBlUMe+7VTvcOInH96in+WdpxAiZH
adesMOMGlsoFrukwH8aFJ2rZ9QlEFqbPux75INn+ICuNYpTBlZcvhdTc3gpNmYHAUiclHhvr1wtA
4ecOMlSpgZ3ArBDmFop8qKejEX1pwvF64HJW3skeNxubyLaOsrvW3k7LyfRdSbk4twIXVt4wqIjr
oboETdBrULzU5K51OIgDbfI1dMDa+rQzVC3ZKjWOq4pekicenNV1QnejPo2xu4OcpgB1qhbhNm8P
vBVILddPeuuoX3NKtl5Z/Pbn5Dp8yWa/dxQCYqK4/cSvV9Erihx++taYAX8xWjoWZNJ5/F0Ru9pD
BgNd7FggIkZ5cj80wsNMsu8W+WWczxcrsQquROSB5BK2FoxxAVhzuNMq716RdtJ0UEF27uMa/YHb
v62GWEAuy6xcg+eAB5ZfObrGx/KdgONKznZ61TDafmGHDlIUAtIv3QJeDnE8ia5ig/brzR84s7UW
mX4+gy9NRqDLgcUShnBbBGx8tNKRmMtAef737MEfJL/VBgsEa6L1T4v4vT2LbUN9PHeJ4J1oUH3d
9pTpxati8kyG3LlVkbWyfU+imzCMEL/0zZUz6y4GgWV8OmO9EcoeUzZcFutWo2K/pGZpp52Zm+Zw
PJd+iMj/yml73eMLMgTbYpzhOBMsaZlyHR90jyGyZUk4Fqrlx1+1qvVg0rzeTNhmODNRcdCXp5L6
DE1XXpEOFrRcycSkSSYl+AmNFiGhsp33y6xS4xmLAKoLY1uxFsT5Fmc6WwQjQwUohFYa7mpY9FVW
TR0jkqVqJTJoXAC3sp31qVnf4HM0QVqqUhhec94PssnA0nXI5B5ZN7LWNCwIH2H3j2/iqw5cBHj5
zON4qosJ4x64h2VmHcIgdFc19jlv5DvVcESw/pV9GvEyQNsFQqLX/eRdL9PwvLASild8AR3YFTtP
62lZB3jddhNSBii0SyX42LpRtxvWkJNL2mA0bbmEUXEycxMZPYWHUX00/gVTU1mrLMivKUevIQ28
J1pm+lWGfBMmUfT2nB0Tkd+BrI3bWzHDMfqTWnZo7T2nK7pbNJA7iOsfkvawYRkHEZaA978UwB9z
BzQmt7oqG5draAbqVUEGvFxoCpyzytbC+16SaK04ZSsF3ZjxMWEVX/eb2wyeqIFBuiQTfeZ4mYj1
BdJr6NYbrE9M8xguGSVtP2PAreNKqpiHxSITf/K5DcyzsXITYKMNrED1KIdrlnEnAPltsKfa0v+r
zLCU2mhuW5a8SnkZFFScMLhXcIbAmYamv9ZV7cTmdnuZE9tCC8RpCBce2QRYXwoAUZbq09/dfqIB
GzkE1oFrAbRi4GYXjZi3Ld/f8GmLM/IfFO/JPDDemOkVHEgSfhkzC6QIQiNImLIJ2TBZRrSXK9lI
uaujpZiQJUbkp2heGLxfPHRw+n1H41D7Rf652Zr8ZEAx3qQJiEZAltF6Gja1kXIckbjJhXH7kWdl
2TdziFuh6VLqZPsd29rNQHtwxJDvLKAecVTSPwzUAtyBTdhzmlvERWE5RJZiP3YymprFf/qEV7cl
zGs/m0aSh5SK73jrmbqey62Pus3BQQwu9bN4kKpF/PVwabdTGpVmrVdbvR5YimLxReV19elNSzxH
Tvo0q+4pLm8q0my9IHYahwUMojsZiVKQCcIptZcS452JdIYZyZROUZEWXPv6ropCITeVdWLwrmpP
yFMO9fVe1YCiqNvNgu2W+r/m2tcVgeTQNJbOvDUFmkDjv6E4iL7KQ98iRmMjY972U0wxFj2is/fy
XaLmDdfNPrWq1ZmnZzUfyZBsdkeSdY+98PfLygLpaQe5GE9CDtsTHb36AX6RH/XPyzBLGcg9MtbB
x7kvR9UDC7+HHDMIHrPvUffNhRXJywh+TiIRgvKhTzLBX1Yz7/5QRA/TXz7KjGmT3dFu90Q3+uEe
3FQyiyXTt4psu5a8vTRyzonsDcKhTJUcVSWw6TmSQxM9J71Rc/cOpn9DUEJLJ2kLaiLGLHXTiOlj
VntybnCjk08GNhzlPTseULf/8p9IKUb0WAHnnNx/5xlAopLLdKaXjt/9CtH9lx3IgSxXhLYmAPQw
nbJaTU/1QSvbxuIeBwBbZywfddsaXoW9oFl+3LyDDD8V8Gt0qiarqopmsevJAWxVHOGmH8LBiA0C
kU99nxa70soXhdYsPZ8T5COllaCusUAskVS9v6aswS7hAqJQqLz+40KIpszvrtE31EALr90CWwY5
5o9XBix62y0XZWO3fXlD7Mnaz+taVxSFPMbAO0WzDoowSIU8zLNZ3R37N/lLjmQXuk4cSk56p1+v
Lxr24ZB+Ur7DOTD36fkm7VVPL1jCy//g/MJmTqkEJgtH3gROL2Hkt/3gQhPWceoF+SeppwfR5XFH
yym2hJZPiXtYgB5g0YFfNDj5jVoMimticjPPVstYnBXg4ceMUZGvSODzN7zI28obKQqqGy1yeiU4
WYiK9fbSQ7/8KJIw6OtxcyWm/25PnFJ27mK7m5U3chToOZYx4hzkg/xGeLblwOhvIf25yG2TQeOt
MLdrBLL0r18ac+ReWdOVvPvI/PFpD/DRHtCDcX+18U9hiV9KLt+pZCvTRKavSvVmHNeVw7CLyFLY
YJSwql3XInWzNqPN7hgUT1ZsVsv/sapm9gHXuQEjpBhkgEUJw4e9GVWAtYljCwh2N3U6IwZM1AHP
khlou+VBhQwXTEIiuJP1mpoHU3uVmB83zX2xpH2wHCt8cV+GXk9tAXjh7erdInJpW1nQBaRJ5Xl4
Kf6SYHNepFWaX+CXGe1uhNPKqbRopWXU5RTTAKqLt5Jq4aCE7xMnz+YcEwloPZJ4GV1B3bdmh4Nq
WGwqShDQYjtazzoichLMKNGO9soOvcdxiKkAirR/Oy6r8NuTyL+XPvne+Y8kdLxLlLmWUHWgLm0k
XuEW7EVvEonm/2SJDm62H+/kjEOiXT25FRVoH1/xUNsZI9JxMXej4idsQKULbJnHkkD3z/oL0WYf
4bPrYpjKSGOXB4/9haBqntpR7PsOkolPb+DGElrBlbwWmITn1ADqCiOgODwgdHgl1kZOg7O8AgcH
vP4JsxvhJUc2bbe5Csvixsczj4GtNhNwszI4Rdak4b+0SRgIMMfnHxzoKxGi+6i2k/niCL8h97jn
tF3+jMrp9GpAxvpISTSXIa/QGu9tSsh+mX8smcbKNCwrLdzmsWAcp9++LOSQ0IfejnkFdZBdbJcM
7mbPuQK6ZIJZaNIPrgvRcgBCWEh99MqWfOIAupLUTMyOrSJrU+NhSU1yfKPcU8afkLqU5uoYCE+n
7mjDP9hsVj2NWQp7ezZKH85V1IRaz7Sewbxqbo1swT0N5R44D0QO7tl0B9+GKydC7shZvg/AplR5
HbZK1OVnJ4UzWW9HOF0ELdgY2h1vqSKs+Ft6vQ7x2ztIbqeTMOmsFe/m4VCceh9JwA1wvY3CPbb4
xoOr1DKDdfz2c9vP1JoMZMq1YaPhNjXgqIhOHc9metiEYVa+1uX2KsblSLL8neLV5/UiRJmMHCp1
3nkTu1l/C5TaUVviDWlh45w+GfpVmBaTuwXU1ORMv2rUjpwP5EauVTr2iaW3oFn3fY2g3zI0lgNx
weyCX0FrDzt/J5FxovZeR8Gf0+wyFUSIs4bF6MI2/i+SsAXVPU9SAgnl3QKo+bzd9UYnS2Zsodbe
XemFx5Zv1wLoe/93moN+RClADyDHhTQdjBIUc85wrcByCv/xpvGyJi8Nn6tApxSZOPApL+hF/vJ+
IU/9iByok8OtD1XcMHnzcD/XlO/IzgePU49SHsOsJf+44ak/DPeU8p/mnEYUv9rxUq/L9aqHL3TN
qxhMZWuE2zwQPhIjMR8etIsznStmv5xiC51B+ywR/Aw2j3sEW5NZrb/L2OTAIoBVH/brUR1p/oHQ
Ygq57Grom9R49GAwTYyyvDB6e27cd1zrs2c9xCGFVaO6Iu8YOO5pIDkhbWO+xcaQxZraKMRxFGx8
FGkhrmi7pB05bKTd3dJFPoz34NM6xgY5Kfb5XjyIGb6Q+Yidm0OEh1wJPSSPOsFRzKQICMi5QB6j
UeYkJobg1QmWf9llU9mv2HUQlNYftJuza6lj2ta3zgjpkoxf8UmR9OBEz9dTdnMWp1sq4Itx3EZ9
nP/lYQJhB9z76KV1IeYIqbZXvfG7bAfwk2IdBNQ6KZtQLYJdGQl/W9eIIRiVqm2nT/6+j9xYAROM
sltp/igMsnFV/p6lAOcYGLv63CgQFUP0+Nn/noN6oDx4hMWdGmIRnOIbCZQEcCo/qnFUeEabH50N
QFnLmBjKHfyn1tnghevtDg6+IwNYa3aC5vtkjKdTQhonGxnQ52WCpJnbxH3CmaK2hIxtaSXx/ad9
CrTduyDBK5JD2NmxSoPsYMloj5R3laOcqUIIWR6EsEFzLNrDIFCaa3RV0d18fg0thFI0SBSgGlJG
nqCGYTC6mJAfoOmwwhRy+eTSbH7YNQhA5Cyi+1uMumPV43DkgH2tevBfGmbX4DQjQa8iKBZWAEwP
LE3oFR+A5m1ssxXP5ujbKLuea/OJ29VikDH0c48eB5A073R2Sa59/6OS4f823433JsVeoJ/o8XBg
Sdvmz/4D6GG9IyBDGsibj7VxJ3xfBx53CmQt3DqAUc+5S2DXMPx2Fyv3oG+lnKKXcs9guRDISumN
ZO44U6ciIJA/vYT2cuoKaeoh+fopCYwaoacq7kIYH2260j/ltEW1iLWAYYyiDGR7HcStcqZwcb0P
0V2JGWKpdOI9wdvoeFtJqvDDHwPuGiZx8hmEQ1dvxXG8AGWpDlkH4bh5l5zPa/kmTABkeBozOftx
o0GIqqglsb75wccavCP3eTJCpnCIL/1Mu47FRqaYC3EnVrwscwSuCNGT4QdzRHfmE7fnMyE1Q/2j
X2tXLuLN73+1lgZI2LZXF00QSLujIuh6QRGp00v9/SAm8+vQ/rqwJS6VTEWMGpsYj1nGPoYH8U9Y
fATwIOVGJGV50rxrlbnKdZKmlfLGshic8DwR4lo4Lk6k+6rLw3b2b4TgncDkSe/iBA+lNvrr9/Lq
XZKOQZp5azFzzg1r9B5PLEej2FV876//Qm0n0c7agq8L8oo5y65r9SB0svX1sWYz/tbZZmLbXFcw
/OIjbeGc9gNf8rwhBLF+qfSDggqC3ZxN/l1fg+RBSqwwajvaeAIWT7ucUizgZ+6wjWOSHSkAj9fw
DQsb58XKmJm3b+NHwBD4V8i66b5q8nl8zqaClQFEBw5+lUHyiYkgyFdgkJEh+xULnAbR+GLjcvAf
pa2WluFEgO285yV+pQU7BkhdWw5ggFyUwPYD/NRncU47wSHTAECL52D9XzVMetiNteKpkZDwCZ+A
VDVOLpbFxJKlrG81icmPkY9PkLjjNwLHMIb/yB8k4AJucR55lnPoUGyZpw56iW+49pcvXxBsTS14
k5ZNaerIbCNFQHH4UCme+hMo7emWEqeM3t5MoQu8AIaycDl5oPhXx9ZZebXQaFuryg16S9WMdv7p
cNMsltDNRUPTkuuP8BYETC3wkKjCcBodsp+drWoZpfE0/pMuj8Eyn+EtVQ+xo9AXHPIkkd7jqGKP
35bQ1smahJnAXMh3OsX6lnbbCw8KN8nFYRilKT5kwobvgXyC18KOLGoOX8j7yKTcAFWeg1Z090V9
7c0IyDakS1zo9LWFY7a/KeY+USFXu1N8NAtuM0ZDAZMYkzZkG1avLDYSTz/+iKWhUlCn+kCHGqPQ
RHr6aMv0V6XW0hfR9WoQyujNGtJ88qkBW2riEmO7Nq5SeOvNfK69UApyhAnL8gaoKKy4VCrM9sne
e1kdxxJz5R6KWORWARylcAwFEnr5Ee5RmvmoaG+ph9Fmw9jO9nxPGH4jk9TNjKsxoFu5zjD89sNQ
1/ZaFcpSMhgRNJoTFGSrz4tr6nPBo7+6vE65N5rqKtJwC8QycqxAtWNoDV4ryCtWeVhODlc88aOs
kkRCXONw5IUgWEsdPDRR7GewzsFKBt1OrQzOYQCCLTMz9QVaLiUadFnVc6Ni/5nVG28aAciu4C6O
cY5lTnqghO59mDNbi2cMHgarKO9fkEDMNRJFs+Bq3+HVlgn/UWfOAWZIDqnbZywkOYJlRnIW1Stm
vfT/eJ+Fh97Bi9kdCguA2+QjmSv4yt2hZnlaom8h9A9Ifp9h54Pfj8nuA6cyWZfOMvEEGXn0bt8a
Ia/zNc8gzIZxKiJUzwBf/Z/SLafdzDOUlCj+NZVldByRL96PWNiqGWq0ySzyfL+RsSeY8D3JoVEs
fYkmMwPNmSsxqEPZhxsm4wHwH4357S8Y1XPMGhxfSQQbjOo/Wsx06wLV/JJWH98pdqMV+EdqqSXR
CpYwnhtaHMmG3Y2OvhpVlqO7CcTqJUcrC6dWwl6120n8RLQ3uoW6zTg2eo8J6RQCb5fnTkyM8LCA
aUeF49y4x9Ckdk0dA89FcvpX4JFFy26Ksn5lInGJnEN+0cJD7onpURvMNbdWPI6tOrnaYDgFCMAr
DQ2dE4FsdnMqCvr7RQPtGj1ifGQ1O4N/5FUp7uHSqW/IeOr9wsJuNvKgOAaLUgIDwwkKe8mVbgr/
d2XsmW2OfJl2y+Pidtop7uE9c3AsZU0f/bN2d/zVjhp7uoMRElIuplGpkd37wTP+WG3gFeigBpov
rjvm3qxyFUce/RxJS2l/H24p8U/6II0nN+P26eYrSGlPSQ+kjEvB6Ceq5qD88T6DV+ccGHrYomKn
KqzkM7U8ws/P+nL9F2GNUt5VvoJPt0qb4YwOfjuUjGO/sE2dzhn99yZBc1a0TcfS8b/CndlpirUW
PsuO5xu3YdBzPcOy9k3LonLvHInZA7MFthnMM74+qx5lOvyrZnWJ277SLfLhoNAhaJtnDhkhXFYJ
A6FlR3v+6oYj3fpJMPI2EZVqQxMuCQxigeDwGHUKEgeIjnoAxYUPL6XTA3llPMsj9tyhU/zHcc7t
up8LG2W0IO4AjQA1BwuPx0a3KZgbrWbiU4ExB2cs+gSNC/vCSZmWVuSG3XKp3XY/jmvVoy03Wl5M
GObf7FUBeY/Yhh6WBFzIhZibFh2mifRDPPUnaSamWL+h536Ih2gTU5W+WxSqH0dT3bvEOYkCacHa
NJJrZpaOYJ16OYFpvwEI9os2JWEOpWOmdFBRw99wkIMiBr5HB3i7GwBhfvK0IAdtyOBR6zjFn74o
52p3WkRHcLGqWeIgONkJh5+yw7H6maqbrZiiAxwRKxBopnX9Xfr7W8cvdzz1tCxbluxhsAo2OlBx
kFLcV/h9vPjTPHZGBkysLWS3Ax4QWSsqZ40tzrNvcZG8OPA5jWj2SWb9pcKA6ijwtlcQ8/EnvNwm
hkGZyZJBxI+mrtKpwt/rAKhqO37WAGpZlFr/l3otJ3FEGi1aoN2tAKHEhI8UGvd5R+k7pVqRGKx4
4nr3R+G6VwoG+0eHk2/A/luewWqhnoN717HKvSZiNdVEYzyZ/x3id/kzmWthMuucDW44BdXDOzhf
1YW7FjxfnkpxUcrW5GLp1QuGwBBIB6/XD+1stZnFgrUSsoCqzoFr5IAMuxumOgTeIyvIPAM0yFXZ
5Qg3w93gpTUqvrtRWZIucpaalgDVcPoFtmJbgaIV6MnnsHzCBfHyOT4b7dWUxDq5KC7KiPzKWPy2
2/smzz7N/vItLSW8bnzDfrqHkqk8r2BOCQ9mz7IkokUx/ZQYRDw9jD2wj2aGDZTK3JmVVKfSfBiz
J9izVgXo1bYgtmLYEfmqUbQcubxtpX0xS+l/M3rHKTtUYYpO1HlBprLqvZjMemixPqtb+qM7uZ3m
jOZ4o+BovgOZpnHbdX6aT9MCarAV8920Lld5oXDAslDGSwA1EpSgPTQ1pY1Y8iz8jM1qgLn3i47V
0hnv1gij9NqLiTIA6U5K/UGGoET6hS2da6sxixRIflByypurIqUmDvWy0soxY5mZV08jXVVjTh0e
HY/1Ke03yRc+CFZu/g7PXFUxI2pgGUm4hRIjv+CLzf/4Bu2Ezf1xDDqTMC9dx+kIPezrY2NUtnAq
7DohkBKAG/fIU5Df7f7AA5fYh+OAO1b9oycYzZQfqMX8ghKJAnYztcCjNSJG4Dmr0THhcL5J7uUN
2nw8pwVGErGctRWgegMUBxg9AsDHs6i6sXme2gcpXL430X0pMmIybPhB/6naK0bcH3PLCmHBocQP
BWfBHBX9cUU88RH/Wp7Jc3e+1t3RrxPa5NjiowepQMV/ccs87DCWYtZkXgvW8MVYKfJe5cep8/1C
ywEacz3M2LqPLoNhpWjUL2Bzbf+5vutoJifrQrpV78XX74pMxN0jFlJJnRlHFwdpxb8NYWeuZP/g
+BD0GF1GjZOo7U+UCwh1MTs8AjNqBIMxEru6WyCEqSH8kb80TG9cn5Uf/GlohLNaZleGyFXWlKo/
Pw1o/WynnaG30WUmdjUgkOTx7VJMpw6Ux+X+SASNOUASrtHLLAIqDVAu0X+cDVq4g7oFJQCatJwq
cN4UlD0Xnq7gNz5mB6MDvIEAhArXA0DnAs25nzYfel8OCUIPlUOjtci6ZkG5fomWssdrGlq67IrS
o9GXcz9XtyU+Dqm7/e9OPHL1dbqIYg5raH7AE6yh20CPVnTLH/TrscWf1AeteFegDLZRsLo06uWG
VNlKkXAmiBvOhY4FCZ1axelGjHXWAzwZ/aOaE+DuIMYN9xDYlhNZ7T/gBoMJpSIR34fJhtRO2VAt
JDZf46ij4zWuj2St9jDXbieKq9kTar2tnmPHINKpwlO7bH534FznlCLuHOv85+I/Fr3y2l4yWBL4
KzSKa49DJhWxtUiR3bvg8H7WpizH3zDYsvWK05psF2gBYuivKdt9cDdDdVaw1DQuYys4BQvh2XHs
9koX24Eqz+xONwC2qiDSffYWCrga/HZ2VQd9m4SLanbYiZXwyCLdPjD4feRScsAE0LUIIH46KTKm
PY70lN0BnCtDQcKdgdzxB+3/+ZOUXv6obP95tNjwuXcjQ+O4Fy6lCsP7N8oUgAXjxN95NFBDbWoM
WAnwCpNjkBKCXOKMDyRIzpayLqf+rxZcnqbhWNYJaGQvOAK5nOvgENmRRpJFU5K9ypHGDN9OWfpK
BZgu50fxjP8HkWsZpSyIqefvm186yrq672rcoAU36/E3n9r+fELMkTH2tSdItjAt+WoPp5QVvNTc
6b5wx/7I8sI9rKX7DmXrvOJW4a6ww7shOfU0/GuDU2mEF76WZLOweojzs6IpTZh/aZUppUOZFiTX
YqrvTz+bGoB1/aV/v9c2FYGeEHfTD1BvzUGW1zBWrVPxCpRhGnnomlS1CAhDJ2NOEVuEkieRxWT9
MgBpd+rLq7vQHh7Zw/E9fykkP9EFGxSlHQsR6vWZYopWychLlrXLrqj/YwY15k7iwxfAqMVIacCK
eONcYyICHe2q7lUu2B25QlTnKRWZWl8R8ZqRZ0aTq7ml4biMPK6lV0a741qj1Dnnsza0Q1OWOpxN
F1cTiUy9bhZonnO4smIpZwSZY7gAejbDyUQd8Mo3A4Nk57sTWu1RptC2XXBQlKTVrk3tlDP5WOa9
55dvett4qvOAo8UhKler5cmcbRPdvrpSxRUfrpBNNK/ST92gyFFFriGej7QQxdQz1UAgbhnsY6ig
lB3EhTSMzozRG2lr5nOj9Y+5qW+gbK4EeaHmdEw1aBMfUI5gZ5KhCF1+HCnHzPglnmeEGHsDVYMm
ROfoPPbOhaCLmMsHzTGOxSEyM9tyB5mpEH5JkNYdQm3YqZFLMi8kgR9ls9b31BZOEffzuv13dOLs
ZppZBeY04b4ZDplRQ8r7NpOOeFKmzj+t3aragNVDuK4V/eb1RgknEj3Sj1K6dJ4yPQovw/NWAeRt
sO2dAjTZlyCaXuCkdl9SI1G9Se5hauY9s8/It70daC+Ce+lYnDfh10Hi+rUlx2k8l6MJhG4LULuV
J5wMyCCeaqoJOhlLXHjsxCJm4l4idym+EM1skKDMPQexE84YAuuP1BshgZB2LWwgdQg2ate9q3oc
mu2FPDbJbjOnu5Sac/bzZsKg/ooLhy2kOZbjq6Z97SoBLECTHnTeOzjEWRI4zjs/c5I8/k2TopgF
KVMo5TAU5cGsn2LAQyjKrCR47FrCOQIn363/S/9Cv29UxVRJcDqHX/iSlbqsjOYRFGSIYKD4W3zl
sY4e90JzelLb7aKK+x1gefbXAvWU9zueQcr/L1PsUipH9yXKgK/pthXYmma/lEruSTGEx8lSdyt/
Ak1nkk7UYFDHyOBzGhaBHvRi5BKxBVR1foM/d0dJ50KFc3bM0r9ueuWtiR+yF5m/VmrhgFLG/qM6
gljDLgVcTFP7F+Qu8obbStNx9AwHRscqSq1GLIs60+GKpetPmbmsuKbrxzLuOlqDWAqplyhRe05w
AiPX9A5OanprL+tX7Uv6/0WAwevQdG+NJCKYe5ANMITjrrpQ9XfXOhiL5ep/SBNl0H2hmHXpzN57
spy+qkH0ZzssVlvLKuxiW3nN51IKD76QmmeNwnG/T1YpPmhdnj/FeFIBSBz5/iPJMhrcRf1kI1sT
7GD5fMN6KsIMIrnZkOh9Ov3pGjyozZVFhODbUBSs9ILDfYL/YDJi4WCrWLUd6ONtNGhAcZ0bdqBm
m0NgkDSvJfFRelUNYqJBwHH1nh5juv3ZWDmbGgKMisUR5tvQXZXBrwhLrLn77NMLesj+jgeonzG4
FhoNpgaZ/k8DuseZk35+VdQkL+8QckbCrOaktWk2XRJp+A4J2OyNhPS6A1LSBf0HN2caCueKSUq3
ib3BdGwrlsEJBDStIa1S0TPMAMeE8XPJz7WZg23ll8Hs2b/xb4LE+VWGgZzPW6xHxb99N90IPm81
BovXktM5iQ0dM7PHt8oBj1jBfzK/5hwl9BDDVm6ylbqmt2S5j0mEmeke0tTfjDyOZ4YXwE4UGlLm
htc6/7Be8y5VgRgNfWXLivlYMUtJt4KlbFabCM+qCwQd/qKzso1nqSfdbMHmwc19+1wTOcNmwtXt
ODRUVKsoP5MSxyoyw0/1q9o29diUlfbzBODe3/8IgGHX6xSp7A2AopGj3B3eEjHRZbdO/t9U3nq3
xOlAhYNiN75J65YWsFiUdyEfVA4jU4mRggDFvPgQnt7PdEUuv0bE8ci+339FUoE/bLdMYgPmV8BT
bz4G/nAIYGJSUS9pxXHmDrZuMPOqcBr3NZpfzuZxOcJvtDfb8nbvEtt9e+uymD9+ZyILLqIECLXY
uT3KzXPzDxxf6SbP8qzsZgLCPiretbZlVeIBPeMIprj2OlvC0U1IYwxcGD7SEsCeXQURT6cGW3m6
I+8RKs77VMD7gJiFvqkMbHFAo4fNUHBMoQyeEK8RcobUmh8r6+BL/oS2bEkFX0OQr+rvhxbQs+h+
wJIfnJTX3sG2+qL3dyBYE/RHfGk5nm67ggAGL7bpXVapdUa9Aygttc+UeBvTOMbUWdb3niLlbFFU
MUGZ92HgVu5KZ6+LI29Zi4MJG9UeqRounwzXDyJIIEPvTVVKbMljL7nh+HpUrGMaZCuKv3wRl8MB
phux2ocCRIu4DezXkPasA2PrUUs1qEKBbSFLO0W4OuHRoL1iz3FI5KKQa8rPtHuJAr1uh98RMeWA
FKa7llYGfS6VzbR5taBpIKmDL9BgXLSSb3IUdOO363BYpypPtgwAUghihLT3lKKZjKJbfI/lIPln
ix1ULC/nHGR8w4zPBPvl7XuV9XLXox2xwO/MOG4E6w6OfkkcH0OmAKlsYx7clEHk5sIvWwySUmZm
XOGa/ZUu2FdMHiuCXfk7XcK2BYGMoHhOyftUmfo0OaquVDWm1im0A9aovczJDSABRfFn3XhfrA5M
bgG4wrsAriupYdSpKD4xBxRwiwLfY9iBO2xonqHoi7RlAHsWlhe6sx0l3BFac/RcvIPTcMibKlhG
FFrsRyLgndGBbuT8QFCeYx7Tmg+tS+wBkoGmLB3ELM171QUH2aa8eIPAT9dcWdqp3YV/M80UyLIy
V01A8W28y/5wgCooKCPYiNjxJGwSiMpe7sPBHsikyrxaf7Ixo1bXQt/J08zBC99vwa5vHnOZ+BHY
z8WdZrXSlgyzcaBkn6k2Pc692eGMBtiNSvs6gu5utimTFVpBaBHbwzwQuSlq5FmTsxgtFmxBhHBv
CB/cyoou7RhXtcRmJ7EjzhRpWv7UHKexXnAskQJkZqIyY4WWs98iiMGquEOof4yC2ocHJSzvLuJp
P0iWig4E/iLjMLOKw5RUPUy3XuQoNihmVT1ygaBv4cUHu/FFyxs/QX908oXTnEBkAqJ1oRTDu7t8
AmvoSZVdv6Q97raTLarpWAsNigR0+1lt6tJQufqAZSiKMlz6fnoREUL7naLxNv8Buep9FWx44oE9
o80faqfzu+m0xd2d10DwerTAw+8U+LmIe7YDFb9SjueqHqI4Zdho+7IIob2176rV2s0rwLQyXG6P
7SIq54WH31KrdQhKzaZ+X8BEyBot5FFE1rYtN6qfzXKSv/bIS+pWmVtO1yDPsb0Q+SnO2RS8MyI8
UpvXK+blCbOMMiZ+dcWk+DtFFvRXatMC3DcEdX11EKIgKe5KqIYLhOcNKPrYfZZ9+z6355ViaNQN
d5exSNNEN0B8rbmzWv8q4jaYjWClQttjW5i/byR+OJ+ou8goIHnUw2hIsCQkc0dK30MARcndwva2
kPg9byZZMyhZnW+olcokOWUMcCsHqNAFu8Dx3FGikJf7edL7MBmFaWt4Borw9KLz07JwjQH5D9Q8
pff6zakluKBDdEUReQNnFRdKXvtPjj3NkQ9aKps4zncXuWGwxrUm+rdQp2c2GgQQ0OiDp+Kn3Dit
SmAATmBH6wGTv45W/TDXI7bd9YuJU8QR0yiv/mO7qSILEvnUcbojwIaDOuIDoaTXfCJlWXkutKLS
v2TFlhlv3lRVIMnPetHjJ1/957jzmaDdEIR2CUJVvkGL2YZVMqpCWijzKqMSgDXfd0Js6EyA9e1V
QPxFduh7cIF15ZmXVjayS2gBqEtBSTun7PqDeemOzWkhEPUuCITDk9lWdDGfC24gDTr1dpmFM0xq
RcxLLkHmF0foikjOGBaY+eGczynbPcQEK8zsA0t3Py3/t/7FfbsYZ17OCFKPplUw/iJeSc53iqLG
bXhKoejfD4OiyUziH6wllbmeJZznGxHhOneCUYxiJUBPsEB9ODUWw3TSDZVr7tGc+NYMFGefct8/
BChEEokiOo8iXWrZx4QZLG0aIESCRYiuBEDFrmGmTPUbEfd3jnwyUso/HqIBIVHtMH4tBnhYFFFl
hPohXpOk2Q8u5BI7sBgQzn2oeYilKoCdCP04DydDsGVoXVBGt5Fz8MhehR0nMEhNoGm3HS+hy5ri
dBA6eZGDWLWCjuWXjmZkw7YhwgLctiQMeHJoJDbnqHQ4qf+7FLRp4T/9RUgTIbTFG65nP+DEBFYF
xTvQidVBBwrGiUiu90bTNAWiJiinl5T+4CKiIw5+aUWowrQNlwOuyC4ZrxPU/VBr/bppVHtV59O+
tQLoDYB1GxUX51P2CmCN3A/J/GU/IwtkkhB7z9vXZ8XrvfPdMl3xTck2nfqw7FKhMjtEggHXzscS
eNHM7Wsh82wtByNfR8D1QGedDz8GAxkIxsDrexH2J0ElN/CID6+hQvln9YMr9KLgyXU1mRPC4OgM
2F0e5kl8qFrgSr2zfs8Ef68wpzVB++7HBIQGSmhAMEUlxnIrhPl8c9Qz3CziJRdinYUQvO/nZWrc
NVJVgdFgtu+xlTKedHWderTj8CztJL282z3wDSpc2rXBJ+hdrUhKMvlqcfEElBBTNeypTVfQwsZh
4JgrrzvXd31AWuH20SvrgCp7IYKEJ08PwDDqJtmJqVoaSvep7N52fVm90XgdiIK0VjPhEVLucMuy
1lD6LSKcAJloiG/Zhbe4XcEkqKBc2MW1f90mxkdK4ZhSfun1WrPPAaK2enpFZiffURaHaZ1jZEe8
fwOA0ounVA73p4+uYwKAcEejFbigmEIzozI8L3Yu0c0WSwkSGitrOjN/5qipF5meRImzSeFH6UR6
hr15Mh6leug2XIkUh/NygncHbPitkSpH/mpdVpKze1UsBcxVxdfO0By67cVuTaK4NPUtnzhhQFRp
KR5xBuBMZfaNI7IvvGXQrwupZMZh48T61uFhzaVTNH/mNi4rYH+oC6SHEZkMEd5BXOGFS4wodsd3
deq5cvqOa9PYTTb8nIs6n8K2l2+h1Xifbg3OOvFMzHyMsMSS2DpsyukOVAnC8I+gRwl4i//HW7xL
oOP1bd5z/3MFBAuchGqLK+3WyoUcjxHaKlKSj/tztgeu4l8KUxUNJavlH5ojeTHCavzVOs1E66L5
G4IepxkT++9q0j+O+ZhFa1V6Mog+rmHmUiSHlnPLHPKcjcTs2CUX8tQiMTcJf62KRDtl5Ean0m//
XE0iirmc6I9l9go0EAN4LML+XvfLjRaJTHNIdi8mfYw8GqHG6VvB/BE5RVSTs3HKiWIArjhCd95t
JmrtO6FzbeS6yH4IXKSo0FEBgH9pC6+s8Nw2PjX3lraYXFkpztIVLokgyQBB5ykPQNIzImAkVTJd
q5Vy8XCpMTDJoZ2oVNwHQ24ZymLqZMCY7tGxZUoI7lkjNjoF4N2Vg7vP3C1mykXJlTfRG0GlPfvN
cxXfNYQvLSgr0N9MEYPR+gD7B8SuiOLiGsdyus+cH1yEYGUAYim4nT9b/TiTS0mBPJYcovS6iDsB
/jTbxLTS9jA+rcdesETwmiZvREPfwGD6SdIIfr28LgsO08NNYowFevNiA551kMTOatL51wP5eUfR
K1z1V1CKZI9bN0sHljjUr1JfNomI/cmJEh+FM8VPKnL8oL0pnR3USxgy8L86DiHAzhWULpEBYcng
pLMZfyZSxq3mC1jE6lkRMrfpdmgEEp5OS7J3BQNS7SqeJwxp5Kww5uNd6ERvgUGPUX3xTkmoI1a8
cYTswKSUqG1fQ5rDvVl0TAlHdhmvoYj2E3SRzDKg6qMZhQzkYz84nzwsJCzII0Gzw1Jqc1hs1AdL
2cf2pbz0BB53umqenYiCA8gL5CZbuCYv99BCOln46c45/YBOijpCM2F3Fi/+UkJNndgza5BckjrB
Z/BeP9Fgtsqr7I/hKhB+oRw6PF0mte5sCT5tCiGdJ5Jp6UqI1qn21lrs4Q8SQPSnoW4Q8dydu3Aw
AbcuabJr+F/FWpt5KfTGg8Gv3cY0TJa9fMmJuIE9Ko7MOmQ17O5u+xmdrB2YlBy/ID6A1Ql+l2jT
cHU+hWIhHWqsKgxGEFhXHCtcfh6SMOBFbV/HYyGI2GyfzeVJ6k+osFHxE0hTgaGY8R3zgVyp/X9J
nNNIwYTcM820soHG26fgdM4TLwUts3aDtqiwxlYxPn8trOkS3FMxNYZFAglWlf764xEiF1jtfT1H
tm4xEtq0ceS70BcLxO268m7AXJuduXHlZlwYS2Lb1iNFpxv+H9f4UPe7xGlum7bUMLzKEh69LKG5
ta8nlKSBKmmGSrHKsbhYtisSnFgS37ruULC8FAjYDIMMRLghAUwBzxdrJxEV/JFisITVggGNmcYZ
2vmqz4yRJDA7XbJCiSsOHVpcZzONdTEzut7x84y1jdNf7uUHKTy1NOUylq+2RlCMf4Aoujz9w/7m
ixRlThwSONjalpv7oxB7qcv7X9MFG7a1sCPOYDXd1/sle8UAgTQn3e8XabR3H4vnBjO8BJ8Ai/SX
taVZxo+4e9KT+jzikZNeXE0LGnyxjwcwX/ZllsZ0LCyrP1dvMkgB8mDp3UuBeoTiE1jFv0/Fra9Y
/CI+KONAfIpADARJukXAeu7gbt258eu3+uF9ukgE9Zj7bf7Yi0RTgh5SRfEhpSf2KPjcmDYfKqXi
U6/Y4i+QJLRv46KGY4TVGctdr1jepjeix+1aWfvjEyqLdNzVNHYLuOf/ZljluGFg2PCA8Juxw9JU
wls0y2sGEkZcnJ+Ea3oryj4WYFbcEhz0pk3Vi3t4V2ZOXXkHo+64K7Ym97zg94uHq8+aR1JkvSVF
BMVvoU+oOpxMyEPV2l1KQTaIvcJTi8WrdRHF6hSxp2Tcpg3YYMQ8heITBEmG42SJZTBIwP5iP1qG
2peArsWJ/+2761DEvuKpT5/QL110xXCghvURtYqbDZuONDzOou2Q91BWXepjsz7DK59z7fJzs0yf
WPgK4k6PwEWJD9TT4Lkt1gveoeITDKvu950IUlAydvrTfbBMAG7VZTS2EvRmXrNoc0bUucleEHTA
t2/JR2ZFs/uDGPe7N8G/922dFA1vnLomnrmNGbkvsWIzA7KH12WpzNdB630qGN0qVDkyY281CAGr
kc4+UIA6elDy+EB+dI6sG4DlukQA6ildRb6S9jhtJD13idpFNPD6lHqVMZHmo4GowETWGBLxTf6t
Cs8C180tlH6/de9WaZJs0fXwhIReDieSJghGLTb61GVnN1HAq3S/SxS+vyuXwBqb3WVIfkwakP8P
9EKbWoCW51VG/taFfy/8ta/dSmHU+TNNpJ4HBXX3tYLiqbJC6+7Pa107dtJWr6wk6ISBNkXqOlwq
1wulEC613q1/+WaKJrEXkfzcNjTxl5zPcagVM5O+TL5IDDUihAhwLyYQBT+2CQinSna9YbzMq6HX
EQvIwYQc50/tKwomoa+B1DXAnC8uZl1FFz8LRHPqjJoAbTQVplwGt8YspY1ereXKJDEtJ+xg7NJ1
t1dJZTHbOVKYCKnL9nb21LhVzKSdYkgfKLxub0wC9VD708oNsbzP5Czg/8mBee9hgoIiS9CfZdm9
7T6MPsvvuB+RRI2qhoOiNxKURcOfqR8q9N+Eh10KcTUTDh+JzfXkcbcScREeJUqwEheFm2L2DLiy
Z9ZE9XXIy19p6dKFBcd3Ql9WXWrAf72aq/wup/EYi1+J+G+7BnLOQ7cnMPjcaMtLWTU7kKiBy5If
W6QvbmkAQk4YTlJIwWQm25EhQxCg6viMxtSi57nLogIIEDPb2oGhHPgBkizC0HaB4AteUtE/i6l2
tv/6BWAMCYxEBXdoxqwHb0M8LDa2Wi2RPk7+mOmdh3+zT4xLlHHZ46bVf64AA+H9NF8cY+xEpk3x
foVGSvES0cRrmgyLLTikEMHoTZ5Fq9tzLyucIqUcgOn6ZB+G3VgC+NStEqmu1SlJ8ckbqSqZhNX3
0gCEKtG9o5CX/KLycuXrtmesOsNEZoFOYCxAhgmvfBxwGs1rjInstWUrajWXvtXPERppVBO/ydJM
SFLfXHKts8R06sI6FFHWttAPp+I40Wtz2BCIV1OlMktwn34Ge9iJeQU/lUpa2UUzkoobXUGWxSma
XdIyisNLbp/YpPaIR3AU8uyx+CRnCZbHOOFZ1xk1L2QHi7xC5jd3DNj8bWVsKtPi6b5uUpC7e1U3
ZOtaRfEiqKoPLAp3nwvwDiR7iQ5hxnRyFY6Ysr/w2VIOH+91hIPLXC6uYzieJ76dD8CnLA4pcdAQ
cyj9u4STYJ+wqFbDYIdXgrfZPhgPX1v4tkSDRnPe9A1lsdp8LJ39yKQRIVlln/Hrk1mcQylPy0aQ
bx43fzWCZ3jlCJm5atbtUhJLxkjLGOWQitpk0ppMQ8BA/shaoBeN0+QbIWb/lEtDH6oMHNB0eK+3
WlvLJvCzb4DTMm2HzqgqHkytr/Xt3TfuJGFX8RL88MZXxlpBW6O3YvmYszJasYEFPbmL1548ZqjV
kPHMB0djhIAedUe3hNu+NZVTQles68hgeJDD311hTpf7Vg3YqVESKIpw6uuMY7w05u/39H8fd/B1
AAbn2LxM3EiVqVEhFOnl4nKgOJ+qHfGQ9hFYgn6BXhiVn1yjeHEPbd+ox6ngSLB/DIMW+LhxfcYA
Y96xBhaHBht3/SnGx4vkfjvWCwml6D5MWoGXA1QZBYbufAOyI/z+F82fbquayruu/VHiNSMOtX1I
/eiw1sp6M9NDvczEtS596PZFtnlVlaBcBJ9P7VBHHrqtEfycr1i0uF2c95ag19B7iNBcB/7InVnA
vLMH+0jX/R2CBsU6w8oZAxPlNy/BAplOZUHfdy605hEkcF7SwYtyPAO/ujKGnsTBfSywg9a37p5Q
PC4/ALaEp0jdCYrH8Tx8KxyihPT5SaWFBLQji9s9FcmPH2yHcWZBZ7avD/lolqHX9+NARfrfFanH
aozTNCtK6p3ULRt9ariHdKL02N48hIYSHfozluyoJsiy5ceDgEbT1tM5PKY7wJLRaoz74TPFTkd2
ZtqUbeRs58Ke+t3A6HiJyiy/GhUFhq1q5iIHRXOpwIw5eNpRgL4Rwe7oicPSJ+FlXOpiaeEaug8z
xV5ZJ9wth8XfkH4JpC8JRhNQOEzoIYBMbvYohzBz3v9N+fNH6XG5J5QFgJ/DbaUdIbT2jV1zwYDp
h1n3jrouCfNf5qVvxa20nsDXE6ivCpW9XwRru6ER1DeHcJ5ca8y2mSqlGbleDKOclnTE8BnS5QxD
vfXCzmH5KoEl1SnzE9LSg+N16K37Ee2YksE0pb1PVbSGver9BpUQoe8sW93objPnGle/+7eQT7aG
3//NA+dCqg4NlR6HG+l7cmv74GtjLCThThubxuBxRvzZXtm9SKlPzbDl2z9s5adjyeVl+RP7NPmf
2cQJAQPtHJKGHZVUw5v3NrZ4iggGHlfr1dv0RG0c2frirUA7mhbFejmlPZZeGjJ+oRVOlKob1+0F
OMy4Li/xilwbxiC+5WdVcVzXVSo1MsmTm4LXXoZ4dYoC/FQY/XXhlJcFBEKqd7l9CDJBCZQj7fCW
LWCJJmuTETcegZPxX6P6tp7jq08OQ0SaywSPkkoP+2lxX36rUxp92HPLElrmla3oJCuFSgg5NpQH
OF96uvy06KCg0D3wE2O/DEAckcR/NmPkVHo99cPdalMTOhJRskx1HLn8SFZ+BMjbS7/eKOIvkIrU
wJ++sqZbQvPQkF4JGW32CpTjqIfS8hxSrvhLl4t3Soljmh8IDXWfEoBuMMHuyflWQ066cfRjh7G5
kkAyDzVdHyg3kPkqY4GEtoPhZrGccA6fHAvmISmhw6TMQjxKIJBGIDvhML8ZEEadc+ge8mlYzwZs
vjRM2GQCTqN12mA+CrSx5CFDJNQqoz9YwbFHalYPO676irBlwhCfKfZiPiZDggObc831AMqXUj54
fwxHyZlVed/G5aA1/TgdaOqmHmTF6uktWo+9KPR7WWbEmAMbz8jY0rciq4WKUzAFPClkyJc/fr4B
gezNf46SLonj4nyCWC+cPxoSmSmQajD19oQZcr88qAxeWY6k+JkvA0qBmZhO2b89wD/blini0hC5
GxwF6Htd5Uqmu0MjEPvfdC5Ml98iZIfKdIs2eb3hKferEYUaFspAU0jJv9+f6q7TLwAiWm0JmvJw
/sdqAfeoBWeKHoUcQWzAy2ULWhz5aWszZRvWBxZSlNn5S+wIiFSxLl8CBQq8AldGzME09GWd3wIF
Jt6+fQTJ+H20FXUm0JkL1QIfJVal+eGRjk2sxNp73cg8EjOzfRHu5V4aTPKi0G3Rc9SQRSRCVmBy
E0VDgJAUVgipSiuD4fhemZsdjo0h1lEPovtSiKtc9g7+TLOLeN0kjZuHSh1yNb19QVTW4NRqChbM
fJWV7r44cM2hCZTwjtjuY70j4phakIU0lr5sT5BcgBe137CX1MBVx0cKGFMwCB0J0tgr4Y2iKohy
sPgOQzTby1voMxvMD+4Vc9TPRa17nxhfxZm8FKN0XDUyEhqwUs2BzEJdzGmaWIvHCkIYlE3YaRM8
HWNTZV4GBoBtYMMyOwEhL2e2zkBjxjmUMEfYL8WXZv06wH/SaksLDmdR3QWixbsPr29u4F+gleju
fvhykcMLUY3K64Dcj41nbaBfdPLhtRymGWDi8hM1eL8H7sK7LEJ7/23/j6Wbg4BkKuVlF9hhUQrB
9tlpueF+F5Mmq+OM9/fYMJMGqgw/0ghNyUmqq9HyOCwYhXatzNw1AYib6iRyISfr24C00daKGFqJ
03VG0QzqzLKKnwrEo84PlZNowB3xm+4zbzZmn/VibkN7fWdB9/vAY6kBG0fTveaFg/XFe67YTjfd
rhDrLuUYj/ENdojWujbMBBspjTMS3kfQMZ660srFYvf8hrtocmqbHEIfcFrFZXEBAYzMbZIZqi/Q
0hKFI08mbMcMXqfxJ3y1KXQtcN/cyoGfs6Zu1DK22P/AUuw+cdbTxjaO42tTLp1yjN+WYayIJOlz
qyXP8HpmzJnvYqsrb/4D++yMW3FEA78Jz6uiZEccqqWmc7ABU+45Mpm2bee0p/zKngzQF+WrfCwS
jlufv85zCCZOR+TwIPRo7SXlNPAnvihj/wxO6hfis6ZgdFcN4uOlVhMFjr5HnLJaEUfs5sEQttPk
OPRhPZbcaDGyEVf7TaEt8TWjvcyPlY2khToJ1OqpSff3mxY89N8/0eVlSxoGCvE9K7+To9TBE1xQ
KWH9IMjH0dlYUVdZZjv2G0SkIgy+TQEURkEnifNAb1epJaoAep9n4RRwAYPtByTWgGO6wl3QoWjb
kKdAms1ISJ35cSNPldvskITrPin5pjm+/Nqw+epsEFiZ83d+qCSAX48T57PQEmFHMoxQMckZidWG
RB2VRRANFyIUV95YZpn+4/AwJQ3sXfd4uxlDayH0gXaz+rIPJUQ3WdFCQNQ1lrLLI/nvCMQOGyuh
msBu5TjsqEfuN/lwiENo7ozSGLLyhAUWquScAVh4/E5kLhyrUwi5iLS5lFeYTaJqjB3mpIwbf6pO
BPyR+9QwZf9wee4/onIS1ZKzvwIsYcpjDpGD6NLSiWSDNIbFgnMeuW6IDBR400fuiTJnlx9wmL7+
AqVOD2/VhIFvE+2F3B+nxysFAbyGn7r/iqQe988X7q+2AO4naNu3e96wz22OdNoTo5DhrN73FrPs
Odc6/1PdB6kyvuQ68EEC84akLaCTotkRnMaEsT39XsOKrOXtndk0tr4rgKTizrn8g3+TR8iVIteo
aabiZ4DykleZts1qUWjoqHba8VfSjFeUvkfqHAkSzZY/sA2ReEpPV4Zt0kGc0JPjmbkfayVOAzcx
RlAYjj39lkqzj+6PndIH1hscQ2VxNZMgexE17LwySBqkyrKiaL3aSFp7Ri/sKBOL0mN4TOYHfD8T
+vdw2PCkigC0dDYVvs477P6Nvi/Chw9zmUHPcAAe1A4eF8ImKCQ8/MW6P+cSnAAAxk47HjOYWhxR
pPr3MxZyVteI5NiwE2BE2NvaOmmwvYnBpxdaOXw1Wnd3WUewSb9wMn/nI1jmEl1mZ18mIbWYe8sh
4yVdVn6q5vsry7arojgC6e9sRrMWZWA6YpEwNlrm4eweqJfGSSsdpW5yKS1ShuunMAUPexKmo1r+
/WozR0JdyK3PjROxOt70h46/vYoZV86/Q85ARpGReKdNtwZSBsnSQUGRk5JtZYoNICdaJDsC/zw1
gT9A2qwlZwvG8c1GyOu5Dv2p64g9OTxG+vGzLBIFal8oM2Ize2dLBWHDOXCraiqnx2VOSDDzK8Nw
7AwQMSMs6w9rrDzbkT9u7MihVax0tXppZ5ONqL/1NCNmbzYohOr2PEUkw5ERYFIVl1G6RK0MBJDg
RkdTcCLRkBMSrbEpAxJhlCbBJLJtkGJMI1EnCJue6jf+zmWuFFaVUAfpvsl3mLS9LSt/SnxkIGQX
4OJkG1Ljl4fFcyzsGflr/pwNugI9TrlrxW0DntT1FLtX/XtTG+TnAjPTyh2ofL+BClp+ylQU+er3
OB6q3pbYfTfLcLBkupmczoDkjJ6U+D2NLhuCDYQ63I12l3QyYRG1dRzYdddufUf65C/f8ePHQO0D
YgQ6qIyJHMJOE0U3A+Gtaevlk2cz3sKggFPyNGWPGUEDLJAFpOHR0aOmVtzP2irxu/TJcR+uVzEv
C53oLbXC06bZ3kAqpjhLTvmy+1C7pOZTxvW53FTqE4B7UnUnYgVLzgCFigG7r4+HJ/MosbMLxhH6
Oiz4KuqsRZu7EbspFD6qh+VI9nfHLlYFGXrEy86IclWwEkwb/hg/UWytO17M0FojB/AwKfjTrFip
U73gYkBGeGb12p2XELCLNhkqI7lwr95Hyki4oUFKGKLjs11esCSYGccHcTnZOiN0l+dP4Ywkplaq
qudlT2lSD7kkykxenNurcWcvY68SeBcaIMRiiaGhqh5WBD/56cCgmr9WrkSm80OrJoQUUcRDsxn4
r6cWErMxx3t3heUSq8Ezi6XqqqRuKPCqk0Cn3wi0NBR92nUAFOP11G9lkaWFdbpc4S/YzA+cfZCT
tgnyrUAeaOynMZRm7IJ6OxBoVH3zLVPn17MWX7TBxMsew5Z3EfxhxbSjcoO3lyQtT5Jl4PPBipBv
QLCrv6QOiOhLhjdHyAI9XHeIWDChwWCzD50MLOC+Q/gKShTF9Yl+ZM9P0HF2paOrvxddeiDYjlLM
Uk5RcsOWeM48NEFbsCoKXzj5jtiMsXS0H47Mna+gE6y2j36CwVMPUFFbMNG6BkYqBFoWEzRWxAEJ
PvOP2L7qGzrUNVGPcXRKxKx82WzmlW3Hln7z6NsmI5NIkzIYfOKWRvrAKjBJi4gwFpk2uyMXwm/f
/wbIMiAmjBlzCVYYMhKgMv/6jW2iXp/UaoyKCfwZzGNF3T2UwktKUFx704qy2cCGTcA+Gcjx9ZXe
fA8f/zW8+z1b6e3ELcQ1eMTFNgyqSkNweWucpXMV8OAynR3vyXzSkKIc0srApMDFAC7YW4IDmtuV
STEMLb+EIOaEYQGCNrY2Ap225bTKMHVSpr/kHdSs0cNGTRohVKGBx8hS2J815t9LqkQtW0Vp2BRx
TGFWIS9K/DxZj7epv9tbWrFXuO7vP2Z8lQQ92avLtVnhPCJzhGlQdeTYu0LgsGyd8GP6Tisro3MN
BLZ4UwyI7juLrTzet6VHT0/PcLvGtIW9+oiYl8nh6yozu19kDItrPhEFAYShA7Oz06RypiHrrIgb
+niiKPNYMYZv4Ge1mEzhCS6fO2dL7MIRBQholZYcQ9wNUcYvhUlZnCOWzm5JnTaz9z0Kk/UX2riq
/YizJ2aQk5O4yabKV+JjR1E6GY88P6BEjuVqKxyMAVh5zoY+IhuO3AyWA0bhw3Q1VfwkWx1pYtu6
x7lREXHgM6LUbnq5h20ftiST/7hICOli/cmrh0Ixlx134L4sqB6jmqnrTQgq7rEPN5BCEoPrn88O
ePSSeHKGGK1OH4PJdSRIHl/pdMrXMh+P/5FOeiOTP376Tlrfr+/w06eBJuJzOTbeVUZivgDCFDNj
+N1ZKr0D9PSarTGMZEuadSWDdKUJnXgUL27XNC83iRTG8a0pdxZUlbAeTfMRBbnBXW+g4QdM0wXS
DgO3WUnKLK35mbYNqHsu/z0ta/AK4gCi3Bxcli8A7xPFBpJyPK/B980juX1zhRRBevyt+Fh5xmf1
SpAi0E0QYyYTpbPdWhxPo9S8mwXsMerH6Nswo45ghYkFA8fec4GIDHF674MdAhp1b1Tv7daMhir8
3u/sKkx7VMkkdA2TUW8tkGnt2CDLlYPjGYv6prpqTK1SZQyXU5SPzpwZRtALUMuQXH+Bgo4UQPRl
/k/Ia9lSIJPf+L5fhBhq3P0xCmhl0LrYuhwIg4UGgsFb6yi2nwRkRCkTC2ZgR/Xm+nZmvhQAlPA0
KLP/j8Eigggm+wXySkEH3haGHEOjBmGjNCGJgn4ArPZa6hCLmv0E/aJiipE7pMmctmqRH/Z5yBWM
VqqBAJOuP5mfEhQph+FoxlCNLg+V3bl6czQy9vcRVfX6P9kSt3FqRiQrpVwb7lRumIJ6HDNFf5EO
LeSS6u9m0uBJFzbE3wo0mKAHa/6NeDTIdbWp6FaodsiKgij2xFHPU/XXAXqTd6yQNfLH3+Q3ZtP3
GsrUf1Rv+S9AAj7u71wIxhsyL6lV+0VxZkQD7+Q/VDKEwA3sAylKEPyWYOA6WlpSpulAEOdOTVw3
zT7cHsu8eONoarCmc95qqvri5jE1G2zHR7YABvjQNs+kaxO24i+aC9SdJrOAHlczOT5tyOCKa1Xh
CLSTxmn5STAb/7Uy/A2O1nqrg0g1QLDx4u8XZ1P/UAjVuOenmtg332xaScv5+GTjp/eLsxD1xKdx
FUBp4+elES2NJK5wHYb3Y1tY5G9aCez/6485NSTYZnunlH9uJ+HuSPxP8x1QhpNEPaW8xouZPZLZ
ylbC9Wma0U3m8zB6WA2rME/zVCP2CqHssCrTUFVR9ayXrRM1NAlPrb/g2zH6I48TnkmESw7Vxp1Y
vP0/WB/TzEU2sM1+ZuHoAvgK2IacV4e58hPoSgG5hgFsSToOc7BS/h20eonrYildXEzvxkR6t1fA
2iRbPBf7Y8zCdHd3cdLggS30uYyK09Pyjgv5ZVzkxtW3OuK/9dW9hXevpvnyj/skaH5X3xN6DAKB
cWB6SLAsGsKNjdtkfjKNAT8P1qDY86E+gu7VJRTMrYC80wHdRipJhZY43OY8re+ujhy3Ld3hZIgq
Suvzos5p3crvb7c6BpY7fDfp+KG5XlkATmRwxJDU68DBiECOy4HZSh73Z8dWiXusuMRzKLhiP0A0
SpQY5lOQodZWM1Jmmku32MsrueWDqzjb0WIIyJ/TlOeSbDOWq74lYU90GOgQwKua0XDRBAjyKAIz
a/5pa+hAAeISr3NYxs74gz/ilGNnP7WCr+hzC4b/GP+lhFpe+Bqpm4fd/ug31kKXqvvxz5jel46B
LCBKnto/Yh6J1ppFzwHSaEqQ7nrKO8CwXvyrCTLz2NHcgf8RpjXefVkBSopJSNyS35hpZ+BZD6QK
EotSoem0ozXFzxYd3lnJ49dHv4hZxa+wEpemwmTQ2R20QEZy78SaNHJeEwerQydSjpZ7IfhjHX8M
VmkbEPOwug3YTMZ6jfc8u3IQJQHkuhlVku9tMwXjLSH/4Fb9QhoMEBkkMsj+a1jvjYaOoTabHVK8
1onPyxU7Y6Jnt4j7zMEJ4SkiGZTVwbisbYY+k6OIDl11RozwkiZTPHVwRmECgaeFW5KbBmhGIpo1
+dMF5rJqq32XtUyoQlZEiu+mlOATm94Ye4QYS6dFwY4PsTwwslqOqJtN1MTOb+vPndVgzzlgLWFI
OjTHgTjSaznCOrgQUmfjnrIwIb7TocIP33T3wq3ENPmCHooegbjaiDXlcq267YDHGCTYFw+gxfxQ
KIBNGK6L32YWJPDl+xHlpiQ6wmKvQsNaJEmVlwJ3fb6nBPt9aFRh8opxHca/q3KUqsh1BG4Ddp5P
ACk8kPl2LnT+/n8s5qA44abow1DNx1deaNkOjnQ5iTHloLfXWywa7Owi7xMvxN+4kLgTSUGuRPrP
XnMineR5BBdiUCTzdPgFeq9ebz5i71RyTB9/y3VjuG5FyUnZXtgt7m3SD6LgTYethiS2pclOgUh8
V74fhozPZlkS/xJCvErvtTZjAUM/+mEheI0xIF8eC7JH6qHHXhydo7glvAFYP/7jF4t3suKCHf7G
IxY60U0HLerJFClQBRTkfb7BajuT6Ni6l+mDsfhjQz5QOY4bPOO4Lzr3B5gjrw0xpFyxLTLi0H+/
iFnv1nszYzvBSiEA01COBJ5E3DSd/YUXYfnJx8t9QIT1Q+7FOgrweteRmtmlUiLTOaHQr/osOt8X
cre5d7mwHQ9GSdTJ0CaxCVLBM9Jetg+CZ5XqEXtzzutNA1QjKHc4mn8Ztv9+ZEKR2NU1NTknf/Sb
/aT57fqBs5cXg5hfmqICWLDyMVuve9MdWSLP0oRkTxBJUbh36GVM3uD65EdERVmUjOkc41LxuU2l
YS7+jsPXB/JLdLL5nP4h5M06u7zlBtWSAsqhrLiJsF5JiJWB/CD7zMLtAM8Z1vifx7Ci/2BD+UtM
nmdMnlEddvCioPwKDY59AcDWq4ehFL19gJRLd2jYvdSgPonT0EnS61tK4OFiOcd2KixsTZ7CUOpF
5Ym39Vo4fv6/rSMa9BWhHV9Jl1m/1oQshdbt7UUQJxY3Um2MrK82oeXYFk4iHrvvIA0umTXChyjq
PNdbUAQARCBjIeGBVUwAqy3ol5LTFw1V9fXYPxjWxURWFTTEEtCuL30bto9rZydQdazrL+WqPW2/
8oiHu7+ZJHUhQD2UVRi2XttZbIHOl5yzPKGZBt7ONqcu5/+5RV5nTsgHT+d949yTU139EIQLMhGz
Dbmt07yMpnD77CthUseW1MVrXdUJHAy4iTPJmh5YNZCSO395Uw9neme46l0AGPMDjZX7WQCEU+3S
HKEDBWZ/hcjGZXI+qdDOs44CQl0+YwMEQlZ9+wr7iDHG07F8seF6ygAJSJqfzpBhtLIKAG0qFvV2
4cc3oY1fxPFBkr8Z3XIHZwWA6XNIg+PfaDhML29EZylWGXwTNJFiJlXmJssx+BzZHV46kLM1WSxs
8RcT2w8/innM6m/kH94dAWONOPlirLBupmmqdRbWdo6HLytpGm2xZykj5tkSPld1TwUVlP98N38Q
Mrl0WTwQh4N4/S2Id+v0IYjzxdIcbmdgz4e5GvTyutc4FR6vIAX4yhm0Qwuy9RTIXzGxvtenWFau
CzoO+XppECrLVayybU8xSAucxnF5EWIm18VkN3wf/tiANONJ6BE/BA9Cz50NgPqPPjTcf5aW4OEH
9KTVwAmdqM8Uf4JCTT0v/RaxDPLWsbLU4Wpj1hVc+1UWh3G5BFrx5jjgWxxtr1/5KkqbObUxQyql
8yyQHZBrT57PY5NHdiMRHCwAe9NN0tzcdeHWUQ0HLU15CbhZGSPjnM7x6sYZVIY96GAxfb8/1H7N
srHZ/D++ArKbR2BhtI1AyXrHQyS3U5Y4/bFpHUclP30ApKyzBy10E9ymBji9NgHAi2d/wAdU97KX
hOdjR+WmiM3m19K9rPLsTNYWJew2YB6ZUkp1onTT2pm0kbkaKy3hPKkI/LiB/lQCEh+LPPWCHGaL
i43HNkki8TK3laqJf/yibIJyp7WoiinnQRm9TkgIW+vmQOfO0OjfQv9vsaay2nVrGX9BrD44PtVw
5WdKtEE4SgC60xz8yGK0u7SnukBijDlliRXl8qXbUhnR02QPtSEqhA/f3/d5sKKKSwUj/svtwsk8
eCy8mB6D4/EpSH2TkEV/Ya6BU+kBHhJDbVxxs294Sq4YD9iZEdVPKlcyTThDiSnLNuU8fFf7gVeQ
NMn4AilJgJyko6fWowlOky2OpNQEBTQ0oF5x9SOfgL4zdIXYYgFyEGlj2OK4PHbrTcYHtP7Gldnb
wy3286ZJdP4hqzmetDtoDedWpkitk0Vz9MWmWTdJ6FaFIQj/A2gFh+TlkHKjxPnNO0UxPger2vaz
pEL/8YYbU+CfpvkweVIAqQNN/kPXOgTuMoxqllu11SpI8FS8Mlscd0cE9fLsgrqteayF+RVSF9pW
/IQg67tquNRTPHi0e0SxmteifqwCxWuS7YznOXGLL+1wyavrXZqp2sC3TfqUWNpuIa5SHcTlfQSW
PCH2hqsGREX6mupyoZL/mr8rgxGtmk/MtngefUQRNOE6RgtvjDEiNxJ7r/9sujR1n6ZVfoR43ZyH
ho2kei78fLGL0Ed/elSwXw0jm2l6BM6gfBxA9aatlp05TAp1tDj3lCJf/bL6jVJvlFcNkinbAjur
xfvwrv70xifa3yMnzF+M9Daja9XUQBigNOuzWVkAd6I+Od8+0b4hXzGDIVGO/MY4JtBqSGHLRxZI
pmFjUviLVqDTBNPRdazhPN5DxJcswqmVDkgxulTKnGbXDOiaA09uMS2calsIAxMakOtVMrfkLJtA
gtadb7G8dyAud0S4eK9c8e+kNNLNOm9QQfav9M42JrenqyL7cYfZcOkLH7grA7J5xsV+yo3rOOvd
Qym5RiGHT3yg4m87QWTr8P5gProoI5pan1ugZNtCjgdYuUU6cOAdTBHVaLceejRd+ZB9KcVGIbyS
lK6xQdgZLq+d4lMBPjrV6s7FzvwIUkqoLbkf+ysQMHRlQYgVftoSVGy+oiUw03glKayznCroi7y/
VXfYPhQ1FYjZ7i/DxTKWAqNOMsk60KD6IGkcKCZr6r+p68aupDCWouxNsnm1xrwv4WTbhZ/MUvpb
R8fpZtNIx3wcsuLwSBPeVqGsyQWT+SEkTJKF062icWPSkpsJRFqp7iMB0XsMcFGjCK+BqwH5s5Qa
B7RfMQHL9dKcEvBgIeQcwyV6To3r/EGF/NgBNKLHJEg46o8aHG3K3VwAeqxtskzZXZ8ysGuU09hJ
dbEiNlCR2nJEG/ar1lXmOy3fxgL036CL4z5UqoDkhU5x6H0z1oZr8BZEuPHl3QAPgTVfVFuZ1IoT
8mOHOJESYLiDJ7Lbr1zC/ZUmZmZWK/+4QIuFyH2AUNykaTyg6no0dJyHIUilXAPvUoCXYVBUlosC
U3L/TNgbfRqjmuWoVmoy5531iZJC+AVcxCGnfMZ7X2Lkzsm2pKsQ4U6xvpsq7tj21m44mJU0+csl
rie1N1r9f3seuj32/nYOToWjlz+2krA1ogSnQneSBDpinL9zbb6JADS8WJw2zEnHO+qUHJwego4z
OJTzBhFT5E+/jbk6ZVzzs5P1DprQsjvw/H5XFhKudj32xKuQldqBafKFSaBjLiVd9BJzu/nW0q0c
KgJ3z8E0/zW8cWjEUi+wukdmUdUob3NYwH070fZEXdakelzKgLRAaz2WdN0WsL41Wez1Wg4fdiIS
qADxhLSsnhyDYiU5p87E5af8Q9wJLjfO/83xpJxm/el6OoW1gLhaJRC9yxT3AalcGo7S0jtrqvdq
stMUPQ5G8EqG8419duu7iwMNt1tGVoY72YdBDtIYGmW/4t7e171WHjttdxyu3t83+d52iK2iqaah
0xSv/VRh2Y0N3CHvxfVBIh6yZHISlzWOt3PfypsOnytLsp4BC9S3XVIBCRoc54pNHoPeMnhIcNUd
MBZFuCO6dsnnNr7kF8HO6X05OtBiEfeTb3UW94CJ06gbjl0kFV/ZXWN/15XZ40+raaaVssdHLiP2
vvoiMg70ArKrtil3fwIzpSP/PBsRHcn04GAM5aDhU7JA5cAtz4qs5xrRBBZ1wgOKC9b6WeJOES+t
BwVVCKRaAOwTCNfckRLRCWcR2hLk++XoT4D3PK5yMYTpFt6bqSkU/QAyYsctduYQng/tUUnGDnBK
4/GwcXnNUUnLIpiNGabG5zY8f/yVX31NsjQMmTZJZpz84aU3wjYIQdbMdVJIjb0nxRzhP7/I/roE
b7QrfIQgUE/cC5x5wXMDRjajGKwDkBwKqfD3fq9CZ+w7puX3TT5zfMXxy7vfL1kwscufSQSOA2U5
X29HAk2HdNx4ZtG7HeCCaJ+Xqegs0nTjA6fXxjiQzVMODIlngy1coT/QCK+myWf44TgGE4S1o0qS
h/pWOh+j2a0E2ovN/ZmiNcYV2T/fenybae0R6GQsioWbjZG6RtrTZPTUDZxjtw6On2KltPHqflhE
o71/HiD2ronmRNzrWVrqIfmBO1A2FIXjNyvm71NrOcs6Qk/72ZSOtuufDE+2Au5KmJQWrlRHezZK
Ukt/wrp02mJOGD8QDvQJen4jqMGgswS/bKeWCG1EAZyTP0BCiEw8CguzfWXXqZIRgvTCnVKlJjZs
T842fZnih5SXcLRzzYeYnLzggrIWk4kPiqtPArBnh3yIz40lhBx5epGewOTJ8RhsqP85OITEt7AT
P0mqFiVkhpriKsxf75ODFruhOzMBveekOfKM5FcaIFqG/s6ety6zeAPqc/WY+uYP7yS9zZMBoZCu
wkitNdWOeS2Vpe/sgpM5zYyrrmBf96gwt2sF8XfjdsGcFH5iO7O5gWWRm2XFPli4ohbUmgstB2ge
xR9haT/mRTDovdNC3/pKB3EUkRfL8tF7neOS/L//PWvuQabA/GMCIv76/FyY+JQuL+m/Fp3X7she
1iLku921vvNyqP070OB4j1sKSNavOriKlYhPUATx5j8k7f4ZNrjIQn8EmfUYY+thrmmfNBY9xYVU
a+6DWN7WLMcuichqqkVoNbUlLsyPAi9dDnh0tk0k9bug9akhRLEXc8EcBGhimY/Ky4sNSpJs/jTb
zKYjnWL2qBn+KWWauBP7HY2MsdJUYcsHNHF7Gmka4NNee+2ycYuQF6nfKtcBHh3bw7y+oJSx5CTQ
Jh88DM0dp0+1TfzkrtLAE3AZKVGR6qfdWPwiqdFgRYV12xqmUk6aQvJnIe2zsjRfVho+Jdp2MwHu
yYRvndjyTKQdjb/nNNu+I0wcasBrUa/J06YgYvt2uoDa4PIkLUlWDeJDdMIq+egKeO86gH50cOnc
3qhRpx106tq6ZTQwJQPqjTeEeaEXQddLSRuN6bpkOCLENdQ+Zzk79G3X4yFFBKGd39Oa3uLnL4Ri
TEy7HfMGW5KJyGOIw4UZrDIMA1U/4KR9hhjjUnJs0UvTPe33ys/P2hpK4j0p/Lrm+IMGkkGh6Ukj
0LBv3WKXAplnaaO/sIqaIwc3bXVlaCXvV/KhToAhXYXBFIrspwUXGV+pHqQf2E13Rw1tFcwCuIdH
T4fKXJecEJKUCgqsPfFdzM0tJE5NAqTImP4K+xC1eJnePwf0SXAnhjvr9LXLgsZp2OqaVqQj+KOw
9iv2mVEEpk70/kGss7BSMLBCTRmUzZEZe+aAy5sANUyNuW2IWIARxErEjkc6t4pzzYlvdf9/v75D
r6mpynkIxRQe64pe4I0908GQMduk81+ld49RJMXKmYmlytklacjACkGKn2HL2gsruz+RYsKo64jm
JJoBkskgnEskkuE86wD3cUdgT1ZyLQHh2d6MQ3usClh+BiUQz5/Ip9Duq3rIK2evapOfApyvmCO8
xVp0LGCCEjcw9lHhaGVhO9Ion9T+/2FNIULB2kze5Fh3g5NCn9j89lIZFGqV/iXJukLfRKXX6H5O
Vx7YaAKwtCjthTLQ4hS2jblKg6Frsjn4e5i01KdmBPh6TRPD9S4zdClBtEODyZLVUr0Wj/BHlbif
M4fCYsGRWksAxJOFSNSJ3AbcRXAONL+a6bQ3hKsnGDCaALNUxyWV+LNiT7jm6NBtEe5Ecomp3JFa
gvspgNmtdfBvRqsPgobvVco+HqLkEZZmgAGdNuaHp7tS2BwFV7TpeI7XDmGqbO33OUVmcMoVtu9v
p8g9LzZfNbSt++g6/woP+6herhsgP35jADRcnH2htRQ3hGRi48HWDp95c8jBK/pIdT8EhMU3Jg/v
9FPBmmXKuwAyVMN2fTvp4PcZrefMMAXJtp2iS8+mcHyquadZ8RKdYRrYG2oP553cdOucRId3z+HL
Dk4fqbnmBhkv1ezbQ5bLQclmxtFwCgMdCTlz3KUr+JbQG+4Gz1gkHNvSLU6xlLke9Oa8iW5XWd0q
YBFTn2HFTXjVZFi9eikAYn44Q0bqfFH7HiOuN6ESqgR76S23ezzZMX1CIR221uKHdWwlFRxTuYcE
QDxSv4WumLX5pAxqV5xLXcWkTXUAnbPrm7dOMEtgGk0a+SA18zwXQIudkoshLUaQj9RFqMh1Ddm5
mno8muFlXIuzWSQUkB+/Q/QozLGIxBVuqFkTYAR0CBKeXH6qoXTdTutbwzxQk8YXtumnBeO3X7gF
bK1NDDRoI4bB85p1f/nEE08Hb1BNHUQUmR2KTSteWmRcJ5gIiavDLfPtGh96OcqKGpOgHGDeWcNn
Nt0wBPBEV72rTXoGbq1dviyPl/Y7u7rYtzsDZHphricX8KzriCd3//U6Lj3nttojmKUV2Mv0i/GD
eFDzh9oIBTJnsJ20zc5dbq/HMqe6BnzvJmf5jtzP1Jay3s1IrTc/ROlLvwSuq7wJAIDqvDImH95n
7uKjQ2Ifpk9yHhQkQ359DZQZIN5QI3JTTqxNviqc6hqR6uCiarvrAFYGFo1hf4m/P8ShjlN3j9mp
pLAWb53FDpO+wxB6H+tkHvN7Ys5UDMt8iJ0FGNDk3eX7+sTYjcugbSU7CILZuledD8ieTGAb4RYq
abqy3IHdf8yeeHaFheh7WfxoVQMItuhkJDGFSvnpZdwPQNF0DhRCcXUpTjbTDrv5vCJYLUdUhy0r
p8eKo0wY2/GtXtyVO8thA2yPq0pqdihIuBqrx5iycwtNcUxr2UPK/0+t85lvE2DwZJfDg6LzCmmD
th8Jz5+AMpeZoU2jmiMwF9aXSz1xuL9TsATC9DVGRaJrQmv1DiTNsJvNZxv/D/BewYr7Y5ou2eTy
17nSSCOU9g8PKW2ymkzqQbTCZF71aXdtPeR1CrT1O+/ZCJ9aL5uul6u6aXR4RXkp6UEP++eM/A2O
QB8r7vfNRteKhDU0kIVHAZNi3WOOiE6H6V3aq65xkCSmA/Aj8fe0Yio0sFRrl782Q71s3dMTeJs0
f61DeYhJuLQLLqVsDkLk90CAk4WCtO8OdU2UgAc3mrU3FrynsAD/fhwFMqYBeyu+BP28prr8PEl5
uB02HZXmm5wrGLV4dUcbWb5rnAf1L3Ba656hf6y/Q8/VGjJWejJ4i5gJUvELxtfhzI0xvBNsJNOd
8VfdrQQ72BANQo5oQ2dY1yyvZI3zLAGylNNqEADgB+s2gbR2jnx/wtvm+eLOz1y5IuoFhIn7UgLM
S9ELBfevZkSWYsFCX2bG2wjcESBXJ0TnWBi9PxJbdldYBRXzDuQ2Y2ecsbBBn9Rtqf2VD0N6Xi1S
BPuxH267MzOvO0wtJaqHi2kzTQ0sW2XvP8uN7aAJvM1futGt78ZqKgch2WPrMiRXmlos9db5ROFw
RWpwWfSpeKN7Ic5j+wwG5DAKLmaePlCnMWIhgVc5GmxwZsdg3+7K4AXIfFWGwOjget/4TiPd1RhD
Dy8WS+j4UovthmXPjaokZclXKm9m3lL9/R2+LfcIl4qSDeO1uORVx50OFdikuvlWlMRipzQ0Rubp
NdchJq/9btx/hiNyR0yUBxtWMMD0x2JuSAA+Qt3IOd2qcZ+sIHQGTIdOVoVO2LBDRKMz6QtlBWbu
6xbhmBGdo1bgduDiyZgVxiPwoJ215vlUPn2IYareJI8kEDBr8WyodgcC4JPvjRW2K6KIWpb6B/Yb
t3DlW5zj/uzvn9DjqKe9i7kmQGdpD5nZVL1c1CFktSpBIlY5icZqg9XPW5AhBupp26QSnIgJLQas
usXxyuyrSrR6Pqr73t6n3bDP5kgJVarNXdVLRLLdjmpvQOKP0eWMjSgbf8M33wHQkbo8TeWBWILf
brvSP6JEXB3WPu6ET0orrbLswYDq3fIar4yPlmQHnYpz9TcMIxGz5kNyAyYFii0wOIlUGR0eUE49
q7VcdgEWjZNXSnEsb9hnVSujTW+p0bL3r49Rm+kZCNU2oYPIrBdBVeJWfI8PwmZF/zQErdS9ztDl
YG+rTd5+w0YOH7nDm5rQt/9MtC5xFIcUFERpfnMTFzObAbeNIRQurMCjkfu1VClpCHWzvxVbgo+2
mBATLeLXINcZoEQkki1naCVnDbRfOtdqU4tuk/LSWXm3pYPWWRidIfB9u7Tzt8BqtZPz7s3fsKFl
kjVvs8z6dFozWJXc664ByLWN8had009dX+dff9PQ+A2QD9D02FV7uFUqMQzSflcrYVvxWBsv5a2H
9FZoDy8aaYjImRTGainKLCWQ6qyK7IVvqkk2oXCfdIQ18MNv08Pp+4o/tNK5iTUyrkHnrJpIuLmU
iDA6WC93RvnvoT7buJClYKJWmAKKcD9qvB+bk3vbh3lsC1bBVS74icXx6O1L/royp4mNqPLAo8AC
IO40fAR1bf7ZGjQq86YOJm1+DxvMJ8uf/AYpq0G7fHC6oD0S13HdF6CXdlb32SO8UgKVHy69fG0a
NgJaDovbkk0EV/Q+Yq5NLkyyMPEXP2XlvhTTF5dnHTXqDRsdqgKMH/Z5GouNArcT++UdjVPpTRMc
/Z9QED/rRFlICEW72hBJW3po9jIjygRqH74DqOXSOHa26FPRxv/BMC475JvDG2OEEziBnhcrcRH8
wEZP/jSq0ewORozvT7NL16LXPj5/TGVLw7hkhl5t7dv049nYkWzVkNAKx7PqdiRplEs4B9ilpdx1
qn5gLj/1v4rTjbbxZHWMZeTO51zlWzxGDJCsT6ncbkqj47VlosQk602GKxz2rw10ux07kEtAUhMQ
8C0+68zEhUvUAKpy/1eDuw7AtL2J8lt6vv0u1A6cph5Rx+cu4Iq3NV/DdrZudAnMajH1iVaQlqsA
ySrmKvVJxM3n75MQ8KGZwPWSUiG+b4kBqVjVWUzJHh6ll72PZks3eBNVd69yNBIkXN9tNBnKJ9zH
3UVI/rbta0Qy6TYWxUmmf9ksOcl5LQuk688zt0Xlbl6g5Gc3qcOh0QCRxCI/WEc+9n9jsE2a6GM5
kDcYuXjwF52nH3306oywNQWMS9gcMDgCGVWpOl3vgigOnsR1ohP/qKEs8oFBwcXUC4RXS6oQ8dSX
rN4OSESPTY7aXcOAWfn2ydnGVSotNz5MozsT2dkoS+JjwEDogb5W/ett2bS54j1PM+Q7x5/uOS0z
r8Tm9HQlWRfT2tCm81XtRBmFRoPyGgh+ZDnyN9AmHswGZBdQHG54QX/sWeKQ48lTjF3+WBRMVlhH
Qpl4vVEeKAAPBl0DVr84BupEFjn2WF59ozTkMWMm5XNgOKNA//qvv5K2XBqXyBKrzcEg6C35xkc4
dXkz9Oa+ar+QMxfvXSS3T1EwyC/hD7EFhOop6IxZLujAlw0rjffFgK9a5jU7yQWOCj6/PZbiKvwB
pboyKoya7R840n2+Iv6LoV0DP5zrxFScnSo4GMWllMU2I0YUNM36lC4I4xPWaHkvnaIkc7ZFxqqt
Kr6xNC2IMXZarg4X/HbbvjlpGBGtNgmqwq9UKJoJdSBScNFBsqlitOP/9ldld2tK1V4b4Yl8av1J
b8gdJZEmwcad+WAN9dYABHocggWotcnJm5GcMQuIDXQ5+6FaY3sU+feYet10+vSnzZtDcUIX2SVD
IEojwze4c+MyqMNXXRXr2A5QcDTR0wqSj9YIysTYpwFbxZdKgCGSJ2Ct5bePIfuOit4E1k9SHLaS
ToOnQkbxv9EaCsQuV/zAwq20lk/h5uilQxZwW4nwyrv1ozTmUG8F0O8ux84TpTpbKmxaBtl6uzTA
gQbP5hkpYL+y1tLsDYbOmHXUEMBCHTpdh4LerlBPREpbby9C1jZqFaQuF7gzBB4BnkKLhY8Nhzn3
+q7oOjrbHzV5z49fz24/BQvXm8+5Z0ivHUYkY/3Ot+kTERgTk7TjEdF0isOttZNvenLVRJBm25s7
QnWnf/kdAlgjNPK5keVpGHu0AFDBbGVtJEbz9/jcYrY46OxfGmZotdgEaFty4l7ZcWaIhU7nWiSQ
p06W1eOr8GOzw26dcLTG1/IOhL/QKdIn98Qg1SBgJOALltROeIeG5uqGf+vsjOrQ5m8mXf6vstMg
tBwqgcg+ICMTck3akiByRcNZ5uYqTzOoCIwKYZd71dHVXoo40xEX6LhdztEjw1gTApHD4wlkFkcI
HKpxDt9T4KHcblUl0LS0DGIS91iXsg5mun/Od4EWG3Dt12onIXFGHCkf7GF7+RO3dJAmRdI5H+OU
IQEY+xTAyCSt/UUTUYgpCh9CG722uPuQ78GL/36dOqMBs+uz5jNVuAVu23mbCO3Xfhac0hZSLtIs
eRFdcD6Uj7TURVBco0q7VKLbwSKV0wBE0trOr8SF50emiKnZe8cVJQEyIznI2W44NUrAl2kCZ/7d
PY+dgsv/BWKoHo6yn+DCuAiwmEW+zoTQ+kQ2b7ztAU3VSw4K1hy8/NeFA/RHPuFu0ej8y22hnGDf
jc3naqGY8YyB28sJLog8F7s3oTwKX8NdnFV3MH93pbS9e9ckXGnC4Ezir7wJUVZqm3QnD0BvvT04
GbtawAGVWSxyzgGny7JhzF9KkKzccgSou16L+kM8XP0dWSGp8MpUqE8FSgycComaplAEzJLYv4YI
f2q3d7kXjHebMmcgtqQFjIsRTj4pX2BXlDg3RIcPIr1tG4l7y59P2mxDAyWX28+vwGsXnVCBf9Ui
0A2UTc2B1R4r9Ta5JvITlNEAT0cG+P9maqltrtPxQdGqCh0ib8Fjj6g7Wlz79XD9O+guW3ICqY0s
GC8uLAdLs62IL9GZwLgEl7XAFsDX1c7VXE/2JiVmkjtGKyP0egYs7nUsUczpto/QkZuSnAb2rtW/
wqcMRf8QGuFCfaScQIYynqyamEdv6Z1RnEjN+FJFiMq2w0//08ABzYliI221gmqYhMhA1UtRxsK8
4OCk1Uz5sE5RXgqHrV4lrPYeD9NnRszVbHB/lE00J+6H7JFC0zsZMZOt9MoNksZ2yW5UF7wNmfzP
HwQ/vr6VJ6zIFQtmq6HovdkSNVEMPReNbwVFrAVfAmCyTnqR4wjMxP6IsYUM8SWiUnb/cjRQ3q4b
xo8l7hlsOg0IgK2cQ2DYEGAsjjODHxgvIp/LRisBEPg3bq55QEwdqAK4lhDDihgukk2G6hVPz8ax
So77Fg6Q/NmLoRjK/9lcDXfX+wG/zlVlVNw5fBAoE8WvAB1vlobrK3d/r7iNEL+mMYFVhYUDA40a
YllF45Vd2Th26EIjsTf9koFqNAj1vmUIFlq9Nog5sMiYHr1RnoOIx21nGuYJwzSs4o1oB4/r+IE4
T/Xwdh/h3rFsRY0HMOLjWX1R+gFrtYw3aBk0WvaY3hIYwPuu8kEDw+R2QUbzOY4uzOmvDp6JHau7
bDQ4IUuG4CkbPfpGyYOE+zek/IJbJFAUbnCOEuhAxi8Cw4dmtUOS4L0Yz1OPctLIAfAbxghshlhi
NwafhI9yLMSSggIDssOnwkK5UdqRHrmPyOd9TZDEXRlpufSn5rLZnkQ2VcZhvVviKDaclVw33Ed6
s+k8qrgxAm8uKhwfBPmDGlknq0310j/EbCBzXNcwyC4nk5Kz26CY4sbfqBurg5UZ1u1/ETr1JFZl
lW1j9athy/FMcs9NnrlV6r7RB3ENqjp6q6J9M1iHIXB8D9R7THWdp9Dcb5kcdGddFq/ovWPwx0k9
TP/IGLuDVCAjCAEOyoGkw4cytilCFWoz6XOwIVDZgzBz4x9yvt4PKmQoKw7DsQfETbLrYsQ3G+/H
/4Kmgb+FaiwsFtgreobwlzJknCIN5XGu7R4Qb6Uqzly7ypnoypGxpLAMRng4dPH+WOQQaOMiPY97
pizcM/EWJqy5BQxu4Frhbe6fbgbkOHiLem6VcxmSyN1/h5pqTkKX6r1205bPeshayiblhRkR6v7W
TmAk1foc8UCVksLnph5tqqHMnn3IdDRtua7sYIL0u7pYN0XiXuuN3y6oRnyIuE7EexW5A9QL4Gpm
pBBJQWtA4qEaFxR4zhcj7qMPrajVKGbi1zr9cWMzN94kJm3l/rX+b259lowtzaJtSAqj8zLQsgHr
n5qBu/M8USbuph3jInFu4COIwBvpdDaY3EZ2qxH4zOBoe4bsiq/f+1kT9TGjfrfo+Mpukdz8LgqG
M0mZWk16HyOzIoIkUYWb0jOpqQaztau8T9lbMNIUwfOpxrquV5ihuGWLAgdGv1PEvar8RBBwoZxN
o2coXj54RdKMMC7O/kxqJ9GC9/hf9tB9N/PD/ajVq+WCVO/ymyj0cpNEiXwFlhk1aV7ynohUsU3m
WpaRp5QAseqZ6P7ocfINc/BDgKtuYj+E/01Q74e3aegKiZ9HW02EUS+zG2sqMcT/Ypeqs7xVJgHo
P3ghYECZiinYML75TkzrvrWk3yZZSeRH7VzgfbG5xotQ+chkeesvDRU19NmFGtYTZPrwj07BUagS
HD+rh8P46yT+vvXClW2yMqRFyZSQK0PFKEJ/QOJp0+XJJOJTTQErHxjMdD8bMLoCGxBPq6rZCaii
6gsTrb2lOZu/Z0Cx6gfkixiSInXDZDYW5XdEY7BtZ5q0dspAraZcpN5wrjZr5yh41SkUCSh0Ct1C
I3WxMP0SjCXKd1I90+tZIvROkKa2Xigira5cphlrg+3BzrTLCT6aA3fZfFMAQZh7AZGHjLQ1qC4e
5eGwX3BuGCUcur+FRVu//Tb1j2ZLn7r0yaQouqrZ5wJyBRXhWzVYaqAZ/tUwcj/9OxdfU6ZsQI1s
gFVm1ZmOv8JmWNsd30jnW4csZ0E86yHHrXLdlCo+a80WPQm8drD/5GI+kNkOyhUdbpxcZALDyP/4
WWTfIV11ni+/Ogd9aOA0tjTQ1qJSJTfyGleFyMPvEOhgG1BQU2k6sGpTXOJSjmmMLXsr+J6pq9rt
hBNQ6rGqaVmZ8vgWAcYtLBhqs6vRgdJV0c++XJXRaNPf7Hwj3nZuFKXxrdfgXw7dgcQeRtJhXA+e
0zrU91fXl7yFVKypn2vL4/qdymFhJyCkK/RzyeTYP2blRvGWNAqx9C6sDZuv8HF1pHTRE50jpZzv
cshB5jW/rgX+7RotEimtvdKod0D54m5grWC+jfU8ag28XcHPdyEe+iRPOrx9H4BrJHci25fcwrOS
0J3mBQgUK3CXnAhMbmrhlOcT8D8fSBIgHUvp3odhyYbjatiSlD/qA3w/zsfCEkuAi2UOA40cK1mE
ezibnLtOUyZ/ZKPcMr0WK1V7I0U2lZIXX1peyR9VwioArq2Xd3EfhH8n96OqvVmAfq4elg/2e3VV
Ahx/jHiLyJNaIu/fcG6x5gLXkrSmM8Ebls2g1a8aahLQgWhbpKR5cIniA2VY3uFuz9qaQ5+VqxB1
UsmX7LLYRAyYEZWjTEVNGkmkfC5ThQeseDdR1VjcCRMdTXicFmm3fEa2pCppTpUIDZDntFPDHjfD
W+eROtzzrqTVTlQMvzIuYx674a8GIkCuEpWuNqd8TCsepx8JKyCsy+ihlnBtNmSWu0XaQryZpcMm
Lz+oOe3jYZ+fqELDKbdS35Alk1Es5n7RwIWfTThqsdqIDoXjYQL3quy2lsGewFGtcIpWUFqSh9Pz
15EFyEU7tzqwLYxBIlcappef3IyRJs2z7dNHIcCj1oBpeg4yAoresYSoxBsP7vFpF2qeEdOO0f5z
NR7VRuoKXS1rnzGN6VOCmTev1p1oroxBXB3QphsYHE52Yv7Z8xsJm3RAcTPcc/QQMRW7EbvIgh7F
OTCuU3dkConMi4Q6ggbj8eSdBlNkrT/3JzRXizRprwKW8ITC5b4PET2Ky0gFHVWnlAM9VNbSd2vz
g4czDVU0NeMUQGCKM34nS+hxMvH5qTPQ51fy1DNWxmX0AfcdAEJAzpsX+5ioekvQ4+zRMblUXozb
2eFNEb8wPo74YCU4oV1RKT2y22jfRkWqjV0l/yODAtfWVdp7gzD5rUl7gUHPqKfKWaoMJuyK7jYK
lsVEhvQl/x+spEl6kmfknHMd4ucc6LWm4DNW9lJakCFLffmx9rs0bU41ccGimDwF4rjDSoJNNq20
TXwGlkFSPWtceRxH7NhnFn8JkBllPCvJuSJr2sbvGXSETGn8yMjWdA0t6Xeeqx2hl9zA0hfKlRaz
HWeBaljJr15APem5AmQkNKmap9944P3oKEAWEb8haT6NFFaFVav63cuRtr5EdtSOoxl8bkmDQZRe
gYWSFi3GVeRTomDmbdx0ev3dnt9RArfeBs2Y4QL3QwnUdIttL1/FXVFBEtfekomzceHfFfM+ypJ6
ikBLMbsL4wp5o6tdcfbF87egYO4/cwLxE3DbjGRo36HAg/jZKD7MfG1ecyzvIcwePgl6/FRVamnq
/A+pKLMHjRZeIguPse0hBtfnXMizEBbgkIDgdxu03NuyUI2tf08ry09X0LtMzXT3LDY/Kzif4PSb
OxIjHzlQXKI6g4jqtyY+pRScPuTKDyjl6+oFzpBApJXuOiAqwRmix4NwyqvtL0q8NSjGpiLmEzU5
jBkTw6BxFS5E5G25P0Y+bc2pTE+JHuABDFHDEpx80OPTY3Senq2b7szL68J3bNvYYiNZ7z3E9ZxJ
RrcpkJdvC20AbQlBSCoPsatxBtC4v0Itsb3a2qY0rKRKPZcB7cb8WKl1JFuqA8lXxWr2zXWudRzO
XMBP8P91GwsBEt5Nt2AW1HT2A/hPmzdKzyMH2antbaeN7FpqhkNctECBCHHr3AyVunJEVdnCnB47
rcBT/qZnpZ0RAL7+V6C5n8hRiRIkZKPFSqeTSaTaGcbBBUnMFjNhlgg26o28XHfoELrSjaNBlXGd
sjCiWrCr/3WeIivNCXKK0qH+PArT3DtQBduOggSIiwqu9n7BSJxMbRNLeWYFsSjQVY2fZ2ykrCHM
4v+IQX7nZDRD7j7sVUZGI16HCjlTfyRSC6g23kIJDpj3stBTkB7Zs6+xxUou1jfAmfXsFr+1VYQp
qfiIbGh3iMxwMgtfiryynAc8BAsECGP4hZGboRrl3deZEYYu+/1lrGwHKnq4atbW1QHPqtRJLNpe
8PqEHe7LRrXqLAyIJ7qK0vpzLRzFzAUXxHMhRDlARvVJyVQ2eXQzuZa8Z7BVf1qRC04662eEtYHA
SEwZeuO6ysGD7A197m4d2v2+DTQx7q+cZio3/4qKxoxEEz3RDTBHze27u8RVVBO18B1xX+uDCFwm
V9tFL6K5CftWKZkjzpCIK9ak7juIO5w6U5PBeiW2FNFXo1PPl3eBT2xWcvNLVP/V8wMj2Nwv8nGJ
NBL65nc3zV8F9F45hToTEuL1DxGEfGPVxjdQdt81T3NI/PnT4njx9JskqFawuuKTmUpidvBhprfN
fDGzhlJ0rJhSxLtsk1wRGWjj/OESrIFH66O9PzmSroWiIlf3nFOhflFiSl5JoGng+iu+hTIN+t4O
3Ec5/Y0Byr4SRbcTmASdpYmZ+WYNSSFQzKYpeGM/gQZlclGp3fFWpyYt5ncbCVgW/+rIKUwpxvWq
ZmyPQ8GEt5uMxBfwTCOb3oCt8heQRW/UXWCLKgGlGJoj1vlGIK/6tHfc2lPf68+pIbRs8kT3IVgI
kW9MjGScpV9T8p/zxS82jEt2Ff7sVgXax1NYhG8BwHOLBvJu7qsZVtwqGDNbVBz5DKI5td4Ldelt
IXBhDocQv1uVBikRxDMbj29UKYQFAKitj8D2M/INXGX3bukaVSwRGldt0GmCRP0hOifNu1OKo5XE
RH57e5Q657TQ9Gl+hHm7JkTBAe9WVofHKX4hOOlBCoHojd1/WGtccUbTGXXn2TluNrRdnd3BGDWa
05MvBh0rGQSqNNq/JxBoeNPkDqYM9lqEVN8Py5kqbl91ADqvKedaw6HhswUDy2SDzoOBz9vWZH/s
iRpiaPi4+gyQOXPuYwjmNkZXCLTHwPmpU7snDKKf7qjcmcjaRZ3tLNQAcjfHpDG90NYT/8yQjWp0
SWQAKbF5SnWpG0mKSTdr1yMwfzCfXTHpWIWun4FmUBsUSUMHkMVh7VfRa6fdrNPAdC/FiarNbvFa
5dtMZEKzxRjIpp6U1gSyOFRDdHEZYaxmLxT88lSCSNuxrcD6sv7v5GSe3m7yShltZOfzJ07LJZR3
1iMWepnVCHUWkwO906PKPARp+J7RolVQZ9k9Dn0KxAOMI/mHYddaY0PbD6Q0lx1fap4mmnunfq6n
ncu9a2I8M2angIYKEX70o010cv4oYieCeNqIXdSgqk8iIakVzKaCRxcctQXPRPf5JB9FhhKshCwX
kCYdBOQX6kPGB/HaX/XJi7UOBPVlfH0tiaBBqmEN5Oz+cx68j/aXY9lv+Vqd6px8twkR+MB3F/UV
Pi9e9B26DJKAZxQoo17PfMRISrjauu0yXtixOA/LWuNoLaij/ftxJNmLr9hh7d0pv+8fmZ/RzY3x
kbhsH5cPDGCvid2kUrcD0rc3Dfb8fImLRmNBnTxJxVuurx7pwgchYrC8RVR9heuwS3i1Uw0hHvdM
c36dLEdeR2uT9OJQFAMSWnjnpOkvJRjaqdylMWJbeR34+NHMey9VcrqcPPFbSDudA6bJ9YaWHPqt
mqw+TWcDLrt+1Umks0DpAC6QJ5ZatCbck1xBRKWXrlcwrw3BcvCww95zhRbFDSoJ+apH3yK5KCOz
2PUNLlFZccr87sJKBzTIYfD65cPYAnsRN65dd3gQBFtzqB4efjgH82pITw9011s1SN8i0Wfzm0uq
TKpbrC0PcNdphqkPUN681Hgkxlps4RGEEWxzBCeoeiGoxx5g+pHHMRydbxsM6/gVFkV41X6wkQZW
vWUS6ipV0hDYnnyWLVHLgfFD8hGxbYpGFuXPPSxTYUnpXBTfVy6mOo6d39Mdxb8XHOQE5fNvgBJC
9oR/Jcso0Nkad/Sni/jLB0TIryl9XznyJcOpMz0ha/FtdrGixm6Ex2c5+8tX/Fwm+MZidfTajP9R
uWq1AGMGfG3trkfEjkHaTyS+FPK1XFg1gmqOK3XqV3lYCVy54DRgUQqGD+a64GJJypApUAfMR9wG
Z42aon6QysQxyE2zd4LZLFnmT4UnDdBocUPBEox4TrwnK8Kteyo4agCvJgDd920XHDRPM4OtZkcB
7n1YiPJLU41o25osqbuO41RNU8sVy6Ei47krWx0vr9lryYISEVjElaDZ6ipUGmbVkpzWup20HWDF
4HLWfFMIe1r6c8ZFFWZGNvt0dE+twH90iqyr76vKWDaOWUYnQvCHh+xlxI2JTg1zoqOPqkMbuvPn
lonRgczB3HS/tq2c0TQrhbx6bEpm76jsxKG5doaSPLPU9D5gDaM9qXGM4LtJN7zc75hKKOh7qkbJ
eC8Hjs1epJ09s8vLvY+m0b2lVe1RkNkqm4fWeUytbKQR2P2m9/0K03RW3uGDYJYGqvOF7Eq2HOD5
uI8Ya4NXY7Rb+YP/GbOukknWRJwbchGVjqHpYfuA4zsTLHpYBUTdwDq9uobpr9qIMUTKAXVbVC0v
C6j1SZZEMmgyDWSo+X42juLOhRHryEcn7GuOb04SsVkD58kGJCjPb8LRSKLrk8zif6w1N3z8rIut
aChLe5IE71zcZb+draKjcMZjfHfeUohxgt/d9sbVdLl7KkkRB283KGd+wWaYgbsDksAW9a78nHWJ
ByfvGAsuMnrm5vSSsamF3uBzkA1kIgcRiRgZCucm8I5L+DyVBaKDi7IUMWzYUCTtLFxxqJtC3bWM
8S7mn6NF7TpucebNxkE8fOizpaEQTypSkcfmtk9o4GiDDkVStScM5KuyrbUl9pOdqKmMKsVg0gFS
cDL+81q8OUeYx0NVXhzlMNGJ0gsXY2G1KiI5WIh2mJqN+Fsxwy8f4TPaf5cDXe98dvKiZ6KoEDQw
zdc78BurXNxbwFW5bx5so+N9PcBm4QST75YjXMnItRbh40EujdLjqo9IOMmG1qhJQxN5M1iu/+ad
EDDeu4DmgqYnpFy4B+lcghHNPDNtamNy7eyY1X2W2VmX2oMn3QhrVeWpZPe1BtErDhhB3QDp/aUi
bUFdBwUFJYgXWEAP1owjhRW15en4ITgEiKyJgD4Uh4kNoGa8rzVa6iy8JnCkWlbMYz5DRMWjiD6e
qyQSQXRphSgcgbbKRDFka6YGuqgrZtcg6W6ezXDJWp+HG+XcN7XtUTJVhhNTfuO5lp8snN7TQymP
z3aAPTutVst5sso05nKSq+exRV7Fgtq614Qsvu1iRO6rqC2RQ0W8UXiNpD0yfLSEfsUOc1hTJMaA
tUJ+wNk8NNw5TVLSOgyPQeDakR8g4vhYVv0VO+r24r0S8oaeGpXmEKOrluu8mgy+w+WFbVXqMrs5
OelvidVNGh2wjPGyUPJdeFLBjmQIcOGlCpqSszLOACJYzncxBMPTMISdXGzhWgpnLLWHHm0F03p9
ika2XF0XIbJDHXrSQ52EbG3lmhX4qNDv039GlosGUukfsKfGlsTpAzpldIlNE88T4P9SkwNkVKRJ
vcuvKP5QgnSfn/0HvyvdWI9pWM2YX/TydyX6i8WWUaZeePAgKv1dadN6Lxzz0CJBs0n+2mD8Lpw6
sKwRziI0jk4evWpI7tta8iFPj8huJ8Dr+fEWe/ajRDfOeXm+iAS/Q8OxZzlYjZxRhfkNMJBwSAsi
ZeQjAkwjSlwdPA/dHyBQzXzl6ysdIGFbWEyFZr/2Rxvwil0fPSMeWFnVbVvrLHYAUb0hLPDHKuHe
dBp+z/w/dgtWMcbc5V+5SbvXuTbzWoaPLFTh3qHM/XlCdxR/nOiJGs2afjPu40mdw6mfVYxZMVCA
41sWpAihlzPnN128d+HlhugTTQAcIjm0uqvmEyRTfllAGBlygHLj9TCrEcM9NXvai2rF9uc/+/VT
f+T8BrHtXVXSLeU1DYYTvDaimgl5zx83BaVY+6b+MxuXy0AmI5AqSpQYXxfnWhYsP2niFGGtGEDS
6Bx5bHI3bPIGiMUdFAQif6+Q7A4rloEgCV3UwENYl54Ryet0bN2uoyZSzLKyQppxKo9K8r1J2Wu1
40ITUOgg0Wcj9iEoZvIJ98nuiIykQSjqWdRXYYO0rDtdnl6044dV04jlUDx3BA0tabT+pln2YqTK
rRcRmd1Gtd2Uy0bJfHczmf6fQVeDGAP+XvGWlbT9WKlkErP2pyEbO+V85XnGvClWwX6lzyKDEEEH
/S3OkiHkYblvdjtgGdHpaelV790qWUYcFLR+61DhyGCL3EcxMeXHYMLN3vOLsnlAkPH4SJAo8HDH
SuTi+awcI0mPyMUcDFwKYi1PQHmfQm4XqerTWIoeGN1Lqc+zQDoX7vTJ5QILkpSM0mzctG3G2Be6
tmc6gn4dLYaGqF7Zk35hUEY31WvXiCLWOwaTotIMBybNmQQJGLjlBtE5b74FJqeqpLxq087TMw4A
wmu2EgzXhdUGHCNiyICR1vKb8iSWim2ReLCLOXcHp54pVjCbhWtR7hkkFuDMchbFuQfxg9sFbObi
oPin2DrCzTD2YjT389BVuJUeXYcygZta6s2II3I819MP2E+qoR7zoJ9nzy6W0p3Aw2VaOyFqBlPu
2JSNzWafIS+pzyrD7TmRPfXkaPmQ61L20vTQVhq+YoV0FC3k5iHbzNhzUNf2LpSVrMLChMvWQ4Jx
nlBC77Fti6vcG+GsZlQ76ckUjF/QLy0wkpWL5KKs3R/Knil3q5b+9UzdoUWK5fe8fBkp17gpZS3r
CW/J9ABtBGwlTKAcaFvkYEPJU0TuM0k9w8q9cpKuuFePl9xBFMqGfwQv/dwpxszXcEF1g3Iv2BwC
dtz0GN7B6WraoxfXuadYOH5orhKn7O/S7VIjM3SkR8O61i5j5AcvzoLKudtqCMvZ9XS2GUkhwkUu
yl49FqxV80KrKjVu+jPLNBd0d1L/tvKoDEM+czcHjgcXbe6PkGZeppNbwsUyG/VLtxE1j6+7OjH+
ZPLP0r0wiyb+7NIFqqZGq2aqRQr+PnYEQQohk4oqtREyiP6OP2Oa0wMs4F0RWNVVIfiW9Oa+S5mr
7rGKWpmlm79i2eEZbpY4DiouxNExiY8I5zslaE13AfbgWbm6mdJICDvxD/8g34wMMbrS1rWzExye
YH0Rj7rs15iSAr9/EaAEXt9Ze2LocGQtmJsnXf7iL6C+KNJPN6X1FdWsk/ApCZypa0Lw74Giyzaa
R08YNe1M5BIET+pSCrH7ndEWDSP9iyZMosu7t8U9xfk9OHQmaIWe0s+s8iDYP0YGqipwFT1ITVg7
AdKoaoys3SNZKtwxlTHubzYQBWJl6sWlEHRn+jbDucrSi5SIN/hIZU7nI81gbesCtM1Thn8tgk3l
jFlkqE+1W4DdcJE99XJGS6JRrR394HCDCJfUltGArw6Lbl22vmnWizKwPlD5Tb5lMlXPov+NaOkn
zXs3GyqBlbggdAzkyoLySoFpvudp5hMK+6aNWX7/vcbh7vh2dgHCed7vBhdiJN33qk7nixcFarjs
x81W3EYB2rvXrf+RNQJ7peAbHT9WBb71NPEKjP8dPDSrKjUIczw/0tBI3DBIs0n4BvoCHQmSnqMr
++cNZr6nNqALRw1g5kdMnzN3LRtdJN+RkgiIvLj3ttnNymmxFOpz1/Iia1PrF+/tMZAWDH5/0kzK
BCCwSnIFxnM1qF0asefokxcFjpbgWqPOqxbGFe5tlj/RIOlQakuhTYfJTN14u1eA/rqa0N6w+yLe
nZsDw5wX/yz4cRgA2r1tNF8hAr7HO/QEw9xK6GoGkAFz/3qczScJxdI8quCtc8qfdqO56drreqpn
wkC0WY7/9iVLql0+xz0LE38bYQDLMfluQbcpKrKeWh9YoqxPzl/1UNtsGqzASZxE2I0QWBpGefM9
0HB7WHQCRSCsR5usEEXDBR2JQyNCzvaG3bgeYFn1Q2HUklzYXv4+6tPJKvL/AAd2GbISAVbPmRFy
WOoPv3h/78+KITXcnPonuC8miCUE+MgyuHvpKldFWLbpCySirlR7VQ4iUHQq5p8IbZzdZ+dAKGse
KNpQFeRXgajwMkkfTu1PAlFZdUYjPpsCnQBbixPdssw2DyBfVzkgC5E2v+iJAEfthFxz4Yp4b7R0
k/4U8oOTHzm8mg05nd4EaURRzeL0ON/l1aGAQyfMjBvQRnn3BFnff1ZxZyxwB2uPOK1WoUC4uIdz
pSUtB69CDMn9Ld+wTNheAPwCitGI9J3dzE42majpzGi96ZyUoMGzX8JK1e8VRRjbdH2DKd1s1Z14
bg7i7VQqfvCTK+zP02b8Ho7an5k7hoB/xumWHS9v3PnYuJVOxn/bUL2VUSdMzEC9O8ksSOJp0+Bf
PogFSx1V70V9Y3/cTyEZgVbowQvFQTBhPm1Z48PutSm5ilXB7xmuuucIi+BTS5rzMtXpyEP0a8F7
dOkEyRAR23VdMjP26V8ca85IL/B5A/mMy4KhLbDK/w1+69IWSxQ+XUt2HxYVU0iDSxyoqvFYIODU
9RTrPsPuSCwn/7pp8A8DJpHdVpdDNyuviQNsI/kZDR30QEwpdOPTfRV/7NAcAsAOkN5ZpQYfKSRD
7W6WgfYPbeQtqa6FDvK3G8kpDQeCMAHMAeaJGefbe5wp13OFBMpzpo1ELKj0x2SCpkrRf+3dewRP
bCZ1jcKYOat4NiHCqVRIyivYzj4K5uLP++yWYtUwMTiY5JCLuyaXD4G1vHL/Pn5Yiq3f+3+68U1j
Vp/pjkiKw2EBbli1W2T4L98gG34SUbDrrh7xSMLTpvvGSIrpbsH1y0hw5kjZK+Sl9WJGkuoX0q+W
Rj+xydP3YzFIfIuJGiKd2dqVNfK3l13P0/N5Sl68Z3XpTgVMITI1CH/wW40PlkJOTA7yk7bfSdZy
AmGCyd7mMjz7wZDP+WsbujsORLlpGzdAsXUYl8eY+T8nXjomHqknz2RRq5VIB0b6wRJGMBG4bXi0
e/t9Cy3+VzwHGDDgHT8y5wHA4iCxd5g79uLy54feVQLvWSt9uQrSDsF/tqxP1Md3D5l0IpLtVtYZ
cFGcm9B42wk+CzyJU4SlspE1aGnA34vULySZIw3RTbAz8E+wzptfOeZas8ukH9/uk/XvTRIRZM6w
JAatf6M8EUshp4r2mjztbr3o8Y98wpKFrEd5wFu7Aq3W3oDvvnNwFUTBIgjoe9owxbhLemvRCa5Z
M/BUpqyB4OCujarHFk4AvimDnTlwrC9fDBETWjm3k4CoB9UkUOAWWokPBOnlALc61n86aRGv3ER8
7KbeN+dJ9VXzAniD5c/a+JYiXvWYTnP93YVa1q7l3EhYnn5KlKX38eMlvCtcw78Sz3iJWJQE6wFd
VSk0fsdF86C9czEUPSFFcGE0q7hhWW6g8IH8jwppTqL1iMFvjZRN2qbwt0J2xXwCy/Dr+tWuveNQ
LP+FNiOy5qZSyQjL+Vfz6KxEBmwLJPQ4sDqHmE1BY9sFtcMRK4p+b+hrCu5m/kAeK8TCjUAggHmN
VfWz2wxZ9n4mkYPFACYuZbzIrrB8OrQMl2ITnhjlcv55jeS00wuEkWyTFs9ck6SIblj9LgZstpaC
n5Tlmv0dN93q83DP+y6AwNyLgMGcmpKPRP3AwvDtPYcLwX/IV8jcqZ+h6ySuTvyS4oV3Ttd0GVxM
hLOiynZ/0jpY6ei+rVhnj/kG8775KfedZyy027cHQOE4sRaFEyNRpn38XAtBdkLkrCOridrmrWMV
E5NDFGhIswtI/+T6lNSt21sx66FWiwhG5Ku8zM/DIzXXhe8ZoBi+DTyoKfZ2Fxy0Cy4rA+RuDTVK
llNe3nBQt07p7TTiTNDln99uA85fqVqBflnr2aKKQ/xeOqJjjhJCDyLt8uwHjS7Sh8nfPLgqAvGi
Zox6VYKK6nI4VmJ1pT3XUE84o56zVJwwRL8LBBJnTB9/YW7Bdr+oGBLL0mkrmRiATS0vQAosBB7l
ezz4WuHmGbNh0EIBYE9bdVX58br0Mfn4lHyGG0JDLVz4sAUeLv5tKDihCY6J6fgXVIIR5V+pnPZn
WmESy5w0CmltkLFKj4GD91x2GSnp7i3jgRmKlVxECZcWjj0uxcc10EpQYIcqDo+ASEcW7P5Gbm7R
S1Q5HVH2KWQ89yvc5iJCSAte3teTYDgtw1Q6nb2CQj7cf4LDxyEUgUA3uVHrkQpi4fjWU9tlHOMN
UbSwTc0j63xhvfDt4yjCRDF5lFzPKHGNGwNEBLPDO91nOW3J8Dv2XA9IM/OUtPII+RhEYUQRw1eS
24WAOGTlKF+2nJbfZMfDsiP9T1B3LaiDFSBNCuw7RJcO5LjiT4yDU/R6hvxaDJIRPbuOKey/R0nA
PUKA7oqz/vvZGLFnZKMFsLtHICy/StRR4um86U/PNfaw1YEi4kH3W0vWap6plvmJFQ5/aCZfIffp
CrkcyrkBlkF96hrQJKT+Q1OJ4pH8D0zit1M4epqGKAGRj323Xv1RezuctRZ+Y54pJMpUDhKNZD0j
eggb2ScozcKQMn3uRCeFC6w49QfgEnt7vS663Y29WLjRoPcBJhfBVZL7SUk1NTeoa1vBwWZP6G0w
GeZH0cfrPGsamjgKucJlMnMyxnU/mp7s5LJOGiaxWWbkhYR1fS4cqvtt9LbHuo0lSeMManWLVDdP
qilLBEZZNKj5mr04Bd9b7SuyYem17bl2ebuM/EkUtmQpN0vqc3Z4m6PBKRAdCupN3RxSO4c4XZeg
mY+PzgjM2fEE8jlRA5XgDYwQIOS+mkzUUcGHa/9JJEmyNvtWiaMqCuYSZHLEODfnb6irHnvubHEM
fl4uSS2MUTR/vGNEJkUJskpRkIQxIqIosnXjFUntiT0Pqx/sriE24KKSfDdX+TdWb4lhR617hYkZ
adAjpPc3e/6lGlRMhllOYcjowmuZI8q+/rN/s0ImS0GDrX8gxkhW3n9n6D3Nr9RI5zfnVWEs9SDw
NltuI5h+UhqKv6wAuRdT5e3wVd/CvJoLqxq6OwsSbyhZTN3zuBvgUz2WX1uhyX7iJaPuH/2Xb5ne
wkgtGF0JNw1OB7+rcKhn0eXgMUtOSlTaSwZrHMMxH956LMbzuhq7+1qlb0RlqijNO9nUKFVCpmmw
ikVB360AbKVg+f4HDK5WwfK+XneGLajSXXSI4LrxfWPheTlpDZRFuh0FOzu2wOGVMhvnoHyYp+oA
ZzKZ66vR69Xj09+4svTuSSZADl0f4yyeewxE9qiCTys9w/DD2S+AA5r+mhlbtxBBGkbw4jimFXdA
J/T6fEnNnpyU+hSMH3PL/gNK/BlNTFA7xfin7m+8VlNQcjk4GwucH2v/hDXoLtyRs8/C83Ul7iZO
C5dmfyQWjYW8fCBAbQ1FICNBdQt5wbV85YAv2XY+GiKykBfAP/A00ihWC7Ul1kYqOnHczkjhl1/H
g6YTFz60zXPJZ4q1aX9misvPL2IsimhF16ElxkTtHv3LxigzD/ZnlbYba+gHBqcyGISk6/xEtwdx
plGOUdQ0s8zMOYECUHyTMrPJ0tm2fPMfmaBHLbC7Z63e4BuOPXLfFHoyQdfTTI6NAODdrN/shiBu
OwiWq4i5KLJbzOyXFBqWtgiMWBrtwnw0hFtkkhz8p1iQDZ9Obbq5bLd/gqnoIkLdvPMVH+1z/y83
MObFGev9tTXhxZNIntcBaPtg6XnD3rKvRsbPATFt4mui7plGP5jFktbUOa+pol0ad6+brsyL1n5H
bFAcZpK58cyjkpPHuEfy0ZGk6Yr8mzh/k282EZVlfgPStxhPOKsmsAtC6LsFShuJ/U71IUA3vdX/
zZ1FG3AUfeb2ZjX2WptheB6/oCVVKFkDX4TigvlHcXAtHmV0mJdg0xKB3+9i9JXHpIENbtlgxsNM
vhN+EJ1IPOOnEsjX4Kqvg+do8BiHYOR9/jPHONXg4pHOAZWpK3an2LLkehiqvDxk+nVAJXExoOk1
MdDRhJ5uLbq5hQM98e113NcTNFly+3z4DsWbj0PHOLuiZ/COy5vidEiczWqycMxVAVGRnTDl9ZL3
plsQM59/GOU5XT3CiKiTliHDF9ia94SYuN/+n3vmuT9WRVvPLv4z0IXJSHCagO4IZaX2xoKwDa1Q
4S0GD0KvJeKMm0SOSEYxLq1cBQMvKs+u/59Ptlo7tAZswASNqbD0yBFJQr90eALjYHItbNEswjri
vNpkv3/OndAF1jTy47avOZf/dDozyKbY+7+nzs9KVSQcA9xj9TkSu5i4VRzMd04G858QFuZG9+Z2
fr/y3VcDoIcz6wLeAFuTrkW2iKOsM0W/AQIw20Ylz72fYyi3O9cW6xl8DdxMsGUx12y6/kqJ5muP
+v4MyGAvqMqzaUuqHV+lBrKNDxBmItbw8bfatZrJliamzV9mnbFU3qHuIJb+FXyhfZZXLuwsZhk5
1bLb9tFar4vxvQ0rle3yrQouYBSEhuaV6T6Z3XwKlqG9jU7dFpFjOyd2f+GJVc9JmKGnY+h3xqEs
zZ9DA5Hv5CQ7+oqI7+jLT4PbxWQRsz3OhQ9Jzq+iaQ+b/eAAF8rQNTb7Lej6d1Wt/0tUC+fmEE9D
BjlZzDJLUDT1ze03fsnHsdc1zI5FsJAjwIvRxHSwL1mOvefdWxx6aE4lRNQGHHvpMIGXUkVDVxaa
bQccfHh8DMjtEFWkmN4Eu1WscLvNGIQx2ysdkWU/SFDRQDzeKDWGlA/OWx5j3L8xtvHF7Ty5FU+A
qhj2WfXtMtJTHyVh/AVs8Mnu1hK0KXhXqrpETduFF7tBXjTc3Q5s414tsEMfUv3MzS1MW6GyydGo
G7wpcfRze90DxW3BmghtY7wINkryXVRh/ubjigR+R/bIYQHv7CrNdATi6wvFNUWRM9bikogH7b5y
8JuGm1F3lJKJn5t8nudn/3iKE6iAK+F0IY9k2l2kLYU+qMbiGhHWFmbK/0vnZRtbkBZk9wj7faAs
wh0AughtBU0VOT8ko/kYV4W/FcGja2Imechn3vlh+lN4adYXBOlLkVKBbMq4oOgV5Dtsrc65mxQ3
XxSkdJ+Io8dWmhRGxBtfWZS10H3PA9PHNNsoUQ30AKT1r7xPemEaHykgQylqH+glHMa/DyXzGQvW
efhr2GNeAgVS5972qzQ7VmBKjsqDx7im1ABp7XQHQC0M+RBpeV18ApAd4vbjNdPMSmungfjDWG2A
yxk4hgGYo2Ytl/JslEase4jvdD/+RYxyu12R/msmkH56HD2jB6tI7X5SaqpOZWW+bm8veN+oNdKv
ZxbctkY9fajm9SgMQA6IDajVFBY1Z3niqfoQpX1a+hS62n2zZ39uv4SlxdWGp0GpCvyV6tJQOgr3
1+F/7Aa6rADGthg+XSbvVAV5bF0NrkJMz/t50j31M5SD4O+Elx0UPYt53KBUIRmS2JpjIK5Tng/N
UmofErk2o+Wj5qjXbkUhXuNzesQ3nYuxAwRIBIHoL/d0JDRBwCpOxIlL2RJ9tGPAs8lSSbb3JE5f
w5PYtAtyJojRD3EJW7viZ+yM/jOjPz2ijV4DmV0OXH2XhS06DNRgamQeI68sOM94CM1jjVqWxVQU
OHjN96TQbaDrQuZOEDx8t1bN/rc9gILAh0heH0xbgu+3Y45xR0xCWBa1Qp0YKiz0imSMDzbOvKuK
bYGWV4nG/pEwTq13IcxWEhXXtUluqSlifYOnqiIWq3FCvuZl0M2vt4DcBried0ePHXPEvnOh/3je
MIjV1LqfnAZtklEYHzDBhkdF7E9v+lyRe8Dv69OBrI3vCkfrqGGeX0zNuY7oHPb50W3nOYp5HYSd
QpHJtVOJrnNu7rCLAR5yhbQSgRQQvPIwKwAWMIqEaqZ706AXbPS3RdujNs3ZS7aYgWWwKxxIWybu
i1DQb5Hrr60hoceS8dUA5CwIRNaxyFqfxM9ibA4oT/W3RSnbrAUzN0ZzU/IKs7VG+xv840wDeO3h
TVuPaFzuFYh3wBfOk2T8E+66mDZsBtzdK1rcYBGbxZF7hw+QGAClM5uwvkRoN5DWT3zwDkc4tqPK
NkJFqwGfZP8TKwGdtXzLDi9XOkrJa0z9RO/T6Z/xNKah4aL1o5y5++f1IcD3M08rS7u7rwTYVjvT
5jfEhzAflOyXtIKgJSVJ7zJq6FVpvTkBoIirbszTO4XoeVRGfVK0DN0cbe/+zodpghNu2OC1FdIR
92tNut/bIIn0m+2rQwK8rDc2a6VRD24BqJIiM/mGTvGuIjKwDHhyU44wmc7GkiCGQshDuJhvBoqO
crP1teyEpPpDFaD5bKXDglE2XmLvVkbf3wtBAWj+IfA/mSXyHP6G+TscJO5Wb8mXNnQgT9TraAq2
915mI5c6W7HoYEcgftBlmFuK+pz75pKoZiMQ4u3w6A4A+HNfU36S3v4LyPpjMe9e8pWNd+SJnahN
4YM6hZD4jlxCx1EFiw+2uUfE2SwseSQ60leG1Wdo4sNkPQ3dSKzKWH4mHMe1uspDvrXHKQarv/sC
d7xWURTohK+UZBav3QWUH1/L9AcuHmlVzJo0ME5kjYEmqmPMgU8ZmXpolPyMs71kfQSC32gqMG+/
BnIlCzdjWBMpqHmH0KOHi7SvRT54c2dh0iCfxX1lyjIHWzg4r9Xg0Stvzm6YC4++P0BnJy3ibvai
t0D4a2GT2A4eR07FG5ggG0M+TvnZCQzGqgTst2Wtn1X93Q8Wv4jBS/J1DMRq8i7RoihgZlGLGtEj
MDXVygzBQlNkmz6okRN+LGc7TkVk8ngf+Mndb0kN4Vbq2aFEPM17BccXtWqUTqz0nN1whvlUP0c0
ck8CRAr67zn+s8a0prokL9tuapKKXRVOAfZMFdGYBCxYu0aAAhs1HEQGcFM8JRP4SaYjp17ec4MG
aYJm6a5T7fh3aYFCjaAuxpxiylNpKHNeCydjcDQFzty3oSQgFYlMXwlx1pRmCmgNwLWclNlKQaG/
HsZVG+pNUZxKWauoVHeb/cUbPnfIYGXKKW+Q3At2wGadEz2QwSriGpUAkAhirFh2Sm7XJSP5/3eu
k2jMkOBK2n1QVj2/p2Nr5A303ZK0SYLDdienl3rrfaotzUqq4pZPMoQpaUsdgpdrP9uwB2Pye63/
cl3n/14dcuz3Y3SPBApGSW3ZRRXOg9ic8VwFwLbdSqMwiX62WEnb00kR24mHaPCvmWnrkXUOQ/tI
Ylo5n9BXm9yHLBLGN7iC5l4bOJd4Rwz15fN0fhGloLuN6ZrJQcd5YMACcg24xgh7pYtyxTDdhmW1
wq8WtckJRE23FSHEioFXkECkCWlj5uM7iudG9vugexSmC3EVZuCiI3QfbcWiLtYtaA2EOw+jVpEy
G7RJ2xNYEk0gzCr47yB3G1wLqxD42IYE7eAi4RYLzVZdBMdhnbLagtWMyVtSdj7FJl+gubQ1auV8
BOYuEShqgN6OIE9Z3L+M5/iB5wza6tnUZf09hEuZIN5tfTC30xKaKV/Xi/7afNNx2h5W/GwconTh
VazR2mVIJNyQ5AAeI3knrtPYYnzddXLD5TIE2zshPzCHDKFdev+PncVDZzGjeN4jEs0xrF/jxRoA
HKPmdVZSFxx0l5dvtR/k/SUsanTMbrAOFXBjKtz3LW7AtcfmSvjYzhTvVBdFzZCM4gwsiOabSAsG
MnAoxj+8iCsyuxeKLwa+jc/1pib0CC25VScp0IqsqM7PJml1bLhD0YCkVCDuySvHgmZRibXL1DBZ
xy4Jhluf7ocT5WyMqMSRs5v8HiRttppg7u0RfSFY0+HWBS5kqVkXvxrKRb3eMxQjfBQTGaC3BJqj
ljUZU9+/uabb4u7s70KPloLFjT+tNQddiYsEK3iA3aeun5piYI4MkfOzapZw/E/lEnvKAToNMndl
R+8L3GgR44Jg73Z0916MB02hiQ/a5Np/9ouQ/q6+lh82Yboi6FWTHMw0ls8eh756+fcd/xuZe7kp
6BdBsWcRcHbfoPsoeQFe+AnwOqpCq9/FDugVedEUdLrgDzpSrXdHMC81SffF+UqSmBplxC+n7bqT
LcUh7/3Z0vwLk5k6mmtkrLylaZxLyFkmUX9wZW7Yzc7LA3uOnJk8IwSBUkNsq3kGmQQ0RGICSuuo
E8tXQtHB18EBsVGCGy8s0F9lKBWSHdgRDkWZJayNgQxyfrstu6z7BVQmzUZmmxjyFtwxGZHYG1Y/
mMEVIlBDJ38dxgv2vr0ccoRF3TYBaA/N0KQkhWMqaehZdrVMnyICxFlfPrlKjOT1F+1JdG0vhtJ+
u9Vx58Hxb5w0i9rONLgkJ06c2je5Ikgsf63Mij9JbTihjRsbNGLTr1rQm7jSyykWHT7l1j4Mb+cj
M+fny0YScjVV8yNxgR8q2Pf6hRznqqosVmitm2Cq8ZakF1mAAm3XZLHX9PloZMumwRYYxoLfsYWr
aCj4Vq805aZxCtx75sbxcz2QsS1BbTTaH/+UlW7IEgY1ft28wQrSKdypx0ZIhVTaXgUHVzz07ONv
h1gpVltiYULGBkl/ffEY43KOis6QlvHdyPVJUR/p3Mm0NvE2sUWWKiV8m+CVjIi2mNci3pxehp4C
HOw18+XAfMcjmCNETS+GPsbZA+1SxE3mqCnafR/1daCFoBlvrU1jHw9PpNGnc4mAYXrg/maY4POm
y3X1hNGz8lRCDUCOotf2vo4SqntWsIPuujRKFPjn/Lm1tsbfKs/3YOvMdHk97PURURvO05GzlQu4
Vecl/j+9guqgwa5NCO8hfH8FqvwSscO171Er1aQFxfM21sy72UmKGMfl81PUxmxRqoLQvMrskGC2
y0XjP9n1AN7/gE8TmdRbJsY8gmfjb4I8mDGVIyQIB5djDzw0JRUuV7AM2NIZHO1SOf2hImr786od
sATmxk6RoCXDYaCKzZlIlL/nSwLneSCxQFzzFCkF3RL21yNaHA7YY18teeNB/vp6R51Qj4ZR5lAF
Nw8xWekziKHBzFInGnOaRzlaeCWOXRe3HgJqhH2ORpQ1s8fJuNfnZJoRfW5F+mozjzcWZU3uWmCZ
SF1aJylbOHLFvI59UygUbkTgsMpUi0zjUnhMYEUiSMp1T1OnUiSGdFsTRXHkmRaIgdYUYP+8BM1o
YOTwsDWaA2e7ZtvYa5CR7+wjtrNBRYe+xOLRLZmY6SganYRY83SOYscvNN/BAjictPh9/p68TxtJ
pgWbCUg0mHBPYC0EWgVHkQVHo1hwHdt4WaTLzM+k0vwGQH/vOndmndquTJFR9YgkXZjpc59ZWufv
+4/FMXACJgFRClORqhkKJqAg7HQONIJJLHmNFdNN8Nh3qY5YlDMYLsUL6YFlGv3rzGOjSLs37i8R
FfQ0SB0ieys/4WnTlUQY1w2zNFjxGdUApe25BLPjZEX0ULffD4RO3NO409AtiYrca4Swm7eZXqmR
sf70wilrrxDWx413vgNk+4fkkd2CIxMANNzPkUCjZFyOAvY23LR81RkhAcwCeh4jU+RuVVshGP4/
IS9UOl5hsWbuy/KpWX9vKD8J/6g1FBsUUypnQL/j7ifpy3GjwiSVT/9G1BrCxs1EtY9It8QPYkgm
OQwxB9vHGF7US3tvWWwXGI5FS5p3eOXzBEdJHX1TyOb5M+qNOjulm0vlJ7kpctl+9oC3X1qQB9Ok
cdKDh1+qbDUsmYt41xnbKv9sTsfhUGzj6MRHHsAEuTNlCspk5FfsT2EvWb0K6KLyW33sGs9Az8rf
MyTdwOlFfBm4/dIw/Z6CkAijGoi277mwwHCpHjSCTrxE2bHbbbn0kuf3/A8bMGiuH+zwL78oV+gi
qXMG6sRXEBqFCbvYIXxomwAe5S9/5Z3QQH8QRwcWCtKtEAnuJpYa4xOWemiLXU4qpqBKsJ0PiAoT
fN4jL14X8RrhxGOPlYbLhrqPe55wLab5uV7UZk24HMYHPE/d5iD7Lj5bkEZfrnokcKtIkq78wrNi
QrrdXJv24KK6QlvMwB4ZLgYs6+ed/OtL0bYyjkzZZqiVxRLY1gkeQGKQMoGaqaMBAIAlqThuVKKF
XYFOB+5ic19WhMMG1Z28ppvM3JloLBnNgQEpZnO26ogSf+UvJSY3XqAVTU6mGvQ52kXQ7uJim7e0
R75FRx44hU9USWp63ebLvSYFDiMEfiwRo0ueziW87cxNRcGa9zxlsQzxmgxsSRTrwivu11DdIXWW
+1zQEFGhmhfeTYutTj6eHZXngXGf+DKf7j/2ML9kjNHqvWfwNnLx3DOK7gztEKPl4Q+jTxW1RQEl
CWtJMb2IsOOOtMHf6EebhYi6thasR2/TZclfNf2ezDRYhoSFKZ4hVNzlamlwzlPptzi6cnwi9tgO
cGAdgVP1umoFgIoy31HrArLmgIyUPilV/6rTQOvoMJ0BNQV+9pF/X28XxMBxxowNz6H1kglT39JL
ZhguxniMD6JzuzKVN7ysO7E6Up2JfzhyvOrsojHQMke/iDFU9MBHO1TZxqeRJiZfEcRFYC2DxPsY
aVIPAGZtxEbIWdeDA43zp2YhVxAB7qp9WqX/CWmUgZaQFuMGV21qt3YdWOMwIertapNxhzY2z4FY
fUr2Kkat3UXRyfNZutypRfInpHOJfl1rHiPD77ce3YR2CQY4wWDbZC2D68xjHwTsleSZUtIrRqZS
hAnKgsRpHaBABOgCxe7IIODxOXt2FvwpnFBPVqrjhw5wGXiIFY+REw1ni/purdMpn2HJs9jjiwQR
xucVJ+sUDPIIazk3nW+vCC9ssPnTu22F7enql98JmG5+QlS0nrMYRgKM0nG65+Q0wdGJXtjbNg4g
OuIyZgmICUfm3r2WJbaCTOpGBDj1uI8u3JMi/YIpAhqGViy24ukoS4HbAHOeZ814tQM3GrgsS1b9
tHuLt/+LRjeeZzqAUf/lASQvrvkjr59SLN8bo48EiNQIRd/16crPfsLMiV3FeqAhFrDx3lIUvaGi
ygoJDIT8v363GLrX2z+elWPh4LFyFRXRzjp9O50D+brEw9r1zB/vlcXJ5tXJOMKX/o2wQn3kqB57
mUn3AbQplI7MHH/GZm1MSpvYptUPZb4KCsPYvt2pCqzzH6/R+bHTzMclm77AuRvyINqMXTwayasX
RtmmDw2LkouVKihP0fVdpZiW7D7aS8ZMvn6MaiBC6+N9SNZnpFpwRLFx99pII0cThCgoc/0/YmTE
/aih+9Uw8ZFwqTJBaGKsU58RsykL/xtH57loIcnxcvtxlpKGtFEfO7Fa3CZBseNvL5QLZeX/7kHv
W7/ItQIN7WVxARgnQes3To1wgp9F58nkzc3fnpxDBB8y4TUE82h2U4nGkPQo30rQMkYmwssarJoH
FKPMrfvZfI0IFB0MXVKeMDHclp0825Gavdgg+8Ni+B2ePuWO665gBgN36ovIIt6Vdqq73DLx4hAL
1Ly1zaXBCCsHsJ4kZ6q/IzIdosAQFWNeC0RnRjw+CogeEkWd4pwwd2YNp4qdsLDKeCuVjZ6oVUmg
tL5XCRbxo8l+NHKqfWvNArcSHxT0ho7htPrsOn3gc0NE9+rRJ0BqOf7SRIGss6wXUHYhFvN6s3TG
DLN9UfZprLTxY2J9BGXZkO5qBNzhMlQsprHRb9I9Tqowu/jEB52F4CW2BkTiwThgZVaBYppkZ9Bl
0D7rp+VI89B5gDP5qenybqOiKmPNXQcu9Hk0OE1W5zvI14eXDhW1mQz2MqAIdcfd9yG1Cq+TafLc
/vglS86F9oKnrQ0rdNMmSFRQFtMcYFpub7YHSeVzYNMZMFI2G/Lz2aEGf0hgM2+mDRK3OaQ7j1Od
qFo/odasiZx4HOSl3ij3zOfOnaWV6ydgieSDfCb/HCENr2apmMFFyAKp30kawEBLRrtH5L2JyVBz
6u8599NJ0m+Wt5vqcROp46xu+wAd7G1ASktaByE1wQEQa1wZVicOxAshnVwPopm1FXjn28O2lg0E
va7BEymTRuov+UWKbBBiYvFPHC1mbTBbYhIwNOYnvK32+jQN1YvRsGdQalnFc6gpjRCGSoV26FVY
L4q2hkFqeXl+XZFWuG2mdpQ26caeTjc2+ZcrT+aA0/vK+QxD/Un8ju7v8qlybeZnCKE4Xp0fjL0g
oSXbJDEhGw5pyqve5XsmEoEU/QpZq0SANvfPztlUTpYdBQAx/uxkP11ZqVUKV7ojOQHo9S1QKZJh
ybahdlzyuUSg1s+x3ZDpvimS5M0wKUbx97cxi3LB1lBU7hOMDWBrsFAUF4rxykQ1BMsuajk56qFo
PMQt8AaYxBj9Tvd5jHEr4wd3/mjt3o5F0M8aDSXxiB1I6vzaSWa5T04/hqq6km1Xo+UuD+YLFJ4V
2veXn255DPTReuwg7NM+QyzzN+c2ZzC/QJX/PukkhuoxC5UGDPZ/YPx5x35p5oKHNhMLfY4vQwUO
RRexmEf2N+dKDC4EJfEMO75h7qSr1fyEXSEsJN9jAm6v1/7xqHHjs6j4ORXkLU/UamIV6a2dX3+W
/774I4puiu8ArKrNJ1pduEDaJW8fuEdUaX9ctDUZnWDLVaVoiY0JbYTDWvxrWmJrnx858o3TVhmd
axpnQQDO313cOqa4jK/u51FnxUqRyu5oStLLCwf+sMYJ4TPKW7Imm5eSFDKEEgc1BxqIrLPPutp7
kagRjM6ASS1m2kLItyXjKSgLxS9118evY902EgWvahPwQ06q0bwxS/NyvjWFHg+4TPn6/ngCuZtl
SOTes15Kr+GQ9WPKOMMI4bBaN5KkTAhDKOgY1jzXmXfidA2GVoPTHEg1IsG6J51eFkbQK5bmMrMM
udNX9Hp8VHUIWpXCtw+EPhkGQjWwJOfKaHNXuXNwXe4Hb8I4WdBbvmTl/7FLVg1bcaNQAcDwWhYe
HmAvvKcLpr6URrzj24NiRSJ8z6bMxsRCQ4fBSu+g+iasXL2hJLjc8ADLNtau3XWEchMnw+FhqNtS
SezRchddYu4zUjrb5wbm3PNqy8zgzwhfru6Q0Jaw32aEoZ8mlIqFfENnPOktYpoi6MR+3zdZSyUr
p4QsJoSwBbk6iVkhvUAeMKaBIE9E5OFy9XzT0kQushYwfTIKahkwvZAssjVQIOiElT892hdwkeQA
Ce7zd6tsVl5hHwC+DqmjNlFUeXoU6PjRwT+NdRmN8w7njXm6sQLd3+XlnAkg1bc8ExKqtszkISuS
h/uSZzWaKZc0kcjMy35tEGpGlZVSTAPk+bN/6t3h7fEaat79YdfkRTilEFH4WJrsdXrNA0NWJBR3
DhHw9hoayVTuad6hFqhYwa30ukbCVdBorRLNhPe4hxDOdAIoxeYk1r91otnn/HUrY39gcX0i0lTc
mvMrvvlSDY+f9UaaUjIX85RGHoL+03L4YuNlH7vXIegMLSyI929uM+gHO1hx6HXdO9FqS+RjGBGR
b22YwB0K3oPM8IwJ8PgnoopojmNoajExIOekKehzAMO9f0fJt6qbyf6ZeQhBEQT3F+VlTdcJ2uUl
q00pfY91KtudRC8JDyZN1goLmhJoFjOslYU8TCN8KiDSY1a/ZqNNTnREGzkXVa54RKG0lfTABarU
FLyk48xUkFXGsC0vCI1evu86HXbWtGspN0bkzzERfvR17FSv/b8cUl4W7Gbk51vogMz1ETxt0wG8
M8ummtJdTxyM+oaeJBFJ7MnbDk2GJSIv8IbZpt9q01QhvRiM0QWnfRymDhElCgCR6NvGz9VnX60L
8asbxKMCYOlI93sPdvbNcvUVntQCWuNJWDQnVHDa30Qmh3Dq+g6PqXxJXh5+ZwmlslemajnlhqdC
fsWP6myInW2S5jP5KhZOACOugbNmPPHUa/HRpRgXSW+1fLZjHN5g60fylwe8HE9aJuaufTEYabQX
nqjCnfb3jZ7jdOEJ+PBlYXMfSR62tQo8JvDVzA2RNIKs5s+BBAaq+wcWVcoIoKnlicge4lABUh/f
+qkUKVX1TUIcB6o8F+d3U4TWTM1zU7eiQS/5XuDkNWaLROVLnPZ6wn+N5tsowdcaIEQautkK6SfD
lyr7d1wLWFUMxHlKT4OxzsGFIFJh7jc2ofFNDtJ0lSsmZy08Y03FWJVKPJ8zyRieX5imNpRLsrFx
l5pNXySw7Wu05JFGacqqhr99XkWNMD1LkU1lVW3boy/32ZcolOqs/rfs+4auY7HFdfQXitlNfith
ThAo+x5ac1LUA10hMr1aeWEX5zFbqVX9JNXeVgiKkAnlMVVx3iqE1iMm47aW9P/HBhv+5yaoegK/
4/ofH+Fk7QyLyDe3M26cU2VeiuFsZxvHwXZaajiuDW+crt4vU+pHN5GdVW20rYo32+277oOZA86X
V1gnw/f3RsQgI2ZJwB6CyY25r/K0pOuNksxmrLL3JjcQaCfzZ1aH/8Os9u5j+TTtbY8zKfU0nfG/
vTevP/efN+8B8S6zRgu1DkYy0SM+H87CRsNs4pzij4ANlemMsp7w63pblKTaPK0JnJ78rNBIPHXZ
Jq3bz7HQFSVOqurYNyug2W+cxDtwK6qNeHbi0qqA9Ng1YlpsQ1kCIDB3N3Q85fTWsExKWyfkoTNg
R1ZdrKjvVmbe8LFbYRU1iRCf1brVjR49QcPhkfj/uuEdDpLJtD4wC1d50sJCA0iTTwnzmvpowjRy
veQiWaX+AtkpBVS1L3JO/sWDbNlkYJ6F1cGU4Qo4rALNPm2RIUnkcStd5WDzC+rvja7Mshd88kJx
R5iYeBoM7/HS6N03tXU1a6ExGUZL/ta2VqPJ+Qj+r++a+k+f2f6SCLqkCqEnwgYvtuEBDQT1ixEB
3+zNebbaGWORj+7PNOSr9PEx8wNnM13fwvyu0h5ANBraBXs4LTGgOe+tWqRFsiZrXGUuAXqyTYYE
UL9Ji75ZQ+Y1XpN3QMizdaVl8DxqeLCx5EcsvR1muiSTP2xvHN5oghrNuRyEZ13KHLBq4jlFd8Vz
+W8oloNJatp0OF1bNbTK0/FiCBXFgixUzg5fg4hDnbgbHN6U/AAFbo02qkat44g2ya6SYraGCKH2
AOHWcEjIiAgotXJGcVtd+l62Gk/9va1Lja82gb+WhBz/uFbLfDjiihoMdmpfEMzqlPo+foBipdyO
0QRWVenL+/Z8JB5tCzqdIJ3DPFyzLTBYhug97a+PlfpJt/33MAeqQwSPhQ7N7vJaQmHJGp+7T6Ii
tJnSpKCE8hzrGj3P5ki3d4eu4SXU3xgB1vrgKwHbai8o5wWcZyuLV6fonQ9mFemZ9rI3p+potjpb
dR+q9wYNNSgcGvB0V0BlHsETS4Qu8OxQsPmdTqPOfHoBMTjESIgSHoqmTQrp7m2/ToMx7pr6KQkU
ubJk6oo3Dm5GrAdYI9GDJljaAGeAH1Ppg2k16vkeBjxZnOt3R+pGeJTRhGinBtb4185Qq4KNcskq
DcOSd6q0Jx5mmjdDad50Lm+bLJkQQq9YdjATtuJsWRPVV4mo/0UNlEexFj5PNwsOCSikfoGh4piJ
7Ppc7cCvSYDx0Kef2njZQsWjwXQEWuy9otoqgzmuK2X7kCsb91vvVG3mFaRCJaaaB6pymrE9bkVo
7Z9PulNc36JH6seqo6DtUadFGG3jqkD9Ihkc1HR3LosC532l3XEXvRsguaS/fWrYwndBSj3lo8Xb
H/xiLO2U1wbY0QmNLEKzSJIsxcU5ur0HEZy4Mmbt/A80cFcJiIMLL3wNBoY5/7/byEFpQf4XoEth
Y9+1yiNpDuFw+myrWlWBbqouukI6b2YasEA5SN9uXVuQUd9ulnSb6bt6r/c1U9WbnbA4X7hvD+AF
xjiV5flHN5HAQRrppXSE88UYBjxKaxrXYYPFWI7OBl/D+OPlig31PjzpxCyJrK1i1CYj/vE2J2Y+
2uheTawUsKemfNydq3zLY8AumryM9SyA+ZezDX7125khyTWcJAObL+9c+QcTtLfYBnN9oR0K0ptB
1ng8bzId5Ep9GLffbKXlpLJ1zOl50u6wUgFEimgBQjO0MhPYYpnPqSQKNwXHjVOOl1usRem/eQR+
aL3GC7TGSmV7zPvhbc3XdYrmghQkMmoBRpFqzUoZ3GKR8zMuaPquSVhLoszW5MdL2UKaCNygrYXb
xnTavbzWTBRN7ph4iazSoa/y20k+TF5EE2xN18jBtfSe3Fk5+rcf28L96bjeU+0u4a9NPOi40M7+
jxb98L3eu6A3HlhoPahS43ROki7gDioLueFrmwByTf2vA/rklNAJ6YrzfZxl/fDr8AFH0w13ktW/
YaanFR3Xb1yzHarvomb1umoysdVHtndjrg6cMtsn71nhVaUO9FHgbAdPeojegmMX5apd/JVB75Le
uhXimb3znECpQJcQFFpSxE55W/qajj5KfLuwQrEto+hNqSmyXJB15BUm7nQuyT98WGwqMbF66dNR
v4eFCauW1PSGvlLQWdP9cST63m1ipOPn10w+PEm62DQUYSWOR+0tY2S2aH1l697TiUGm2pWmptnE
qBnkM+nkTLscJwZ1i1VAKQQtYiFrmGdo4V6MRmxZUwQFLBzoVpXx4/rE2OoSZ/8wMn075e9If9oX
6Fw0O+2p62Siuj2g7SMg3O/aNSDUetnd+PLFap1q5+XGfxeLByEIaHU9MqFivIkIgdBu6+ncLJP1
CxlbIxsd8FTCm6m0OS1WCJ19YxjuvrKFMq1Y7eRSW83N7kpWmdb/p8C+yUPkXQ0BfYOudWsmG+WC
ee2PW2p7yF8IPpblKNlv2FsX6OxHZPuqtEiKn6ae3IuSzfmw2nC0a3ZQfkgl9zpRhXMh+4hIaXcX
5lZIsLHVYHbNgaDWsMZxgQaRVbNxnI0NsQ84qLJ/DpZW+Adg3tiDgN+YstANyKa5g8Skf/7XXOkZ
8xNdlaZCRHKzX3ArgpBahpGU7WzxXJxNrhp2HblpP/+3d1oE2nawqy/iX3Uc3zAAi0ABFnmMgi6B
capMHzI7pbgoSZk2q9uy7qeh13jRK9sfx26EJ9XY9akvcyUkTsQKNrYwasnWy0201POJQbX4AbS3
2BFOGjwReWJOmULuzTNbKxCUO67kr71vvp8xjwVWGx6BYN5PXg2L+/ORYjq5SMk8sjmLdQP2yGWu
KM9Df0NhIEFnn199gxicpi1JAvebvdhiERPZKiaf/AuzE0vThd+Zdr0oxxycZ+sdIRQOSVAo3SNu
m9emlgR0xGmiCO6KGa9N5FcYXiP9qE5mL9wC2GyURyWJbaQJG16Soa0BAjXB9ALK3cMcNziXu3Po
mI6pe6De/RgFsKdD0al68/2Un9x32rXgQPRQlJodaWgE9rUKNzpUC/R0qk+K+g7oFM7/FWFk8Ll0
S6nigfpxme75CP5SnvBTNcFuSwYeUbBzlC+4EbfMI6Qp1gn2kvr8MlkfYAGDgS/XODVDvugz+KYo
7imGOUjTblavR825kXBRFbv+yDe/r/wuAvjhMuB9z+mV9Hs4O9AILra83iObZfBnnmGGN0Jlb1eQ
rCvVsPhLlNcnLiGj9kIFgh23u3GwwBnjQ7tAfCs644QDnpTgvzDg8MFHYQKatmA/cF9hmoxpnABD
trPCy9tzF9QrRat+PTmJiqAZPD6SX7UjHSfn9o+D9TkQrVzCDEe/SRcHsjvhd2x5Q8jxZFdQ45VL
yr/IZsMIp6s5T14Gy6wYgygZrwWbRPRndpMiArILNu0c0deZ4EJVji0j/sas00Gg9S1HldewAfsN
9LuZcV1klHqWeho4DlvoV0RP6QujvZgdzLGuc57vZqq+4QhuUbm63+E/iKkUE+MeA+MYV8PNXQH2
9UHIMXFatWoInJ7ba/KLEd3m21lZV+h9trBRFB2Oy+KKxgaBL6mgkGLw3shyhPm4TyhDhS9IfHuq
O4jIvSZn5v/Qxo9yQFMsN+HzOMDRr3NDxYSUmJGHb6CS1/+VNQxTY/suSptig0FscHwWb/bH8y4a
w+nrvOErfg5UFfWMzJs0apw01ENhVVsQzWsPLTE+GT55PN0bKIMx9xB2XBMwHNXRInssBJC3NziX
9dmQZBesIzhdUmzbBWdHsyNNkQLj+4b6TKhxFgVM8+AceZvsuPelg3rkRq5AuXW4WTJrrUD7HovZ
550fSDk+45K3F8ShB+FMBwV2IypTzw+8mhl01FIxW7tBvIGKHaaRmKImm/Iy0p8Jeo6//Qf0XsJ6
S5LENr5LFLeAJK1TdvzP9NeaXP1APObjT/0Aom+rWO9IK8Md+cYKZDh47KV+M4cztTlCWIJ+ND+T
K3JBwHTme+ocq8EZenOJifPyaEZvh2/cC3w3+Kvh44q7K90Bbibn1Lh9DZXWAUeV81xiCSYOtRGN
A3vQ6HKoZE/pWrCrPC0mMJUkbgr21y03Lmv6LoBNf38UcOcJOcvloIEcJIlCeGJVm6jVGpSxBmtg
tI7v00V2QCrIf9KecfA7f48o3+FG8/OvM2YoOyLKaUQ70tKmW97D/2UFoBgrwyAzYPME1TbaHNiu
OAcpqYf7BtoK6p2CwmToJzzYwTQ6ONtqufg9mxuYIzSjAJUjtINVlnhAu1e1XUqqpUGsT2APV8Aw
3thyibKyEmz4ZebUSocuHJlEOWAEXx0P6f05zmnCxJxbKBbs5Xsi2vRbVi8cOIPQW4TLflv0gTtH
+kuL9x6PErTStNapdbuyEuJSEtJiwZgabktLwNWrt0b0dvNNiO+bcN7URNnXgpm2lTG/wVnILsZu
Hip+y44S7sjDsQtTBj/K7zqRsOKAHp8lkhpTjdaa792BsEMcBSwaCEshjG1Rcr89j5BtOaJOvTkU
sonBFGoDMX277N+XKR5nbiGTuggpetwhPRDrbiar18EqUeUu9fwasnj4RZ5G0JaQYH/BcWb9J6da
Bbx28ysqhyAf7ocdK1MjFvbeatxLFCBO3T3cH6UDMkA3MSB88DgU7tr7ePKzt29RQKSTEafXP5K7
aGjL3o9uJnIxEVRY3ymb6M6oY5OyH3VgrF2pdnY29nZkr5uR4uacncJtmXlP7NVthGJAd9CFtbQK
btctVYRqK66DMrmXyPq7DtvbUNuAAHuay0/sWDVbKbm9ZJXBz84Foeu0x4D6iDdjt4nCMwLaQfIq
33kEb8KdS5mrJ2E61o5oEfEMwrCAK3u6vmDxIPD+lWIVtKbdIKstS3llWQglBZhyWZ1Fmeb3NsWA
4J2Oxi+YBMGwFo7Qt6Gk9FdYDOmmt8l7CKJmj2jsbDJ8Psq190zOGL5bOXB0vn9PEYlqXJkmVdnG
Oh/U8tgKChg9kK5AAblcoHtjf5EmFBqdd7NRh9+C9yjxkScy0Ek/hn3P6/2reDgAQdqIHKCr/m+C
XGSVRvnaBg9K5ZwXkwE8mz2YckEpEOAkdMh0Ib0C14m3Ygc/3E4s6Z7WJ+ROxTDv+xcnlVSOghTg
nZHQaLnySZfnyeIR8Iz2koizzafXOgRapcH7nU/OLpKQ6JcmWirtj/IiVGwYoOalU+EG4vZDp4J8
1L/hO0BXmNwD7SNs5Vt8QGVfTZevCRkevSBtTei3WAW0J6/vJzJao0qPY8vxcDzsGORW/kCD6DIW
JiQoRME8+kJofXzKFogF++tDNTTvh2z30/RcQsxzqOwCmrdSh8pY7JWFSbQuKvFDT3jjtPTWTwmA
9GDRD/6VKUwknPIaABrZ6y9SasRzYiQAAtbWbipH2l8kobNRZVcVRQ/65zzK+gZqswoxJdRuDjuG
xCZOjmJdwId/aol9zR10lLr/JtWHtFtXfErd3LCS5xtPNkKkon5cfaPglYSWksSL2UaqknkMPffs
r6MtqtdByE+snBRrx9pEl/Bcam1OCzdpceEa6XKgPDwGNZYp/tTjEsqxofh1SJio4AIRIVQhjwxn
fnUDK825yTY/fXlTgWgupKvSWQp5utdJBEgsUhTTb8GRCUO75vvvxEpH+TzKuZ6A6dGYdE9lerui
iBRqW/4gxFsasgzBOFvQkwETRIQRSUwWcjX0UeGqkee8EC/1u+TZVNkNpdQVhwWG2+a7QJVzhOPu
TDTHdp2gRtnnK1iq5zWrCTyt4cDzmwfkEukNBgjYmsn3NwNSSBkvuRnbPSNU6nqG6q+o6+1UPGYp
RGQLsnmRFeTMqEvWi7+Q5QOjFFFCbJ0z0c2bScTPGtdYxeIDtnVLKuCFWykv6cxjYm2ex1FCq+ge
DbcYBdpPJeY7cgPpM4eXq4b6PhQU0tQfilJT3DRaeOwJT9obcBQ0mqJ8/UcGqR+r26sUl/lpHbC+
WY9b8JR53dxQU1VVXCUL/SZmAM9K+nEyHHUTQc/1qhNZqc7iiWMXTXXDjbVW84IHCj0Fxk6uAimO
sW5BLRIB0i5Toir/YogGPvquymzcvsQQVitiz7JxpUkZAlkgmrAzNOhZlHZSUbRZ9Pt03ohfuTEV
Ig1cmYm6R9FgVkcS0x0DInP9ZAuvj5h3zPRNHEQgGMp094siXBuMJn2+nGvvifcNZTkPrVoH9ZxK
16bj/qnDgDlvtjPq71SWvPVcG9IJY6caoeHsEEMM9KkU0FW52a3mO/QTatx3xRuTjMFvROPJRKnh
Zkpagd/kQQc9JyHPLZ1RzJfrCYX19uskPYe8X/FrOniz0JuP74sIgEDfzo7/4t9wyCuQRn6Gk8y8
QhlEzz6kyGIW74Eo1rrJc1W27HeGWylsrWlA98T+dPujmQyJZc4bc+lcqCDnk9zwB9rvE/z8n9wD
TZ6CWz/4C6v1E3GrkWbSWCo9ImnnMTZL5kBMJmDNvDxXwEaS8NYv2xxOIynDqMQNKM5nT8i7Vvti
KB9fQOoP1F/z11Wag4ZVPlBFw/U6wra4+ej4icQfk+Ao4OCoxlo81zxQkuomGEKV9sDnmNp7Vt3q
XUkMYhT5O6liHsboKLTb3xium7vfTQgE3r8sRNLDvMUX4HkfzV2ATKmdn/ZwdsH5p1s5+wuBB/Z8
gVQlLFLxw8tX3UdNLaAO+PtHv7kyPvYu7UzveydoN7B4hUZh0kzMtwMCohWy6gRinEEM8pS7zg5X
D/TrVurcrDJKyzT4wWX0HR99MtDKCP7ObwZPVwug8+t23SY0kHglywefJGmBx8sZBp4/Amukaf8t
9D7WRpjFsv06o70Tii4yy3TyzjRMrvBFslBy5JlBNfnKVkucIJLLu8S8lC8HA0xyM0XUX4WqF8G8
AcPQielwhAbgSAKf4iI7gseni+oCA40ceFlx1F6Li/4SJIV3r6Qin1LfiIHvlnUV2a2ew0ZBhG8V
LnYCPBeNHnn4CBYuMORhk4g48mLlm4Dbl4yoQLd0f6MksQZiUPkUfFmWBWIgOVqMpG48Nnj32noY
dD4YmuqWky0pdrWfjlFLfu5oyqWKlHcrMwZMq+DnF0Yej1KJtcwfIaC43UEEHypIwtXENjJlQQpF
dAbpVfZ0Tvbx28rgfoeVkJJs+yGxcYq3Yc3IUwouMW9WEM+lBMLRrVW5GyPb0bzKNV8ZPbz+jX4H
WP34spuDa0T2HX38lBr1Ew1Kq/uGkO7aRssPq8+T32xpE5gXoPEArsggwEgQYhdESgrvXxL6iGXe
sY66vYX3pnjU2iphBc1aUlEr/IuEDUlJftQkx6OHkmtKlA34crCIzVX36pHRu/SJXQbWM7rEJIwr
llvXB4T05ASvoDFpH67Zwe8uc57HlojmZ2B+BXknFt1kjBMv2fW7RRCnDMbx8izP6OEaKrwU6d+5
a0QFQtFjKIP0Pj0vWKnw5clOQP5AFbJ6qb2bpWSlKkO7kFpFD8MI42emh8QoWHXASoG7Hbl0hI5i
SomSE+fKgAa3P6ZsEuybnPDrsovtdwWuG3tsP0IFznV1mQ7PYb94sO9QQQda2EeBkpGy6RPuwut4
3ddPlsjMffnpV62EKUtcP+ZOc22wtQJ4GcxcrND2JiRwogkGshkbSlahpXwDs1Qu7f9uIfklKAV1
YTFAuwK+lHskR/yR93eDxhVbDJ/pNZgK51ucdHe5EkfjtKs0hJS7t8DP5QVnzUwTd86MRA679bgq
tbGul+6vBSnRwG7lype/iCyVGzQ8vcFpykfmSMsEF4VqMfGYFEW/Ki1uI4AMzrrT83h97ZakBTyW
032dCTfMS34OPpmoPK3M/Ww5/5Nggp2QlMWOIrD/vlj7MEIkzMPIBsr5jVRPHYRZkTsFUxQD/PlJ
xLenVXscgxfxH7AYHQaoDNnzynbHUWtJJp6Dx4E2a60YyHWsSXr63yTI+x9QZ9TjlmidyRjPAy1H
nLruBYKE97Ug3B8GmMKtFdEdLtjGhu8ONiHD/r6n3xGZ6l8teGeoPbKOKF/6tR0m62j1sbmGlwgC
+HM2G5WwApkEQf6K27B3IJQK+TkSptMj4vzTvijtlSFG4G4BOckoDnV3+OGIl7ofxnP2Hfp7ieNE
xLhQb1RX7tHb6nB+MKuwTLA5AIs6f3zxvOybgLls2fCrQbqor3VW+XXUKV529ELcbwes80+PEqhg
BGLFfIaBrLmYnE3shTnBx7Cy6rPmF3hC/+C7ArLkYt4IIWaBZ+hz/Wn31i+LnAPIjaKyEY2vXQhU
zoDjxMbw+3qkKmk+6cr6llJQ2Kxask7i34oz7+WMHCqZ8lB0CI9fkgySee7Xd/HOcnKBUfQmMXwg
x27wRWdoC8KMGX3s2WFMnUd9lR3AIlxuw4d4Tlu/aU60baR5Jf7i7IETbJG0ddRws25iEAejyQd7
HsBZPWXfh4XzgkEOS8Ek7uz2iHwWRtZmI6PwwYXxXDAF8kfbrD3faknTYJn6QCJSMPC1Y1Xg0PXN
EFuwMavMiGBxAsyLEoNOIPkVZinnCJPdXwHN/TQjIt5VMrP+ky3nV16Jk3ZMWGln0co+zwVQbA21
RBWmLLZKbU/K/oIslGxgqpjP1DdEtGQ1pIsg7pdjbD0fRU/3gokFfb4I9Mlc0PWFZjoecV5HX3Cm
Sy96exPetDzJvgnwGhzhdPtPwhcwkilFKmxTWUIf23YWSQ41PdiyayG3UK8emdsppMocUM3x0JRc
myJIgcLc06JUlkOuZlu8GTBsozzdLmXOMae1O5hEVy4S2GvpP1gK0aqwevBVVa2WVk4hLPIx/Ivm
qJKn1AAf8wuFkEIAWpzONPRjgAxn9ZmOyr553cLwWYF3QIhiGCsNPUqlPBXxS7A6CXP/Yx0+7syt
Na1AKrAWOgVZnIbUqNodiOxtZKUO9qD61VAR+RRIV0H4Ga4Et8ltYTcNvfBZqnDx5ubWJdcE/oFD
rCIU+2h+j/k686YqXmftz+t6DsE3gT+Oc7gEpt3w6KNn1oMxoywPe7xZcK3EXWBTZfsRQBZC6dU4
iSzyYsqCIkpZLI5r21SyBWOlBAxZGkF19b2UJT8PywuwZmBo/qd0PmBmqv5SqorDxTu/dmswlgHZ
3rUsAHyQYa7YUH69vmAE9UQi0OcI4glXMnRSCrO5TMEaNW9IBqnIBr6z9XGReivuAjwztAmwJZyM
hc5tWQnvNrJf20vrCVVyF9h2iEFIgf23oLoa6e+10uSdaSs9U9EEsEdojHH5L+yIrxPg98i6lNow
mknRggNb95WT+mVnBq99awuSg4ucnUZ6KboSyyvQswjQ5elAbaqvRhubgy0Ue8wu4HgDxMjBSzeC
Cc0GHJ2fwMMEQV8CSTi5BtBKfbt2ooDpKhmlpueKlydCiCWVUYiRBGsHUyONiL6fYaCHpkulHq5F
MKzPW7+PUPQECVLAt/Jn4Gbi35NtJs33F9lvzyV94Szy/mp9L4tf+oCNPSbggjRtY1dn0Q1zNqbQ
VXO7JcR0eg+TNWENJs6P/H49QgmarHpdln6sTnDNYjYla0oTpk92h1TcEaJhmidi3e8s53ZRysj3
BqBGbuxVXeeY2/vmyCuWqnq8IjiolVibDmmyKTRDrgqNpc+7tRxXioOio0xhvkIeQh8AxPZqS3ON
x+Swa391aNUUqPzJAP+L7HbJPCuUSlA4OIsRwdbft+adhrnjfvAdnTmTut9zYGvk1K1x9c1QOUi2
V6mKarjor9FdsMf2A+PSjvwxJvJKaZng4dcVATvxlM+Dg5LF1jnh7vXDWXnBHrEe7aEeVykwaJDX
7/UriiDuTJXsYfypGnOEU931IT+IwZPSPPgc6CEKZTXUkwYj6jnlBy0WFskHd4Ezw1K3Fcxn67lS
S7MLhMKR8tvd6V5gmnf/iN95IypEkhsZfMOj2OErIAkS2J+YQhVOKOAuMCJp2piaXeBQg0Jawcjh
O02W4Pffs3Pu/9v1AHaBJDAs7ysko+MMhrpVF5KjhWXyN+r5JXpqGDTY37wJe0SUpad9iLnAk5Lb
K1r5y2acMbA84QheTH9RyrnKH87NRn04jUOxx22Y8qk/ivU6Dt8Lr6C4PmNFE0JsOGQzGNsrffP4
+fxn5SfIICR8UX5hF9gRc9vJiS1n5gU8DXVZEyWP5fCPHdjxTBczMm8s3xDS+GT2PHvcNAzffEFU
f1lflYUSh44cANH8Q2Hknpg/wtjoL34mmR2r3Zc2bm/8kPm9OzYfZJe9s0AVz1dfJ+0q9AXj62M4
uRd1L3d3sGfBc59sanhpbwhgDwy+jD9JiV1mDx0K5JO8caXNDTZ3QiINSDYb48/28OTztBG+beG1
TfJ7BjozSeOOm6PLZYpMsAb+cXtG85n9u5dZ1ibGO2J2KZH4TsHcO+cgfKBPcAPdbBf9aHIuJ1mE
6AG1BndEJYPaCUtodoP0bMcsTY+Qg7jB5dpKfrpdI0Z9CGpQBzLz4FFUMI3V9JMntT8Nu/ypZfe1
PFbD+9OQcDWluMxovztwHYauZQ3QEExz49Q50z1PBqUTtkdBEKUoHRIZY9zrlRnXxoLrRBiclSvX
48LyEigemsHZo7SGChuMdjVUMkaeTDshBclZf8HFZdLp6bgBAIql+aGtnu3EWRZnuvYbkoteC1cg
XyfmYaxhPGwWaUp1wQwbok9TFPobEbU3XHruApnySFDp3PBDj9KR/QU5SwU/6qngSw3JQ/lWkKJS
kjSjEe3tvDWxJYyvNgpH/d4qI+EwHS/WDAb2hocR23t+3t9NqMSouBGkJnta8qWxeQleFjuq57Qi
Ek1xyxuyPTgZcSbHgSMpZHNJZJiwdv7vvS257YV4/6PSsQ2Z/6EOgj5eSJ+8WBwV7UA+OV+7bJNN
dmzzuErOsSQZ/ibc86+xVZRnFLXwLsqV+d47s765aTLg5T3BFIgZEqwaJlIFGHKfhbvRf3EW04D2
3ZbraVrndZ/xyEBcJ9vDRzavi1F4gQUiMid8ZF4vEqIxBWtUtPV9T+0wsaRpza47kuteY1ljM2cw
zd4DCktLSgaTIAef46/7CSnH2ADZIBgfzx0kgRfGgun7PuURpkm4aqVc1HGRa+TW8puiIZhg6Q9K
45VyX3n9bgylLhFqBxltEYBZO/tMfzKNmZ9SsoAtuCmdEv2MEQckNIDgqVHppyduC4NS+m4YfugT
v3LpD5mRHq3bhzSADNvX9tawJpQM0MYFjTE/JznEOo/DGf9NPQ8ijjzbFflLEsfNtmkaZX46xoIH
xhRFhqViQYR3Vg8yGAZkajxEIYR+2wbXNqmdApGO6DZZrJV4V31DC5UqKWmCnKJ+UXOXfx26gj9C
HJN/aiuirZyhb6HHPuE9VUUnHmUgc1EVFwSha1Wm34m6XYVurmrWbfKWZlWdy/kmB9qsK2IUMuDw
ATb/4Leekv2Ac29e7F6ISEkPQZXWWlBgPdmQBhSE/WyHoXpe+PJ6gUCTXJPjC2Y3EBeWF7zGo4qM
gpbs8U4gqy6IAwAa7lgOAENpn2O+5t2RPbw962jCB4QCd9u6hIJ4JjJEaJ8MN9fymKsLOYhMTWl/
Od9i73bsfylGHi4t6Q+UH7dxe4C+R+m06tjq6LQW5ioqKqmK4+QebALAmayhegAkX/B7wO0rWV1R
rs4Lxrh7l9j3q+rk5HgOXe46/vRZ6VI8PnpFdxJ+jV66jih+T4/Z00eUJBRaeLGTRPZAvIjxkBzw
FrnsYnY5VWE11Lco4On4zAcbFGOW/WQV/lf42w9LdCt41v14gc5JV8KxpMStiOF93mM98o1WHUsw
Tphq97w7kjOfyPdktcYBYBnZYLCuWnniEGl5o8In2MfuGxhr6IOt2KEt5i0HQ7dxJkGDjQ+RubJg
0orQ8i+EdyUHjwMI92vA7QDMc6VTJ1LsoX9A7mokHhmxlzU2Rlq8DQqOntHiiKOzlUPHKbWML1id
KX2l6hxrvYh9Sl5UMnkGnozVrPuGnQFPlFQNM54DiVAoIkPEJX9LRunSe/uoVMfNlIQRC35yY/xB
a3yT7yYRAf+Q46BeCzy1GGJ9pKtG1VuncqZBuJdLH/1N2NSvOu8wt8QOzV2sjuSKq5QaKSqYFzrd
FVSvsZAE1eSy5jTdyPJKBBhLGmHsEyA/rgKMXRVx1zDg5Cbu/5T6Sk46F0UWEeF4n7SHE2bYigbz
pJYesmJcyNCjP8XOyfXMyJPQVnAGGEr9vwrwNS+E0YrQifvo/cnDxnQzi31/kuwOBxM8KIp0OCEj
p8ac2YjayYicAEwwDlODXRlazbZ80Lmn6s+OvNGxrhuQGk32zGgau51xDipV3lwUDz6QJh8OXHHu
FX5OBAlX4jmYQUiAnZwTM5zoNZHLYhlsvGTUXzzP6AAUM2s7c6QWR/KLpBb3J/wpKnXQEsdQyHpB
TI3ASIcScGjaYxyYICqtqQJLR5FpytSIXPHVT8JkVse3n2YgiDGOvSixi0R23JW1QwUPpaS61yi1
RFXU4wxTFxko35sXgA6z4VkyuteOeWsVHSi8y3kJN3nSTWCSlO0EhRP8ZXvhpBg+2tIGicQCikvs
cXtidAmz+FS91msibDPKT6SDTTNf9vLvLjJProh/GcERLTdAck+T4FqZNCvT42cCKwMhKbFeOXKQ
Zn6XHWe9/rkEZZaufGi2nTBBCC+BqugC6nPaEd8v7TcRTw+Lrvcr4DQFkOo0O5zuXEJ3FndoM52i
WzKF5k9G/5s0FL/aXEyG+IoweEV+d1XAZ1eCcQ4w7DTV1I3QGoTe33MqHfwa9r2TYBl3jJgrrV+P
lvli8rr9TI5qXQ2uv4duGCR0gt6K25JJKPHG2O3mH7YmNEgS59WqX+6ncmMCmMQ7jEZZdDd0HRGU
DeEa4JFcasIvIkpvHKl8VI4BVaJwIbUkCkfa2mI+hEj6Jr6YG7GqQX8AotvjWk62s8mOjs+ZycGe
1SZneLwHM5FABTJoffM2pMW0qgyAf22fXp8vzv38n5b++kNw7XDNcfgFcDZyMh9PT9lD3RoSP3Oq
PD37fh2pkBy68W7w/pQStSIfIdii62TaNhbc7Gh2AsFFmxtEIybNWEom44WHBS8lphxh+l4AL/X7
LRRr69PV0r4UqJ5KxiQID2gy8w0nmRVyoOJ3FlDcsHT4u78laboRAewtf131XL/sE5hZ0tEzG1cj
a0p07KeTOxUBiJnaJpgfJygQUb1JvrxkXIDn+dwrJMgClno5dwIveJtmhoD2r8OST6SsY3me49Sh
UT1GAxDeUgGxBwegLYQ6exx28+kUZCTQRAm15lAtbAtYFWY3xwJBO8iXxzMu+i8phVnNRP0LR7W6
w9SEQEa/2IQk7G6VdLVGRBDPlMT4uZF201JpBgWFxthIRodTAX9Cmz7ocXYuW8lPf6l1Tkl8OIPw
Y7yRogSuW7uuUAYoPRKKOjJG8JwAkWopOpdqGtH7B2wPVqYBfkcq8oVO++BUzY3bXjtdb2fi/zEE
CubAo9JoZ1LTJXRaappCgFtzH44Lpydhujkl+tFYa8ERYV9WoLugv7FeHGBqHZA1ylB/XThp+0AF
MSAXhzG69mJsnsQYPiA931++ljPhGHe97jUiQ5bE+FJnc8dolodQMtEYajr4xOA7hCNMF5bFmDRz
8j/No+My9k2gtN+oXNnVoBL97Iq4xMx/CLfLPgXd8dRGLajil9Lab9hg3Fvx838qh6jt+D+NxqE5
cbnra/hhzSSwfj5dKLBzBHsvt9N1GD6n2bAS/Nn7OyV8s5zSZQl57eo0ba+KO/uK0jCHwatpT65n
d1+Gt3eIF1gixL5Eh8l58PalTMB1EukJI0U6OKSmbnDgU1T0HE+y9I5SEqA6x97NTBeEybUN6Db2
S3Q8Y8pzVrDYJWmtcS3L6/ESRu4nOpMEV+ARSQ1avKtt0wreORaPeljm71TLvq637Xi5NkY41zUJ
UrauW1E9VGYJf9FbL3/v2uq2HXOUs7p6+2f7tRgS6vosj6I7ILOwx6bJ3dxsJDedOmKZdW0NMgue
c45pNBsB82amLlLNaVtTWgBvMneoVcjxQF2VzsM+9hSMwfq98O0YheunE5Ox9jjpXK7CvMv4lyMj
6eNbQc772RQQA2oOLBX5K+Rc9Kbkx6+aIdO75AiY2cjH9ck59SCTX8WTT7zvBxwiuy3c1PyqF2FW
IeQECZP6tFXO+wIFGjuVfxENRjPsQ6kcw8z6k88a1BckmILBwrqbxs+hXxrFwW2ucV1JfRk9ng9X
PZ8Zw5OQmSV2xh+XEVziWQF6igNB1h7UyxBHghBc+rmv7bWkKXrJvljMcOXAQ4edDlMkmF7638XK
OWddhNcVrB3DihYPCmS5PY3/ZNB0lDGBp0UuxXOEoCGvLsbxU1N9/mjkuXN5F3WVRl3Zh7iTjofd
fgJ4mt0ZxA7NEqyYVuBd+cWAusPm6p2XOd3v4zhk9DFKlPh5M+Ur/Zw4xstoME/GK8hCRuSf/T3I
lRmikgu0i69BWpPChRvMNLGPf6yF0Bn2jH/aQiFXpUO4pVe+Hq/OnfLEd7zc1gEJCAgPZnt+EyRb
Zz4ErzuHFSEcNDtn3RQGSIEsLl40cnaVlpFN1Vm+mnZdoPVFUqBTmiPvCtr9XfcuxVUreg/Jv9Fe
+57Xgcr6xQqWeom9Yk/7Edg7gfVw9GyUNU4vQvsnMN7OGm3HtSqa9qIjmiNPr5sak681/zY7qTZr
oyqT7Z9hUnYtSIytxmF8O17LP27zWXRe5/juXB4fLD5d41mBFUbLJk8TFRxSTLLB8T3t1o+rygIS
V26eQVq+RiEHuoip2Y//eMgJtIbYsjhtVMiTRtVBj3z/ub2PRvaAMGmjZ6ByEQuFIBM8bQknzNum
AcmNX1b7upRA3v8Pzg+pVHhEKb6tT6Q4ImOM8AFRP4E8T4mfcPpKUiRhQG+GvGX07CO1sDihvWEB
WyjsPEEMsDCPRKJ2X2gW8LV82TzkovzyHAsdgr5YZky1fDLrm3p9JKXbvZRVv5RFm/SREbolSRav
6RGz2tZHo1naI67mdCmhiap2n+iSHfiDDMt1phU6Syo/yDBnhqzHZC6oG73Jyajy94fB6LZ95cp2
A4zDacrvZLO7iNt3voPlV5sOQz2Fgo+CcG+fRANjpNnmx23n6oYo7MEI3MQVngVhplh5QlNGqwT5
jbxY8H6W06RVKJZ4uNJAnXLoBUyxa8v0R3znVmjWOLyvLf3v6dPQkTio1sR4Y1zWRJhHOvAnHKbF
dgDSvPZQIFvDIiDztzmi0OfJsKCjSpG7SGofmqmpjW5KXeO9/kDPNGWzTWCVRULDlf4X/bgSigJA
P1N8HQejs1By5ouCYuxH1ec1IDwpOK1iLixp+808p0M9WVCdMallHjCDW6dNu71O+WKUXPW1VPqo
S/eXixSn3wQ0XQpTwO409LvX1f64QK0J8xZlXiwfdVK4g0IXH+guL4s5NsgICj2o1pxb56vHuIWs
NaD4Ip0jJULX8W9cCVQpjrq8uCUPXvAXKul3zCtv86npx0jHR5NHlpWSFXoXlqGnyLtT1W1amwrD
fLy3Bl73LSxrxtaDJYHMSqlipGm5Qf5uLqIjOrW0fWRGt5gztFQ0WCuD5+PCBnjOrGLFBZFcYPWO
VrHw5XZVc9bkGX+XLE0P3rX8R90xum48ojffSL1BWFbNwDdRYkrcq02QF3rNQAFzV5/59JGrD9wR
L4Tei3T5+L/xf+EABb16zT0bIDChtXSkhGL1ZUVTfW5V4jlyIQyvDAzMNnBM1wQM+tR/GDT3wjDz
LBQVTFUhve/0zYDFFr/HE63HOqL8pSf5tRb/RWC5wEF9XJktHkq6EA+MvUWEvplv6KZorVJOTH1P
nfmfFMYlBAWHIexABIxUhapDFctbDhjrLj+H4+w2DsQMbm6cEjErzI6zTA3nu3/mY7qRIpnVNOKI
NXNjZapNZxhjfqTKPXlU5LqFTb2auiFkSdxrgO+wCkP9L8N3w9FQWXvaw2BVrtm7PdCh5dH3OPQn
qoqmhJWIVdYqnNodgFMaN4P2AaJGMQhGhWVsMxRCp6jRUPeqpUjcj8gBcurimFU3IogMBsjup/eZ
Pe1M7SBbZBJsVACeZvAzA/nOl5MPsXczFl79BpsZ8FebHzZV8qKGHl2QbbCC0sHh7pUmRmwfYvOJ
cm5Pqw/IcY+KYSMUIQows760iOwYtc7LOCkXuslcrotZ9Ew5xIWsegGJH9lCIHd0Kki8a4yCMKbR
P3gKVayv73jd1tSkG9lyQz+0386x6j1HisZAXvywJuw70xUyEJzi/hzpaqQpKlQbaTDNfUSL6x3G
upamPR+0pvfuAtH0ufRhnPMT/x9RM6sWOiOHJfT1lWMSlNK1hJ7agLCSKKaJMoNMTZ8vZZRl5hFp
v1889u8JxUa1pahTC9sezxYsYCKywBN+On69kAKZh42pTy7zGy5WQ7XfZqWBq2ArNbTW7ErlCsNX
LCweiJBjNaS73y8CUV+XNXhRsnykbDof3WNX4hPStkT5UlIre9Jv/H2vR6pyYrzwgeWFxpdeO/+k
W427KFTCi1U3a1TYq1cVhc6BGQvasxgXC5DXRTUZQePgeKPNHrhY5wtZDBEK+WelPTO+JKS6kLUp
nYWKTrIfqU6b6FQ/5CQfcheWiisSwFlR2w1/7IQVgJmZE1jLKDmT3VoGS/ZLgc0PqZ1H3rRF8wUF
Y6rGtmUzSUx+Qw==
`protect end_protected

