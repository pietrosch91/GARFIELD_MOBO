

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DIIXDeJza+sKqBrj4qf+gSpQ5HFYwUFgPgXoi9a/661p1fOh7GC1Yxr4QhwzfxxbI2esRkgX+RWV
O70wuqmd6g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tc3vvZL4Z4/k9lIOYWoeVvOilMT9DFpT/2Qg9j3BlHsCcWm3A3qs8Rzy60Chth5nEU3HV6KUki6A
hRQKZNb1v/6vjwTmXalrXjELjcws7f/IYaWgZmjVdYjpJE/aoPqNISqRAxye6F73bRYmttkSLsKA
mpZhym45OoX2lTi2dYU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qQBOLNsTpDaTilOll0jbdzN9+CFe+2YuHpSZBsocYQBx4tFyydxFP4QWzsgkpKMVj+vgHsshU0FN
Wu3IvX6zwtMbic8Oj5a78zbLuCwQAJkzJHVEC33oza9R+KKTeRuoZulmj32txP8npOqkH//3iN6m
rbkJ5ZuVWuWTahdk1WIS1WH0JMwmkoMmZOzkIvY3OwyRzQ7J4JWsuGgUCQP2UiR1wTcS23zdZ4if
K5dX89DOQ5XLDZRfGBzqloRoc2KLKrNKj69bM6afBdivLgfZpIq8pSaRYrb4D4nQ/NQLMqKVQM7g
UtRkTmmMOH9irg/EZkbw+ma+qT3UysisXvIRjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FnYKQSPwFxsA2Tic0BZESWi6Be2FIedgCX7009o+DpIyXr2I2/Jxc6RNA88ViWghN3LxaxRvHMEk
pR+MRZPIxTWv8WVlO2x5IF03WAJs9GAB6d9KbRe6Gs/fOQS8fMMkXpyEq4+6dsQ1yT9ckah4Cdmr
T2dV46kU3DtfOZwlWxk0OFzQSvWXEIETRCvrsGEf/mlDvxo3c99T8p2n/HDBiBrHIY+98bbLLHvl
mVYYFNZpsys4uRT/TVeQxVr2Ro29URGWoe0peT9xCIdU44Br4X8OPNWGJlsWrkooLMv9dYIUEfQK
VsblVGzcgvRtwlSZRK4G7ikWOKojLVBxgIsuhw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k/CEKtjJXdiEV2H3DdiRA6UDxaoZt303yi4S31RTSRFiDtNKXEWX7hAbczUxcDYrAZq9Pa18y/Iv
ju3h9ViJ/yaF+1n8xAYTxusQZdevYvn8leKkc+XbCxi8/TAYj4SQ2bTf4RMijly6zLqqO004hHo9
AbWF/Tq5CZLrvf24Df0yyJWZTL2km1BM5nTE6v8B0iMxEncPNncJ1g0VKySbcBDCh6+IdZeFDvjk
siaQTjWx1gj+MKrM5hxCdh1gK5aVhC9As2wDY0avEH+1IxuO6QhBjnWFKX5v8fUQvgp5zjSufCpK
Ff3Ce0pbO40TcP98XMg/XiCNI+dX7w8S194wMw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B0pRxV4llSbxSsgbT9dwcuzImsNM7Ywl/K0BGEC/Mw/vBjKJqOpZbs/20GVssjsAwFuJAwsuRvU2
DcscqGBWo/UUVxZ1dW+/mhv8EMGY/gglmOl/jSYwQ7g7m4z3an+lZM1T9/p423pPW8FVM8MYisbM
+tyxyBR/MgTmoxWxnA0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EHRObHCL8AfvkiomPbt7c3iNsMF4eZGxQ33JWJrsuaoV9trVmGm8vEcVPWLNhGAeekB73BJR+LiZ
zi9a08JnSoTsgO+46uuuGrEM1IK8husQ9MqNyNGRTbups69htwaKPx1YLtc1M/60smF/b6euaSYM
JSASlMnD29rew98IbsycQiGsHKlati+Itr7j9mPAlgM09poau5yONp8Qnq4dT11PG2FAMF9RKNCl
UCdKh8nmXtEmrpJH+V95f0ogErBgKxxAVi55Yvtg8bgVdXD9OE1BJxHTIDLs/OWMstM7CzQdhFwf
ujlmDvylJDwTSbP429MwLLobIYUiMwfATB7Cqg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
90BjojWW2TzVe11h5C7YkeY2FL7t2OFZ7sHpmI/fOyqngPpUOYZnECezMNUIN3Pcr0qbrUR7RJeM
wtVtpctUUZyzowYY9sGyudemoWcgK05DYhODaYp3kBTBQB4/D4EqpjhljY6+v1xi+IYz8hrLl9gH
SSkXLVrcmVeTJ7vFJRfrjGpPMIgR3Laer3x0sKdWALWbEMj1c5S0dhy0ZDbNCDWu/fC6iHvDkrPy
hAgGoKl4mPgC1sIwsYBhZRGAYTVCVPyG10zb3hN5QBMXBkZZzJcHAJJmvD8R9oRAoqUlzfJaQ6Xp
dCPPjfiBnwX8o/ohC1dJVWK9QW8ne7W31knHzftv9KNjYz7DmgWICTTcNl/6KJRJ0/Kyir0v0u/F
Il4P1MsJTdOaXLoT9B5bf71nCtLlVev1sK0jlQyjSOlFz0gb4Dwl1uhFmHNC6B+KjzFPzpF7QLGr
Z41vIKuH5AsTuWLcfcBjd5GIrRtsn93kbYLRmGtVntEkcV+48Xx1zmX7ZR6yfu7iKRIz5gyw6yOI
Vp/JiQUfNoW5BS/C0Z/sUQWIge7VTlWTg21r/3KsxKjHCXqBumBiQWgGssuNE3q9wb0ToWOgZ5Ye
o2U9Iga3FAqQRIndkcXS8xwNMpm16XiA4h+ndisr4kK1uycjLgjLhKiED6XfWRK7jV1aADTFXS7G
WDA29d6FCBpwZTqRXBzu8R3ZAyt87hQOxnOZ+QSkvKJHK2touQMJh4G4puvbEqcNaWX1Pg7cizhO
lSTsUpvkPcE2Evt5QHpGbpeDmpBZWzvvFQaFAHcgPG0kCdlllyN+b/zjCOPj+IRkj5cMXquVUVv7
bmXlcqCNT5EcYPOqFPADOsoSjcE8kbFrFu5l4aqzZtzyTdLGoaKkboqyR+weGNOuWwmunNY1TZ3A
Cjxm3KlcWANR/Ysb+NQLBesYr2CQzDMIxZKD7hS1N1BT0hPRPrhy1jhec52YfUzw5WRtw2Hwn+gQ
FyFfpVFKogwG65b8I+aWZ31nv8/sqsnYL6PCwaBujeaVfN6XQ/AyF6sDGf9f55RxsLdZ+8/EoS/9
PLVHgXJ2RDLei1Tbux9nqaD9Hb9MalmtyTzqUPRFbKJ8+Ajq0lFJkBu0jtksIag0WnWu1tYB48pS
Gi72YFZjdlwoTJugz/2CD+4PaHUlWUmkTHiTeUEUrrWT0w88alhIWJqne4oMNE8J1PKwgdB3RFa1
ZWWT2qPn/FTsjuCYjdvHhly+6b6lI/Kfi5L0Cbpf77+Lz9cOurfryoamqCSKxfm9eSc1hWLhzCX5
uIu/VcMjfwn4Kf5JTBebd2hEHLxFuDOnay2ka6rKgsgE8hdHICCGoTUHPi1x2emv0pwfeXv8mi+X
M2tfHYaMbQS2D29XUbfdHrfAVbuMIjd4xfh3NJ9lkTnsH5xGBAS1oylBvaJOtBHRy5401jJnTXqx
JyAuxAN8wWiroPxChu/6CSxs/mIuiF+Ziu13QWb9oTgA1PFIUshzBcs9jGHdzmSR+CnD5j0Q0TRe
5qit8i/UO826PKxEdKqfh/x2bkk7ifEdiCQA1TKoWz01Zps5Tvn+TJPCSIXRkeUOFDfL+kOS49KD
3Xop4mLKavYsn3BBSRUhBsIhvQJzdR2X74ZHHY6sKfd4nR4HOiF0pCKSmM1QLr1i/LN9b3X5RiAH
/ORN8I6oYaQWYNuCgEOJfrOJ2jtYOchZQq8AM5s6CN8FVtLk4ll8Qijg9gRmZ/cpJv2qWxEhZWYH
VElA+EHZFxWSRDAPV0suxU6VKCoQnm7bf6xzbeaIcbg/UiBOEJAyoOyjXYlc7NDMm1X3Ge+0Enkq
m30qM34NNa8NGtGlWb0NPd/JUs2tWsIwbqzEc7wMtuE6xxlDgtG3/LzP58vl0n3n4wHBkyT0a7/J
Vfmu5n5LI76BtWaR+fufsO6YdXBFXQgZ94uCET053zXop8Xr2QT6WEb+K4Ldjy2laBNLg9uOzoF/
daf7Q5h7bnz6Wc/5q8Q3KhhQYmBFRcXSmCFChVDscmfCh3kS6nRagjwgjLB1dRnMlucpaHBSlaZp
RdOfGi0HtXtZwmvHPePOYRN5YNgeI1267ip+Z+WhdFjunZkuCXv+9nPg9adHbyTdbGc44+sSfJqP
+mK9P704LUUsgJ0jrXcpOpFN9W/BNrU0zxC79aL5ogQVCf1QKXKIY5mZFTQnCmviGChNzOR3vTrh
HD5CG10GOEugITpH2gAeh/23e8ZndRcGZs4nOhVrOdQC6K4upaGSKvNZ6HN8ugx1h56mK+mWDrlD
gGxaxM8baMs8/l8QFHczYyM0zVk5P4Sbd60hosgbhcobX23MxsPEi2Wyvo3OavWRn2gMZMTZ4Kac
C19MhXAI3EFuAW258mtQhx7yBDkR44hUfKZ3hq9KN36Qjqy2WhqOXymVzMUuAngpmluc7oqlxKEE
sRD89Z6m+Lu4IcqxOeVYUL6W2Uz2oPfd/gAWmuOHAyepZN1QgYK5UwK17DtB4cmmbsLG5A6t0J0A
yLAHl7WViQ7/lMr1WgEPAqDSKt0El+0VXV1LF8mOXU5NTyNsv83S+mr82+W+KLCtAJ5HhoP9DnD+
z+Dp6J9Vcthn0NDTZV1PjK+W8aTxnnCKurP9MUEj45jTjPDJ4bzJP2/Q7EjGuGZtuYiicz7DoaNn
sdQ+GOg3OEAIXaJYtJjzxayL4BAQDSFdv8kt6yT6YDu/cQFeDMaldiXLcRdM71RUVQpUBkw52Ssh
7ZKJMz7xzVjHgfVlVbnuebuOOqh1paY9X2E93tqdSQN7HiAbUCNALohdzCVYGZZYA7nlKGJkuJQU
mtIY0SrYTOs152qgEomcJf8N412EBDwWGfrTaqaG4Jy5PYpRuUd1SoqZCOBKsVCoz3f6Rh4/FFW4
QPsaBBVHFu35As9uAVrex9ffKZZvCaUgGYv8VGfKo8+YZhfYgxQJqUNaD72FFaMdmhp2l42pfKa5
lPQ3kyw3XIFsQKmbPO8g2eYCtA/meCAhYbls7hlZwr0MvAwfUZ3lHsXt5rwP7+SzEMpbIYjE7LKl
wtVA+7x9i15oVSVih5b+he0hEz2wQwgf9uN436ExIzJMtQSI/l9LIEUVecta1fXVGC60m5gnE3N5
+iH1Vq4KJk0PmW64xwcR/jKEpRRv0CIQ1JbbokFnf6sKt/iGhvrYBLr9qfzUPnKctfLLGhVUbd4N
VWCs5mYhn8Ra+PYmojiLoKBuPm1/mRZOx1Xm6MthLkSSq9/hbHtOB4fF0ySh452cOSypD35jZq1j
SOHbaftNPzlLSr+PyKE9JYhDgcueAM5dSUI0ptyR+gilV7iHT0WOBILHgZbKxeXNDg4lacXp3G++
Btq1YQveIaWm8jeALlHLBY9F1rMRGu6zF+G7+27IfOGSKpx++800ZWyTT5kOHC56Lrcs4LHEmERU
z/r8Ap+c8x6PrFAzhBpmcVMXNJiFkyq9C7VoNfxJZ7ZD6g0o8I3moSWYov2haYcxXM+c5VzDOQSB
5UssIpiyvGBV8H8kN9OWxtYRGTcop1Z5seVUlDDnjpRfqs0BTjCOidHM7X0NYd2QRMnfUyPx0B/M
mr6CTfhnalkX/vIxpyB4hxvYbhAEzsItDSacPeur9cLzcOAszLggnYsKTSteC4ms9a4d6wOoca+O
Slq87I1Gm1wNucRXaIl54oMR9wFXi7zr2F/PEOIheknoDnmr5an5w3MQenYE89lNJAj0T+87wQfF
vRg4ST4xo7ExO3bIjqUyGLlowbv9oNBmpv6p4xN06ZI6a86cVAb4e8DttgyF/tzdd+8AUuRhd3ZN
LGdOKedJotccte7XE1ANBqMo1o78/HkUfEkAqjVOhtfZM+WpGgJgjcEYEv6lVqrNYoEd/7UT0mJy
SdW6JJMx2uzVZYi+094bgu0fpc/gKTQCDZwxJu3JRBYNYUzT/Ge/ywBMrWW02G9RoqjTFCQOXz49
8htxIZnuGyYrAci3TvwWHe67AaMd6Td8GxrxP4aAlt7rEu+GB//cA7ADUvw8sJS+scSm7Kf59XRE
rSPd5A+uVWEfTCNEu1PSR2t5OfkKPykQcINfZe8hWULihGDfzscTq1UeDNRh3LSmCEituWOphipI
2dHqjAp/BwXywIUvDNHjnujoOyd7mDI1gLgYfagNcsEKnwGuWMesUYw278JKlsnrJgQiZjiNKfZ8
4KBRRncvksXdq7pthjhBmz/vKT1yspVpij3BjKsvZLzaxcMu+T5OllC1nk+oJ7R3mS5AeWEp6FDa
wrhgSjAExfW+fLG/yTUfmLApN/AZW58AROSBVIMZBtijneC1rzbJcs/WeGyCMkGMCbCloKFeufjy
bLF5pxcG/irHJTjLQXUjFXDC8vT3kQjz9D1A/jbD1DYrs5367SEIArg26hN/lzvtrukdsYiuKdK1
ML/qbDNlaNm7Im7fogfkeayIuA/S4e0Kp/lfsr28U3PIy3tr6uPOSTbfidnmywbRV0BX/7Q/6n3e
Lrooo+OKB2k8UZ23MM0kWoN/UN2JtBWI3Ge8+60A+TSDOkHJd9VOHFd6N81t0Z9f15Xim2n3Ws+h
E71Z9JupPPYcLiYzPRcuazmh2q3wRKEHRJPCwf3pqtBNcQilEP051ep4nGRllt4bq5ucw1AJ3oCG
0Du91BWTqFwN7pGqnuPX4YjGt8kxEPg/OjlA+3O1YnGCmsAeZJlZ3U8rGB8fGDUoojWXrhGvSuJ0
4k9ZPphZbpjcQAlbVgtNBZqhLewqY35B5sAtRsTdOiv7l55JXRRRqjm0Rl/ZR2Em0WXdFvNNDQz1
gVNCH1C2UxCZmPzzxp2DoZcNsvZIM8fAFdgCl27rt5ZXTM9WYWInxbdBGVd0pgYm8yOUWFa1Lw2W
SusfBworBICboYxIVXdUnDa9JhmMZRTJeuGaW000J/DF+KU64b3tudM+QTgE4iLC9S+3xIy0Pwaf
EswUaPUDTQTVTUPMoK6XoBK8PTQksw0Tdm9qlKPlOMERhNhOd7x77LIqhQEKWvCJxZ+fLctjTkbU
f1icZdWLhZL70Zne88BQ2++/GFkUS6gLIn/4ujNe0GBnWRAsDrn5SWL02ZyM3tnu+/exsSm6TAKt
iF/BaEjo/sI27ROqKnnZsA0igvzhFW7HkcNCvO83kh7G39gM/YzHeYOtQOASLbkqXyeDsBgkc979
SkfqGmspog0ViiT9oK9sj574Sp/Ime6yfWwpZbZa+UYIQ8AhyWdn2Pogs6kNy9uMDjAq2w0C08gP
T/rS9WB/+2EuD9KzmG96ollhI/gaU/UUQosdxqj9Z2GRmVlxNm0e6EK25qbumj8oy9ehbGI2r6XQ
OyCzRMBLtfzR3484rq95fnEJ26XyMVkuH21tWzuhMP5fggmmVMEigPZ1sLIIQOty25ghs/P+nFJh
tb+uzzO1/EJoSy2RwDNAbq/SqoDn6RVVRLfIDZiJdDLzddjbE/ysNMenoBDY/NzOrhtUpwmxaieG
4iDhBDvXkDUdk1/5zBGzD4+gbWz01ikt1KErxJ/1Gqc/fb2Az+NCdG4VkPbdZNTOTlSS9ItGCreZ
XllUFSyGnitifmmyKhZkb8ZtZHnz9I4Qr6YEEgUiCFEi8MuqNa4X2+t/w2nosiSh7DVVlMEBFwBd
9mUtSNTf91+mZH6Uuled04gJA+MdfACtbIyK0HtqiEX32LVk/bGDLJ50ohUNXD30chonUyEuhvi5
XdCWHGJvaTtnrFNQ+2Nn7uaegEtFYvfkFrHS0cZab6DJls+VFSJg3EPZTfth48mbfbxtAnn9Kzlo
Y+nTTzFuHDGMesoUUmTin4hSqiFUni6OzHbspm5j1qtr+ml+bTMgJ/9be8h7qaHl8QAlvoD+uCLI
dp2IqegGU4Fws7BugbNnqjDSplk2CNkb1IxMDl2ufEiYZ7RqK/nOSHNFhrRCyXpJQI2j2y4YcDFo
4bOlE65oTTGLjI3KZvf04A2cvoQfFfAk0kavSehD6/E3SKj5LOnxUGYnAMMPQVu24Rr0OL1Jufil
vk9bvJ7kM/C4DVejVDnbYJIfrpuG+uEIpfnzypDuSDUHsoUNLDCaT8QKwSSYg0lbo4CnsM/RY3qB
KyLlQL0S7AorJLwfJWywod1Q3s2lUsoSoMNoL+CNcDq9t3WiqqwWEMfsbe8L+/+HTG14oCvb4usw
lS+6IsOToXPZlLO3+EKRJjpf7g17cjMkC5y9cNaJtzOoMuaJO6hYd1rNuUsktkvVpHqUOPbt4Rg/
aGazk2SGYSnc1JC80qx+XffF7zellG6l8PrHrAqy596dydU7Y5jRFi0d1x2uvYiLEoWJq15L07xO
oK0h2cNXOm4Ae1O1YJq6NSOGwUOZaa3DpHw10LsFtEKXXARBJBTC0CvZomGvw91rcObFvv82qctn
t//fp7Ypj936bHrQYR4e4eBYjoL7vWckSJtRktfZtCcxe2RqDFsjZ7x6ETvBxUTmBkKderB1FV0i
useYchrwplWN60vwB+cDncRRzUL9xEKZdRVYW9jigI8N2yxLxJAUjOnlLGSKs5Ke97Lukr++H144
ru1cIYqNGOyxXfHbdJi8mHuhR9qnfrrjaui45tIFftpHl1hjskTMBQ2m5vqINpt2i095350O1DCT
cCXWB+ZVxqF9yPJR0Da+gx53Wt4eyf2eZZdxNmOw32SeqP385d1dKIzc7yrNXxUHlmV2zba121oD
fEG9nBY1kI36QfrexM85N5fJhY/LIVcMApHWMmYBODUT9kIvMEChgn41NjzISx3IzG6My991sNf7
wxA6NilkbClAY9wgQIe/EfxqnZg0rkZcNXK7DoY8mh2bUJlf+biBT7Gz++unAvllT3Z32VgCpXwi
n8QKbpcrK62O4Ol6VCdUAbCwBBORICC4D5zFx0pH+dImvl9pz/IZIjyNvzTSpYpnVP/9fU+zXaK7
iPz3aA4c8UsCCLZYFlgq6pDLIXg2PesUsYevOwKdKWAIKioOueea0voZG71dPbMBbtjYHRTb26Iz
8WQyHVQ90hpTosUSuWOenoIlJTnDmB51FZVQHxUROPSVyNGiY69fW/WyD6V//bXlUaT4CKmQkjxp
HQJ4KabthqsBh9VMTLIvR2BUXeYfixSZ5Y/UysVexjxnreRZbo4gD7dcR0eyo5i+m/pXrs6Qv6iX
OzYy7UJmVuocQbBIjIjv+dK/elT9zWRbMrNljMQLC843GwEv7YPsFbrBUJSrUDK1WLerTOZrLWsX
fWUhuWLRl15FvUIXYYNMZ9niVF2/fyyMwROsu553sCpKdE7g5ft0Zbu+XpTKNcsWd0OpXO58IFri
SWnw5MrHLVIF20Orpu1PoYVVBp8WSQusDIXFtvO66tnWay9Vf5pol1aqRMW8sbhVQoqEQZMFS6LU
O2op4YwBB+tZneuExR0ZXslkbdscwfj9OeRVXigkJft36H47bkdocmSI85hw3eKOotkCCN61mS89
qpOfALGJxmzrtX31UvH8iCANdQnDQsg+di7x61gAyvHaALCkA6GeyTMrej1t3PhLtijwa3OZ1L+Y
0R0RSTLq2qw4sHZ5TtwtMAmxOZW7P5kpwUTPhy6Cm7KdshtXE2Z8LqjK8j0ineYV/OuPWOfm0O+1
tVdxdHzPNw6srDu5x4mMlYZUlQzVVjrzs+LMCff9MB8g2xTJeeorct1MmmUHF1Rpwg6Yw3J+lEBf
m74UYmFnQ5XHEByEdx+EkcCAPiENUwnK1StT3LNoz1Ee90kspq4H3IJBbcHG+qhZRgZXjkNoTyBQ
BFpueIk/+XUl5reb95M23iGv7Woz+Dwxej9Gk9TQiohjWI5Ck4nb3ZirRzz9TSCtbaT5ZL8B/iiT
tWNfIFPiLn1l86EWgnriDQtUQ7G9u8nwKsQe7lVls4MJObkD8K02cd4OSHWevulhEFmsmIcp++9X
dP37fIJdMlhylqa2zM+YLFBjEC5rltazaH4i5x5n5R1zBQaADl9zFUXTM/TYH9V/YUxIBBTMt6Iu
Wgpp22O8EEhf1LZ/br8IqjzTDg2vv1+WAiegaVXu3PcGPXIx4xEzOOApVyVeKNrcffxyZnmQUgfr
sPgBJkbf/QkrX5SIVo7/uYX+kBK9ZqJKvvNcwy9SuRS493XRa2T2kBCQ72b3KZfZXmTOnBy/oeSP
Xco9yhMGzf7G9SvuOj/rKjsN3tAbRPjFxYruC46UIhA8ueOF1TUEQfN9+c43i1Jm7jM0zGkl7SZc
6/TELSoe1jNoikHLmSRKqmRPOiorn5xBxeBQEZJ2nOxiN6Azj6gbEZIvnjii1fiqBXNBzwid/eX2
53yM1FSNbJx2MlQ3FirldTI/CEh0s2Lx7AO6xVSS2x3h/n34NIsfG8I9UmlFMAK9VGCY1jtBL7we
zFsnZebl/vAnPsF52dy3OT/NnkOKca7cV+uMCmKlI808ZKCvIi6IvyWiHDKWOhXT19VNb+pur9xz
FHkl+VAp+pULKHVvcDypv01/AfcbCNVcr+yH7McJmGjPk5R9eVg8faRj1drMwgSt0rnopzLv3i5k
gRjAmyiyjVrxw6S+5L7KHoexYVhFaDfUWxB4hFX3iH4gZiYZ9XBHubUTi9DoSBYY75KzF5gwg4Xu
fsSpxlPA/Hw9TR7oWuVX71Bfpezd5PsHbpyNMc91TWjqSAKFtwdZNP5kygU1CcUjj2AfhLSvfiUg
5inM+HUkPFvB3b95J/YI6FDBIqSn5y2mU/8xhwwlVjo94OwHOONozDjiGCscsSmxP8ZU3yEu5/9Q
jVd1lveCx6EwXMh2idwTJ2tg8fDmXHHA3Fz54cy1kvwXyrQpok+IdXU1j1v05XibZEhjRYOj2Mrb
+fx4RQ79z5LPw+TPrBRPC90ObC3FTNTq6DZKC44nVJ+y20iNemxsrSIUXHP5qXcsXS82WRVOpyaE
v84Fu0Nvxc9M0KDYPkpMWD3EdUaKSm6VYVTfMkILJ1fK0j56AC02bSE9CAPj3t4xyskck0cPPDHV
hGjLFBErSRrtvFQczidbc0hl3YHbx0+SBgkis/WMcP+Zltl+JpUdNhba0VLj6nMrOAHepdB674XK
Yg+83Z3VCjfv33MPuzlqLuVZQpOVjD7fL+aQwfj+zRLPaE7ARWmUgBsKTGg2BnUgNUrM3veZZN6C
eJOVW8ihZHIsj5naq84FvBRKWqIIZcim+2wGuzMBSX4OBCxQSC1lGmOqzP00D+PsqfqMGOlOukHy
zVIhplugPyzOOVimgCkOkV1KMPAeuFZODzFOIOBhWH8oca5pkvwzoTl7TjnCe9QWdT7F6Xn9+B4q
7KwDpugzI/cTpMr8lQUINCPWhD0Gazi5M99gQHXJ1nM406X3L46H4OmnRhuthAXoZucKB2WrooPd
+dBQpHe9QM8ggYej4lLtO09xrRtmbbc9LfQAHDKrrraddMkcfa+NFYb59NCHIqqyfhmOYAf0teCO
PK0P22jyK+j2SjaaxVKAs+K9BCCB7nQY5XpYg7PSFseUTjVyZw/36/M532BFocyACQ0m+fIEYiDP
C4epF4TuUvbwvD8vNCb/RA1Vys9B6Yq/hudvHkl0RYqHjsoyYeTAtqLLWCErdYQ2UHJ6ge6GBWqv
KuUDbyz8uoqJ8+mWpgH64z20Qxfzx9ehzBflV4xZNng7a3Mur1Yl7Ui5EMdfDnm9xY84cl73Gh2a
NoSwrbD/GaKpQPiKorQVVMs4U5TKB8pBubRy8Jf8DuUPjIfiOjI3pWKz0mcNUfdSdk1p1bbx66Hu
xc7mQ68QUVn8WuVjRNvgJNiJTP8b7eEpE48SQvn9gwg+1dIp7/Fbk274W44AKxrES4Ec9FDZE/46
Jg9LtlG/1yn38GbS4otoytYh7HIyJlTfoMk5ZDR7SYfmsWa6svwMcRGXt/ho+Ixtgqch3z5VsFcE
CeVgW1TePdq4Hmk2LylxT1hyOlcU2aNx0rtZS+aLUeQ4UNdkiFCifZyuU5hex7/6i9OOVpPaZ5S6
Z8IE051ALUK0cHmD2cbqc+txFKXQxHltIz+AWyV0+3JOTmn3UcLjYOgEAw8hLViRXMyHKqka12I/
Y6t15zdbz1JFWQOl+F713lqpbod4fXuG52LMWtPvGb+YKgNXrhAP2KsRNudhOIZzq1C3hkVcBXnj
YN0+yD4vNwv3NA1r/5n2nGJHm0Cs9XDhKSz6xC7YgeLBkvajOIl6znzNMzemb2cXI5P02CAvZP3s
F6KwNlLxHuxwBO+T/B8IFXznFwagCYIqxIHP00F26s9FY71HwPM/0R3ATQyrlAEi2FXVh1C/4WC9
Ty0oI/PrNw1Ia7vZaCm6iRTVm0C23+fQpobGjyFQK7XGHDkVK/aK55LiDKSOzXWXTE8wNoZCGyLv
tnbER/zGf2FN7qA+uhXRUQ+auxSB8w8aV34O3D+3Zfs783Y4SQhCtA8nZ1OLOMCpJT2bqfwa9VNr
sS2TkaEguSsRfcxZlfrHhG9mH5T6p8IARTV3ZvnxhTulgWHiXv7cwVNPtZwQdsl8wQLg3MBBrdyE
b+l8+C+wcKrh4dMsWUKDP55QQlCfJlma41qzIdA3l4MjO8VpC2tGBA4JSbSf+Hc1wtDXFZihCvB9
Ggva2NPc5rlr+WLIrcBZydpNTA+YR/0ubcZU+zEHodaa19IzAVWHt/hvg4LIS0ZT7tcgzYMojybI
ddQOMhqQDiJu1R8j6AM2Dt5z9o4dH8woyqMRK3NAIqTBXzyWpm4MQaH6zWXjVAWBliKlZDIyXQwT
x7a+EVuu1UCVM+7UjntyNdcpIguSDIR5om6ecHuHZLnZ89pQY9p9liGPF2Xew2BSkluN6Myfkj1j
6y0V2aWkROtTIbxk62+vL/M48VfMcEJn59hUCWV7lrNmsTdrxU6CWpVdkRm4VRsAPKS2H8rOuD97
l31zKxwbhOc2ZsaZP++btzM6l/em85D1lqFFjPVyMZZrdQMWFo/w38OiM0ASB1AvgZQvzRNXd/mJ
7mZqVISHDXxdcQnOgyIfQI7dbm5YD3UxHEI8IEkO+AI74PZhbIzvFvXbSCru5yNNR2l+Zjm+M65P
urPZ1rQXFyD/8FL/EmUYn0DLabISpkTB+AtO76Ofh/ZlRF0dFsh7C4KVNnNMzyqjttIvXe/SKyZY
/oPTNl9xAXgyAIMQk+hAy+VkVG6HxlJHhplKHBUXJ5sLq4uJGzeSh7RG6nbd5DLUoPCQ6JaB6uJN
y1lI0v0T4rBe7OQFuXNpG39/Z9C5fDDUTxbphc/0PxJKHwCFEu+N1RkCmHBK9LcDVJ9XGRU9sGf+
yBgrAoEKg9F/xqW/UhFFXKSId+svJzr4V/7G7sjjA95JUGRWXDtd6igM/raYrx753flSWyzL9UoX
wF7tQkC6ox/sWvgL9n/qOpudDJZh307xcnqYNNdrREjf5N1YkF5dYxdb5s92JSBGNzt9hLdUWWKl
+5W6gH8h11tQX1196x0BUPcB4EEQwKY6CnOqvGBzJ57ykx8m7tuOX7wu4wi531s7tM/0Xv+gYMB+
GskfDR9fVg61SEnj4Cww6rub76u7YDa4jOPbsGBJBwurk+L2rKueEf6+CX9jjs4EaQsioGlY7Tax
kejw1S0sqL9+89YII1wKf3mh37k90HhG8NF0vM0nBqG15ngziWn11EGMPGK4j/A1okZmiprdGi1j
PqkUIHr5jFyRHvZKPCcNoysF7aJSELUCSjPBr+J1K9uMfqjr7U21A9/Ek94uU28LlKYe0Jp8HE0R
GQQpsKq9QzcoYl/FqLwFeNeTS4/0losBewWSXmgdima8ZLjjXuLloV8rsTQNJYRJd6BuM4IBJrrr
Gc4TxzE6xreIl0OOCipxlmLAUFZzW2w0Ca7ESTZMcr7tpu33NLIbMUKQPOpzymnDhqWqco60/ooU
LzrtAmR0icowZJTKCsTsiDYbF4Tu3tsO7Z41h5L8adpbIRo9Ofx4XH9g40tdvQb3d61R1GBZ61az
b1hKm6yHjBuJ5QeDJwlcqqdhWGcCa+51f2wMK2quaPZmHvI6CyWV+77nGH2cHPFG+TNqP6sZIWaf
iKK9vu7wPsPeYVqJONYvnHHOt9k2E2SpGlfOwfso7WTY3PUvCP0jMQUrZtEVOu2VHHx3YXW9Rhpp
CbooKYPw5tgCGQ73NYBKFaPEYTd2zkqXu2lr0HoY7+oe7mByLO58wQg7Fe2h8GAOb714SeJaXHfR
Pjr5OFS08HgaG+5o4n1b9DdA19dF4csuyNSpnBDFeIVKDjj4LxLJl95tI1c8ZccwyqxquvGs7EX6
b0qP8Z6lyO1YQerRW2P7aFVr5VpF/gjpO319HjjElxvCC23qJPS3p5yERIRZfNxAW5hXDoMwUA1M
iV2RzOw0NLkC/HCo4sqyJAZXyoaux6kTBy2/KZGlqRUvVGAP78bafJEeeoWX+/tHPxFUxqgo/T0E
mr7foF+WVjby2mHHvtn32/CZElUc2FXgd+9wUN/r/sNsHIQmiGgkx5+Oppc6RPIGxFj3QUhwMyFr
LEBnuhc2eAoAfc5/mP1D7h4JmMoupdMbyXSsH1FNUP+aVeMkxhSQQ3haK/UU2xUZTY3GRciB4a1s
cBEfB35Nje9asVhKzGcnUQmHotqSZvpHNnlGTAUQ0zRjZRbUig3nrE+Xy6MxzuPXWFWjeAwGdico
0/yCu6NPHRU/HEld9Is9ouh7F9Bf8fEkzYF9LoePzbkJgkDTNR+nTFtyEJRDQnkU24z/HrGZlX6S
aiEoppQIFd4f/+MrKxJAqPKaM350cHo2Rjdsy4GLBdadD06vZixdZWJpi21M+vvbHDQ2CulL9S7F
IsAZj7mUZ4FqyAYshbvK6/iFe1nebhhFbllrRx5BEY9CzZ/vv4ocgIqfkXnCIkUuq5/qFa/PZxh7
1v2N4wLAH1xaGl8r0JaVaGG9u3iILwl+o3v8IHC2Zs9mvQPg+gJRP/fWpfjIGpaRbknvrsGJOOa1
nPDdLzW9nzBeLchFf9Uykr1wZcu/Rjxg0T3l50aGucCFoNIYyMJ4qTP5AKoxS/2UpJcfMi0J69LM
zGmq5D1EBFSzpmVcNq8GnRyCaeMPBkHXw/oTeFZVxsP3hZoYItM7DdOyUh/xHK99ElftBHtudom1
PDoqqfc41juEQ4IThVNd4J1Bo8qVTO+KTStQVN6lxCxkxW2u5IFOYEWdijR5job3v5yNDYeH1Jhg
cm3VCaOlQYZCMJmJptxGU07ff1YzH117HQFEVWBKi1QX+OsrtszK0jzcjyJFoJxtXy/2TjdbUwKH
bOoeW6DEAM4426SwaQWDLQ+C0MPpWJRkSk2ku4mCM2uji7/C0sFArx+Q9f2Uyx1XFWM8O6RdR1Y1
JCOnRAs9D8MQ43E8Kpjza1d3ZtUxZ60gz71OQ+pgsa/B8+HAoBs6STCHwts9kQ227yWji4am7TiM
ANg35DMnx6urTQZutozV4Oi4yhOOYwi1Lqkf6VYDmSB4K5PFduYvJh01/WKAnMCgIp6uxvfagWPo
bDSkVq3Pd5Vl7OxZno/sx5BZUVoLMfpGxlXPpfDLnmBrtoOmGpoOKqA3hvpNLHZWoxQ7qjYZj7NT
9aXuIbyITxXhJh5+go/9Q1731lt6CoDzKYeNqLa4Mp1rg4MGjfk0rlTsSQXUw5FGvA/2MxVeoiYI
rmYpBJRyBgYRXw4tSgBk06CowR5E/v+VL18BgW5iySp+QRYQ6KuVSwN6QbgbHctyovO3LX2kntAz
gy1FUY6o2vOloYkAuzvVDLO6w1pMinX9a6Afp8ivYXepK++U9quL+s6EkkJ/J3M8EiSLe3aGCUf5
xDovEuZi3v6pZ4/XObFJV0CHQ8trAodra9HDQbxeKxctihyv0CSNlfuzOf+V3lL0t+Ov8aqqxteE
LiZuF0T+vjTIS14+uu5bh71Y6YPpJcxrV3FKuFxZGmERpluHzMBVQo46MZ/4CRq0JXXZY7l7Sv2z
F2LxVJR6mTtyXrBBye510+C0ptxM3n7NeopX+5Nk8bOVgdfaLTGKdqRcLKEqDG/AwA3buw8u85wa
iUtkmcHT24HOPHGrrPqDU+KjFwBNOCYffA0zQqglDl16lYYRjK09lzzyRr6KdkcVjR0lwlrh+Hvi
yVsJjz2L/fc2xGHkFs59aptl9Jn/pR6cTlPcRwNae0/YA6Ym03WWCI8iC2mP5DiG6/mk6F8Qvy+Q
pmt/vZgNkv0O/h8VVb1i8HIXfnGb2uOxjXTpA9Kcubb7kubYiX/ILhm/oapLunfQFBqPm5SbRfbT
UuwGMkD4j05oOZMVpiNliOuDvBNxbIMO+R0OhRK+Refr0fSYhm8WLidZ+87OLrru9AK6SL0Mo6vH
3pTdpbhXKdLRmokf9Tc9L7T4x8S+WOxM0dptfye1cr2wSe7gkvOqzN7BlexuSzlIxic4jw4QY98T
vJKWuk/YLA7MwM1c7X80efNbPLkcXIP4TYDrDa4/Jg914gevQ9Zw4B422GgkyE+HJmAc0AscpQtM
eDFi42upS5gM/NY16+T22yW2fhWWmhA6349EpkfkmWd8P0Kzhxqh05Zd0hDsioNhE2VJn1LqqHcK
tsTn+4xM72SrB8HTofv5ZuLfZvoma+UWQ4XDE0pG0Jo1uvLoYPWrfIa9pnbtihrg5PvVKPOOfKJA
U9LRFTdWnPJGt+WUFMmcBzK2gh2Ir7RWAFfE9zATUyZ7VJ8jxzfrcWTCIFNw/zGryLtSFHWLiZyh
Ttt1EtmcRi6+CcMi8PcryZ5ZwGlvxNMfg4YBSR3JKW1juo4ij1AUGtpumjO+EoFB8tRQUXMYbu72
bWdU6Rfu+qIxVRKyxH5rqaVuXgUNc2gpOkRkPRYoZvXItUVzTNP0as2/Hn0VcGaOG3B2w7L3r6RS
y6p4tZS4aMu0WkzS0sCn5hecOyukukRgKDmJDYSPcAYC7TwNvWmK4V1+pbX69Bn0/jb4gWb8ddwh
zsCiuZQD3xlYo96c3/NJfwQO4IO4RbppN/jVcSp9wZ3r08EsEiJKAs8eUyk1jPwl0QpeRusB4HvL
U8l9Vs8F3VawskOX78Eq4OED90bxWkZhgURC+C6dOLJAwrjxFnyraV1q1RDU5b35qEiAQOhXfWq8
HRJnqiOpN+BxLtDZtK112BoCAfz7e5tE34SAuKxabaPVfw72BlquswMVjaIhQK6Uhvy55+k+9rkQ
bT3AzeJGBY2MNdiIc70dWH4A5Hsy6hc+VRA/g/YF/izeAXANc/BphrqA+1yE6IG0FAQpbNsTnoKK
nT/OhZjUkyms6gaomqWi2gVXdGIz5xDcCGAwlwDvIfr9aXa/hILlMKTArIX9cNLgdjalyn+Czue9
GVZk8FfocaEE9+rpWeC8DLiifqJwp36x4w0Sgx4UQNqp/GIlZ9aL6Zz0zOewvZi5mBf9JZ+XY81o
D6SooBlaSRbRJYslEKKVikLzsFLQ0Td1aCCdZ8g43weWOnRj3+HbVFyy+arB95y9v6VhJLrxTkd6
zFzOBZijIrLpok8CCwZ1j79iil6HUDhsHOmjvsg4s5L5kXRx+j1Tp0U6jonKtlrt2rrxY6d3sZ91
+39XTqP0jLe1xKlyyZS42twdBW2sCa9nmtHl0DplurkjQQ6A9aFzgeEtyDkKDVTo9zarJE4cWL31
g+gBqaLIauIVHlt+uyJ+ZDmkQN49XoXqtuQipJ1TGONzkrtdEoLM9Vf0hAoLrfbF9DxzAqTtX5Jr
HijKU4BeB6xA6LjTHgAHPFCWunqD2CfeOwqApxzPnOCRbnujaDsdr0NQ4xHfpoGHnOFCmQSWk/mU
36LGjkCd34uNdsoDF7l1yzZXTBSSD/iMQoTkPku8jdsi71qYqOT+TlEtrDYhRONKQ3y7AjYV27RX
S3TbtHM/GCBXXNOPFzGeDcjdlJFU3srWi/9OhG4ac98+xziEldMrGU+8eeRF4tt/wAR+LLT0M3nj
Ln2Il29tHs18GcuN+Lm1kwR9KEmtwNpS/lp+2vx5E3w4LUA3Dq1/NdCVYEU7EF4aCEOlMuslze+7
eZWFy4nWK76G5Rosc+ertaQDP+KpqVmpQi3hE98vliNhDhJqrsVUGTPIHqozfusaMy0e72WRd9No
tcFJlim25KVpGdTqA1o/ujnc0FZEy5LHeh3c523+2CeZfWy7PpJldqnxJOozFyIymXCcHftvntYk
3+5mjKGqW+bucDS/unqDwNthqgHybkyjCGC9Pz0Bsfa33oyDAu6sRWQ3JAMglMpRViwLGtkajoFp
A/OHnbKHPkcmWEndZrVpvxlyzmAsoQUu7ZZIMdXJAfkOe5BTmzXErSV0vfNPCqR3eZfwthrRCD/I
9/7c8OZ8T8nC4M6z1Rsu6gY/Ug8sceh7AwGyrXgXOJzCFrEoZGLVwVcqNG0uI3E+WpnB3RVclbFQ
N9uHsJu6ke7iwMm36fsZ81Ljkm6/kQrmvZF4Chp2hqka9+8qrtO31xHMdQi+LYwLNAP3BN9v5Iqh
w0gFXyxB2rdjP5l1jSxXVI/ze7FN1AuuZgmTWB+h4I3TtUmZs1Et10nibghmOsT44fI833ye1t6x
VSCVGM9xKN5BtlX7SVfTj2x+poeEnRXFOfJi954KESJT/7EkLxpsD6+ssbbMKhLr+w04tyk/l1cd
4biGzJghGYn2Q/OwG+rGM7C8OE0EuL2AldCls+ZnWtWeKqd8hc4PkAGMUD5b5Ls31HQ1TZndwiH8
R9mVhCA/doOanZfU5z5CPzC4NkQuIVjeLWzXatIukk+vkyCla8O2f2H8NAXPopSN+tF3l1gn2V0B
EWfbUEryZV4Gs4Qzy4wWRScAbNuBSaHYkWLPzEn2SQLqaZ+c0LUvf45m6uml0wXd7hS/TXA1zlJM
9JRG+tandLk+m+nzxs6x7ZHIBGsUCaVll/apsxndDmjcZfmvfp/vxN6sFSkFnVu6UsAmxifUU0TK
0wDRtIV2EXaGTEU9vsXiZHt0NHd04zZXvl+Ju+v8NJ9FmIg+LckRcltwawTD5Ga3SWM94NGSb4rP
Cc7GbpdPBl8yxqDdTqoVOWVbcvW19Q6wJUn+mDiDOYwkRiPkZ5rnXU1n/kyv7hoLCYAdtpfH1m7e
oz+1qhlegqKsFkOfINIlXtsc7XmVnYrYCctCGNwqIwDolOTSA7qt4sgDHWOpyHoVBPAVuFopil8f
9uZwgrTecUAgfKhWiYhZn2aD0S7q25cVKjWKGctXSUCihqLWzxxtdGPjOSOmUSKcjRvdcjpYj5bd
b6A+nOgbzYd9XqDDPHOv04LA53g8z+iCN5qjpTqsNfmJnJv8cQmi4/V2yM4GxAZScO4P1o8xq5XD
w38Kh0Rr+m0G4K5TecCEf2znewzDdqwfk19yr28bbkVNKPiss7UvzLNMlAwsz6GKWIgLu8cBEUtT
/dYVPDILqc4I8NXjbGiiz000rkbF0dLp63ekUcnFNBJuLcEF1XNSnK3WSKxR8GKcBuimct3Xxl7Q
ItgM+yo185yMmWg6OA+cWhlfeRNSsQ4DGrxMee3JMLddVuku4Dc5qPlk+KM/33Q0fpZTS6bcL+mk
QHRuAFD6UpPGPtB/adpA4FUYg1aM/dfs/j9DiAAWgyKawd3kZXd2Aq4GcwdBn0zFuudRPYH/nA5c
Xn+GyIqd+4KN4ebWKzJiEVKmn5FfnwT0JKzPQVB0fZsSCBeBsNfiym2BVNzeMjTwjcyh3W/P4hh9
BKkvH9PW8mfsKCoOACf4zJzeRBglu4ZOo6F0n/Gj/vY/67pSMBmiAiwyGP3uBgrec/FTgbkAjpsm
QfTmyQXb4jh4Eagde2NH8b8QqiM3JyHbmdDxCLuPxKivcrZq1L3cVFvZo2Adx/gdtzHvesVAWZhw
QGg3a+0QbPVnpCcFdQvrNqqsnLGsSVuNi3atVQ7Shhpci84ZOKD9E6O6Ml3vzbftLj2tbLueNXFH
8ojKSXIbHahlKSc5Q0gNOZEEdM0KkohFa0hnaP6rMm5nr4MVy2mvVSeK8HBqjyoUi21d/EmhggeN
Q+meukHQWftUi08DIdlrrohzkBkwqRJHRTDd8UFVLnXD1aVZviYgVBDC2H3XZwll4Dycke7Y4OeL
xzHt2qIdtPfe3ex5G/zMWJ1rtE/bJsQQADscYcwJI2sLYqXLxqOF1+IHcoH5zAAOENOXM10vgUse
RKc/UjiI1F2oCcKHk7mp2SR9YtEGvdIDmCkeIJr/IaCbKKgOnUEHgvGahh6tLD62eZl5kbtWAIIo
vo6xaAqRZoCliYdpYr9GwZb6moi/vU5YoAJElAYeVF+g0qcQPNA0YvQRBcugAphEA86KuaxrtKG5
SWk4HuVyhiBf7s0eG04ixWMvZsJbcy1Iqhm2EyHhGmw4fsm535sWeNzhlTK2uf6oW+4x0GVhmBCs
OXk/MHyiIqSVhWXhRPKDLTR//eihB/8C/gf+DSMeLE7yUmsdTviNB1GHW+A53N+AGRG9SMqqa5jW
4AF3ljPk2JJWD63JIcWtI78Um9Eka0uIpVPiQ4svlPEruG45qY+c3UOiJd5LHVlLjhoym1AmJqkp
GAj92WMULdT7wL5tMEBZUiv8A3JXKnPNvL/RcMJJbStPSXEX0QwEVUUqzGYFVkxzS//LXL8ziMfV
IOKuyruIwHnrSEdqlaA1IYOYX+Z4G+VXglyMBKdMAKBLY8ZnxtgPgKnI2InavBSjsxDU8sLUKtZ+
1uxhOtPE/Sej+eGu01V33X8Zda702baChunqxRbUjAx33bDKFwF3Qv+JedICS6DZ1fi3B3+XoS9z
SwOlXOnOuK7ZT2dT00MocDFR/vMYeBpdpXZnCpxaclePCBGrLGvw20ijOcxAyM/DG6YuWB1sLktT
bgWivxOLDn4gbeLaDSSDTMrOO8S4F4pEyEI+BzPYyC92372i0/UavnbS0b5n2nfTT0Vg6YxSFwZ3
K/R2qY5Z8p2abkNOSxBzimXhN2C9IvvbMOujOqoWYCIt2USg3jU5SS5r2g/MiuRafhOEbCo6PK0i
HNgo0KsO8g3dJBIvONbZkNPNJorukHNhIzd5p4FgybYprSSkTZLIGLhb5oHVtAngRB+Gi8mac+YP
W05GdQkdxA2akzxXo2fZ9wI+8fXZOGWWJz7efjGKF9QIa0LC43L9FjimeF5Kj1/xPU82K7pejJJZ
JIk2ytMFO3tuxofXtIzTOf/1yChdXdsfh6SmI2SkBFy/S+Iay4nTyINH6nirHuS7WvKvYX5uMWNj
r8p3kzyV980/NJ4SS7hcPU1S+UadPlLAprMbbVsC2nSLsTsKHblXub6blM+4diPM2mRTfJf/GMvD
AU878u1N+5e/hjG2xFt/BuKO8KdbzIsZgKIv11NofyszwzBCPv9/dxUvMO0v7QfUDRnSPyYLQg+K
qv4zzXDYpEet3OWa7hqqoi5vTMTXtsQINvXNplykOyBUIGkyDmaa3d7x3RpoMOP7MT3lAi5aDdW0
K8UO8+sBY3ni75OvP9dX3zpsM2+JIUr3CVG6ilY8IGbiweQbI2HE2NF+MqW1QADzV4ldopit9CuT
lt2r60ROZ1TiEvggOxN/3EKvpNHXPlBeDZDiuhmd/iDOjdRaOHz/EeR42CRvnJwHWC+gNXUAAZt2
kafxlF918d+CJHOhcpS4aDjKoQ9VGvjvRfnKLl5dGQlgh4dDejRPy+wKK2/vAokd7PITgbcmbDLz
lD/NtlYVy+9VwLpMObSt098ERNm5pRxYs/LHWuLI4lC3iWTcUQyoWrDQSQJpj5I8oCwrMu0N7n0I
ETP2fA0QqxitfJm3FVluafMVoBxqgkjLiq2SMPJHjBtYDVcMfejlVDuyJUORiixhx8C6eR/mIXYG
FPLrUH77NfyrYxoB1Dow22XsyIjKzfOhfFBTQ98FtWnynrBe+j/jQwVBny0jglkfUQcENzoaSj5S
D1juOi7VsHYZgjT/Gd6oG5GbT/GAx88xL50g6WglIRq2bT9EKJN/r52Sw/UxB8ziQhAbsKoquixT
eZiJ70PmlV7S0ILKaQugzUqJElNQ4NKEnKqv+CEiG1YWB+mmzX5/ZDbQK4ke3RyIzMwqYGC//u5P
UD5rXMbXVLF8Ms2Fc8X8FHEEkG4Ifvrxf3pOWlw9faRS6Mhk7dlPToki1Feph4sqdVeioOulD5PK
36OFn209CxbSMEnTEVxsOiiIfJ9k26aYrC4V5plFz6umZZfQOnELbSsDXhJlMOQ3d7AtGRw4XSrO
hoZGkALJaqOwdCfWxZUZdKbD106tuY86NlCJWYde+t+3cu2pUoqzEIrozhWDq87uWRyISnfGZOBM
O6HNNMbzIM+kz8V3r3cfDUCgFmLHB0qcMjLLblSk6D6hNOy08p7e5O+SOccs0hZlvq0DKNnSYw+O
B+65MCU45tNfV3BhFhNQsT8vFuG7gw+xTay9/erMTXuy3CClTqSa8D+uDFAou2YGFgA+kNpQGg83
o83o50FPkVh+hv6q2oHSO6xUnLP0NMHKFv5rOfhH2ma1mJ9IZceVCqRel5vUL+ebXl7fdwGTepUk
+pSD4ZjDlEIS7Jbp7nS2XIK7d0RzCF/FhPcVQd8OqUylBB95tgR8R18afa7IhvbqwGNzKtSiZ50v
KrYBIEc9Bch4OsziDz0nT+PDiJqRGa+TvE58RRy9Ha3wvXRGv1k3vzrbnDV3MVKt3YlvdBkSQkkd
iVOkU4pVNE4F/B6JgLU+o2rnnX44Wq5kr65y2IF2VyzZ9vL6rKqq9j0H7Gg7IjEZfltuHML7u4Wg
0SLsO/Q1e/ySvFCbgvy9x9JtdVKCKzdAq53+ocOpDsCD48wlvv+AqxwE83JqbfsG6AnJXC4Km8pn
6wJIN7nSxCVlcQa9WL3ousCrKE5J0v4PjcBYjwwEhT2cjorTxqBHAKFLrTC0ffmfuKTSsfuXgQE/
qNoSWNo5FqABK4pRFaEP2Ypr/xIgSDHU+IA5BMOGpiB8+UsfkAxiaLlgSMwCKqZxqHshww364qGb
5c0wmY0HIBfyiBHVCBahCFJCJ/GwlfoSzrkGW6QOuRbWQgKuOlHce29nCl7j26Lez5sDd2EsrGPK
DnjNFUjyXXtxx+vVWiTZ8W8yirBu7uYLN335O2g/HmiHN71iGkn4FuL6AioQTJOVSRgPCQjhgXMP
/r4bXjxCuWLw+xbBsoAnYKfYIi5zQYysuEyZD6WCtTLImNHM+SQxR6+ZES+PxqGkUhN18I31OORc
65FDYolLBVbwS4TmWYjU3IbsYeis0clp1O2qtf2ped/fo72F5SzDFATXqYRZYbTN4BAG9aabnr/w
W7j0MVByXEZSDC9ZoJCb/YOVz7MIkwxTK8glUzQAgEBQoSx8Kr9dtHrBkymtddnKKThC3mjbWDwE
rxSXVRuBts9eKzwjvcZy400wGfjSjtgY8AM4la68w0GG7hEkkrwurh43+24EtEE63+QoUvMXQx47
/tB/neLG/y0BARfA5m6TMmGgfh+iO+HueyMSLc1AH0Qp+VgiWTBTA0fzDCenb3FQ0ZRgHEsWCevv
U9XZjlIDEaIrwXhWasyfrhmNCHWeEeMgMHNU8He2aEaQ46Ye2R4cBcn3CPBKmTjB6tWIcfOT2Vu0
t6q7gSchO2ozntvqfY+zV7XN/JgPX0QaQ5/0XCHaWh9eEDEnZK/jP3SnvfbXZlABHOl4pvdJlIps
WObBBdU9XfVHeYkiJhbBKCOo97RN/IQJL2daqtH4ExbN+oSY0UwkRDjA5BNePfxBRhFmyKxjkmHo
cQTS0uiNqh6uJ3GHzpCfD5MpCBDgCoCrTTL0h3IioqBtjWRzJbQktNkBpwUpCbyhVs5YLV/6ruJq
phRY4kpi6dUK/OqVPe9sM3NmehK380us3CnqtI4QpTyoV9vRK2XqXCEujhJM561igcAyR7e2tspt
Lch4AjANnjfg8IsQRg4v4FFUDSArgRUNHmj+F6tzj4G4+uIWdI3K/pPKWAzdgp8oa1NL8Eex9wu8
/NKgnWClXNLPuZg+NdNNYPJIOHaOCuY4vgOcdKdNaITnnQdfrU0Ff4m6TFLF/3SGyjIzSK0C4fO+
60M3PqLCtLMCdN/TYy7lTBnkV0m9NxmoTZ31QbKK3No95hFYDT3dhpYjQJdAN+djVHXmx43edNE/
sQqiBXIPeBBwva7hDO2K7kUjAw4HD+C1mY4+XH/R+8LXrtkad64GkmKTnC32gXVxA4l1k2VXDDYO
aX9c3+uo/d3PEmsaMJ7sOwhmXAWd+HXlmaKusWVhB2XMSAL5nSv/vqK87GI4teKvVtjlRHys6dsk
slCxgKbjz9L7oMfpkUNCcjMDoNGZrLeox8KYkcWk5hokjTcnUmW1BLrDFjYjZ+Nl0Df8mRoSqOj0
DjxyxuV+Qttamo1hIz1uyAD0XBbzRrZP6Y6Lur65nfdFUI2usNTeLdCiApLTXXxr2RxDGyEmNWC2
L/48YCRcGLxUCMzawt9DE7R5mdpag51SUq6MbyeDP51ok1VHRHUPMUQh30D84RfT4qAGAY2tfdjS
bKftnxgE4T8bux2JMIuB6QWBrVd2ZqvfMHXbwBrk+ygrfgWBQA3mzPiKM/kyGE5BINOW5IqONdW7
YNbjgg7XVdcq7dbVFsUuPjSxi2DoIJiG2P8lKH1T+ank/kvBW3l8A0niLVykHaDuztGqJiHbzsjx
G0eelmot/so7PRm9VoZR5WJywUqCsOBFVRIJ3iimP7eFn1DP4nnJlnSqA0FXF/sPeJuRorq4zQ3d
r2PEk2+EoaszYmfMyniYms88wnpprUspcTSUer/ohgAkg6njOoDpHfXWIxqHYp2VYnChpXhF7VIj
VoUvUQeTAmoVfMInbNe41IH46m7CDGF2inumUINDTXpbpjwbQezi8LKLe6uUGf+r/iFhW9POmIkx
MBuV526tP+ovMaiJ/mc8Jd9zYh10i0Y3D471iyZX/u1RsILFeVootCxl3uLmVS5u8CYsfovHSzOP
nVAbWOpoBLXz4Q/CeLBqIKQ/fz4R/BfWXeCA6bbNMklN+kY0aJuctHNAjnhI7iTeVMoFuvxZQuSh
MFf4EuuWATWfwTlVX8oYWu08RuyYZYu40dWbeYMtZbfJHX08NOV8kGpN4YORv1wYUflBceruWWsK
VD41PiDL8egyAFOgySj4q6MyymMu/DAEsFMdVlAUS5iFwox8tvgcKiAHM+n2e2SB965XePoawsAo
w1UMUnehjCMGozVUAYxClnOQQdl4nYBbKZNxOutA56NXBPVL+xfkYpLf1X2KipzfYp/AuWEXjpGS
gFHYS8ebobd7nfVJs0gQowF1UwsYhTbyw6UCG/ZVyzVnNLD25ZMOBS0RN/3FxK3YJ7UK3MLogfl1
3HcqOWiwE6Fqx+K26YVohSfL6+GeTh+VR6Gqw7XgiHi4ZVf4tN4wUoBN1dL9WlDnzjru0iPI1TqJ
jXIaj+klaQcEGFdCdiaa8u54KQBLTaxH6gRTjJQdAACO2OrPOVm0Gd1Mu5L3pUPseqBwLNiifb+c
QaPm4hvMUz9Nh15gkLn9tvixB5ye/soYwmM2SEgh5V0qfWjROXB8XJWotDth4fumkXHZW5n3mu1n
HfXR4w2T2zVHESGH2f9xy6OVVRFIOQ30A5DLBcf1HbFaoWR1UDl1WRPgptTD7pmokBbg7GuJWEKK
w9EXOiqM32UtnLhvy4XuXPr9wudgz96tRQLEeGNbYTI3JxDNDWT7fb00uJBh521UY6rB6udKEiMY
lJz3Fe5u6L/36locHN1MmZ4obrWIpDZdAlYrGYo2/fpmlOISHp7Z0610xkJLe4I4gZCsjLsHPNYL
Nu3c8yPxxKRrb7083NEOikYk9jCVVuG2tOFWESnw0RlUz4D6KTAsNVpxKGB0JJkwiRjcc8ybR0vu
1WaNTrxNOWrpF/lBHWHQrlo7M0vkNvid5lmN2gEwvscTXj1CFZvtCKheesoBUnsZ9/1o5ffD4gsB
yCT6wi/WGUvc1ZpfG/q43kV33cPG3cGYFH6blSrZsusg9/iwEWuOMUrVaSzrr9eiUE+wJaWdc4jD
fh+RQQaXqFjuV1bY6v7Z0FU2XDprvYTNFVYYZ7fX5OgRQuL9j6wP68sQsi4bcBhQGGBaRplsvByk
Kwv5WKXSgaq/YwlSwDhP9hIcnFEn3Q59t2QgPDNPBOnwMVim9bbhqmAEgDoYto4iKFfubkPC/ySq
fonAQBI7Ich7xD60BPsuQU3MVpbli3Eg7hzqPasU1AuorCUWhYcSfjx/Iy0sx2CCdSCd2hoXkfST
NPypoJ1pRFM5PcpXqIigundD5qb4SwVNkGOeWM6wZYmOwd1tX2+RHbizfgrahA7Pjl/+JG4bpfck
RAeFlW/pQfSzsE33D0Ia9MMWMnF2KcWWpwu3sdAGwn1Jz2JMmIAoIGCPzlc581L+mSuWeYtN87E1
DRdqXtuC6v7HKChU96LCEBeiwhem1FWCNT7N8KLwtYkR28l9iRAg+sLrUl7y7CuCRCWKCShmk6MM
Zw/wrvSARhJ70KMQchj1OD/2Jpu+M3UZBtwTJRRKYK05HtcLnli7hgrNjSV72o52x989jVKI6sxQ
/Z8eD7OyIUSVXgtMmCjzBg1lQ5RLyN4M7cVCrrIH5tQRcZFqlIS8dGBjITR2guRh/TYICtuhexov
/w99cG+9XzOknOUNTA6cDmScc4M31dlImRvsniELJW2yRz5z4g1diZ/RDPDKHYmHXoA8nZCpZQyQ
cGAlYes0foPheBcYDOn9V/xBowFG8rZ6gMgw8GBcqbCh64MxvAQez0KkjBzM4IFg9jhaXe0bDhod
yleWOPCCoMmEFaiyXSzhZgZnIF0ssZ8mnwZ2j5xRBRuYtRRyxp0CGbjjsyXXUpSzKhxOk7zTV21N
NXqOWG6RIr9KxSFMHXLOstzckBhMtXWm8//2Ho9n9erWpGvxcS9S4jqs4/bjWmLA+dWYBcSjaS83
WGa6uZKTDv7DfnPFTGBywky0Jp7V11S+wirXEZgRdikhrKBNmno69v6mOUjOtqs82L75OeZSyOV6
4rvTs9xIakbU1omE3Wq65gYVixQTeyPU6qworgUCfCfy4iVz5k8QA/1MiBbuiIJZLsuBlJALo3uy
94474puXT/RC4jPoC/OJi7G2cnCUA1PeyBczNvmJJ/a0pgTVk0tqH5EzuSo92IPl3RpArIFnij5C
Ab78BxjWpmhTitwkVzj5hmAweEJf7gQoSa33dA+r7l1I5XQ5RmqLGCXvOuzc7gU4EF8S65Hc1hXq
FyHCB+j+ulJqZl7Bdhkkr4awFHx6ui8/RYTIZbjK1yBd8t3GeIEOm72uHdaUi6RZgdqDfavaIjQ1
Ud/q00HzJch3rfiUyeQ/nm+FtyCO0PfZ/83SQDRe44tZ0fuzqQ9kkmalOxUK16c8k2g67e6b0SWd
pUiD/BKT4cfQxMgWU0s8EaHCT0ugKnRm+nOoirM+KI+81gVg/6matcZW1GhKzFpCjtJwLDv+wShC
HSvanIh6fkq0YkhkF+8EO2NZYELl5dDcZbNMmS01zkmYr4SF7S4zC/UskqYfjsb0wPoAt1cipEMV
GBBG5c0lzIlkEwRkflsITUfOYHEUJRubicGdyYx76fYom84g7rQ0UBp45uJxKyjK07Mo8+APwMD/
+gtNzL0UQMqgf1Gc58MvE8xWuUzjUIAXcp+emkrmdLy6WExgomd3aMpGnZFYfXsgNeEzXUrfZZ0a
WDFFF0JD76zQAtvh1jymTTM4RJ40MrFKnTkaQNe9R/siMnyk4lZFTLpl+KVzbFUABsk/OIkcfH1m
yDsNcVuxRuUhntxoij9yoW4BiFLLmmmtOs14V/Vr5MDF0z0Mwz6YJ/yFFsFkvTfWO5dEe6JEt/5j
y/+SnFcWPTg4JBk6SGdLwY+oM/7tJYBGf8ZtL49Wy3Dmi1CSPcuU5393eVcdJTgJy6Ai51upu0I+
VVmq1YrYM3e9f/LaWMaB5WkuxUx5lbEOVWyCc968dOAVYmbTschm23gdpFFjS6LkRRe7o996O3tS
5UaJkLYbnvpzCEVzz7EJ38CtzGtVkVB/4J55sv+z6VEevPXS3AxsLUOpmYB+sa0OAm3tGBw9VP1v
k7w4imxB7aRk6ENy0PlR55HfjMvDzqBTmE5LNiRAJJw1Z7pXdg9aPsad28vPJe2mJQqudoga03hV
tW9NfY0XzlRzvgiXRcveEwvg/Wv5ALDeD3MSpsxoDarRLH91mpnEnAxTVjjmGv3dPrTTYQN1lHJz
NC9EnMyIqW6prmeSiUDBrEwDJuryA7bOyD9rowGir+BXLeNhYyIvdIhHKg5eSeE0cH4KaD1Dv3d3
nD3+QVpILATJfws2yqEJcXyeq4uEOnys8yj+EsiJDc413N6S3J1pajAlUfK4rRXnRpRu4l6bK2/I
zXWRKgm35Q2b1RQDN3UgFf8a1t3U6oLHGMlse/7tBTZrX4akp+kVqmXzTlzRFSMNBzdRoWNjuM0b
l55rg1PkIXf7TJZaaE8HXlpTMdtX3hCg/IjGZeq/qGs5wNVqUNNeXJwTnLe3qfbSMWb7ZCgOotFd
mOrjPGoePBkURMBGLosWZW0iwA8bYnIPau486uypiqUwrgctwNPyxge2YaxEOxzRhDbd+A8HnDgk
quu27mEdwmmTsaJPlHHyfFIS2N32N6Hm5b8OQtQPXkwnH/0KhS0hulfSP/qheuXK1bJ1XgsWzBUY
bGvaZOg91Q6QU1wIhJy7QB17cYaLEPt8ksf+DvD4O1g//zznC0R9GaFrvYriLHdFMatIXMY3FA4I
4vO/vT7hrMTFclMngONNjiIDIw6QgRrjCJZ0XpFnUN61fdkwB1rdMLQHWC7a7GXrIcsMXm9/FXrQ
afe2RzUU4RmxeTCr5xIkZDJNBVSDYE58dLXM0SuW6otbRQlMJaoF/A9ZboTBAWvMlIcajleJ66wZ
yrH0uNZqZd8uLWtW2hBL39IJ4oFEQWXywLHM0mqDXaVDwBM2PErMiTDPOWgbnF/n4RFPq2iASAlR
uNNvpIhzwB5bhk/SSiyEwN+k7o9cZmN0C4nNfPfIy942S8c+1zHyVJKZA0NteGOR1P+IrEy6+MGv
02K2jag15sq94VQME54FTvOnf6t9N9qT9DAi/q+Zkyj3m/6Erjoun8PEIM9GLHF7Myyd3V09/MB7
hvgvmuz+6JrARY0VjaPwm0xcViro84qtKTGtWd0MkwXW7TAT8KCzgYHifKqvZY9G0Eharye8owxi
ezBzGKD4p5k2yl1a2e2WRG9SLp/7VEx568IA3nsvQ4MLVF/98IN/hjvIUfBND7DYpKsGA10hSnMP
IryM8u0CwQNQjdCf1afjkEjw0MEMd0c6AaM+vzZ7Q3TSY9Lqu0PwBdkeC94WOrQyZgjTTFVEDpI+
eTGZOkXHLUjWOBV7NTK/qgYFxjbklIw+7UlySI7Jpf6OGdNjsIxjEGif+plf3gZ7VSTA6giu9u3b
QOxL21rz1nEb9MKolmcRzuIjOCJGmvi/m4+MpFqqnhwCG/t4xxjyIpwRa/osBnB86nySgEe8S8Es
ih1XtE5WE/OlNmj98GTVtl4W9x91BmQF2+qQMRUVLC4PE4/5pRExN5Vwto22Na4enEH9y7t9nHYy
Apee+mFWkexRCU7/h4VQyr4pLRXpDefiYrYJ4+e7mxTpKQ6p3gEZuRf6/2k1GcGDcGK2t1AQl4az
BSXlwm8VcNgCxcGpu+2G/er36CAO77/ttsWxDFaEoLIdmFsmIjXvobfaMYtq/CeUE4sO9hG5454g
nINL3kfJkuPkT8Fg4WvOccVteTYSLhvKTEXmesrOOHGk25BfhJkLS5leHsSxeekcgoMrCvFKl+jk
Crp+15+ibiMsWlKpAJZ+H/jVzKjuPrkrJG+qF5++5GUVRv0ZDSieNteV2kBr9JDW6lERsgGopjK6
v0B2mtDeKXU+JYAsQ5kvNWtmV2Baa2X7oB3VgSo8eCU+vlS4l7MKb6pySDppqXRBqL0gEZfMOa5a
mKD/Ar26NoVmGdzGpMC2O/ItGaAy32BcuJu5mrcdBKt1qXjf1JPsbTMZWEQXdHwLVCBwrU7/Of5f
0gqxQR4J1sFhByRfUQmwiBct1BKmSWCJXqXFMAWmyUJCC4WLewuLp4V5HsqTldltOfwOALSp0JST
C6yr+5zn8AjfxngwAbfgZv1VXc+AIgq6R/J0/5mlyFLtsALGJx63mRZh9pTkrQjkF84mvbbCYqDA
TcYH1PKpes9ts+LuL3edmvG9Pp3PvZdlaNgb+BkrktU5I7IG5CTXUDfcFmX7goHK07h4bDCvh9/H
KvrNUaNNcH0DSvPBTx4XXlaD2dbTzReMTcH4LW20jylmmDIvaOvlfrEO4bpaiFzaKus6TJzqfjgj
BAb0RFLmHaJmEE3/08BmnBZnpP8vDgdrz983hE9Da5ArhK+zlU/kmlWT4HNJMJ/fCn9ZfqvtdKQM
wEF+lPUjycz6VyDp3tGBEMUScm3B25q0oHscg+wh3ZYCmEKrmvZPjtuUc+p+/FQZpwt8zgJGIHB6
+okGoFzDZjwIWuhhStYsAwrEgG0Ox1jGDFrYV5B/2Taf+mEvF9x3iSBrhCb8Jwskzwv7vaiDXOCI
o2mf+erf5pkgWvsggU5Rm0iwyzFk32bLu2z4r7cugf/fWQzbMcbIUaFLilvKw/8tTZfgR2gezaAH
x79n3t+463vm16CS0CYYVJ6iNZ/+skoU3kraSLetrHahPuBiYUGwzeGoSUWhDKE4OxFb0X2LpOL+
F5K7PulzOjxXIIvO0LgQzm/mGJhWKAjG2iUKMxM3OJqaYl3U7bYaZPFlg2JYgnyaDnAf4Jv4MfvA
0y3s3mmQ+AB21VwApXjU6bDBe00DUlYC4jFVKdy2Z/r+l/enqQEsLDFW9vED4BIuEOYYjsuFy3KH
3nlIWg6VyNhVHf383pXA2Yt/ekIwhg2vKoPXCEInrFWPsnnBdvPUHEWC1LjajFCAWaBdjEJ4H1Yl
Z4Dfi+KB/yP/LIWi6asTZdORBpauc4o5iIoQzktByav2WchcW2wWY8Va2zMK0N3PXjVtt/QYI5d7
b4Vptb95twWVOr2whY0bk7x1EDPMKjb1Jm0g3WnwaQpcLOeQrVHFTLiGWrQVULS41yK/YAmajiIy
NXPAPw2p0lNUDoSN0ch6OZqUwm7MnlOlgYfb2TWJpvwJAZW9cwwQk2Ynmai0Th5urh4XyA7lGY7b
bkFyjIo0jMI+iulfRh1Wf6d82UKPfCg/T6qup2JCmInj5ZRyfaVVC/5Vleptb4LxIMVuY8uHeqpO
v4SKt9s0+L94v8ncWT8uAJcpzHv9hINuXfhIVamkmM3ZAs5L4kSWkdA10GhJ8qi1WCQwbfBu8iJu
hv1N/xlgsRfA4kvpi/tAhiWr++VxewkYKUa5ylJ+9RGWPwCExBgkg8lQfyM0GPt+0gwaruNAn7+x
ePo6OujSqUyzYvPrRbka2MC+yFDwN1sHLVkb1/lndv8evuKK1DPnLRKB0QWQh8t66S/XPN7g5BNA
n1f/wgR3frmyStLH9kUTq8Cg+VIvBSTSxAotvVRXyaGmL+RzLWbxamThg2swJ+CHIzdHFmjnnVBc
4hISQyTRunJ3Mj5z0MSTM7EgeHBzH6ANUdX3yR3K2hSgikFrg/s7n+E0L1/+MpE2kjficlo97anc
GqAErPGcsZQJd3XIIkM6Gpl/+XPLB02RYBBB6BWj2OsgzN6eHLU31KKVnE43uuAREpncn3BQo2V6
P5GoV9EBWJaSdspxLTPlHSxv8dqSA073fT9v88gvalytOhi21FzhWNMVLeRHGgUZbdYlBoOtAtiP
AGMxOfMCXfFCZKoH5yESRg31WR3fQBIHi84WyuQJTVJUhOUsXuJjSWn74UyHcXD2A0KtyeTrGoUA
mPmzWP0/vQ5ektZOEXHQWrr97e85oemqiYUv/JHn5fbW98dhpJchbjCyf3sNJoidIISbZurau6sX
nFeWh5H0rnsGZal/e4RcJy06dEGHbqez1V30HtbWV3awyEryCnWDjITrbd3bDdoSySV9ATQ0qJbh
P/0+Coem+Ad/Zqc/E4VIdjqul/n/vBv+3cgX7ekmyTzOIH9m8PdR8XZWX+QnOlGHU0qg4jcxnUOF
u6ABq3zezbtwU9gMYIuPaOPC3ljw1M0ir6HZAW3U/aArckw0zav8kSx5FQuyHnCIGkEMSR9wlOTi
4T9auBUcbJpFD9BjljGusACFWwpNIFI1lUga0pHbBz7sv2si/ammkBW6uR9qtMuMTBPshFTwNOiZ
bbMLeY+XecUyQ9cmI+jEI9FcbwJez3JC/bBh/sjrKw3ifQWb1TUbqz8YjBVobxWDxtplSJ8brfNU
FPVDQJcjKRj/PdHlPKjEFSNZbKn4pWAA6aQdTG1+TutoyKi9HzmvneEa6wECwvYXK22PkHEbkFPK
wzRedfDEf5e56us3UfDJS4oUY1ObM18GMEi+IR6SrZNNid8VNVNgcLapjLPAXK/9JbqhDY0+PA3N
QpGHxZb4cTVAVh7jlMnxtzLsdgB1h2YznWFgyEOpom8pEaZFpRACRHKkTfmSCFIDmulQ92cBDsfK
hl+1zwO4rNW2Xf8Ohi/3CfUExU8M+C4v/MmHftv0Okh2Sd5vpIZpY4XYlLFZjEuWTIqzvwPZFFsy
SD/fYhULk2zX9UZGbaS0Bi7VQ55YDrKbgTkRP1c+/jiCwcPP6AMC2CSnszHxhWG8pHZ7JnMF4W1z
mH9VgYmzEYI8W5B8Kw5tok4i50Fv1p2SKfh30HhEP+oWsNO9o3rdNeANQdoCs5Uhu6R2JzRU9qAC
F67CDFyaAeZy4JNXU2LTUKOEq0kd/pxZeBhIT6lGECN0Ph1n/dtg9StPxKuVbm/dGDDjRXJVODYr
ez4Sk+HydWvFk0CIeRVrzosJ+YXzdKP2GMYyj1LZmDHzzV3pLuQX3cqD5cUNofu3ABDaPcP42+PI
W8JsI/3/VHvukELtEQeOQgtV2R0P37UU8UE3KmPMe5v2VFd0+123QoPZzt7B9MWil+MyrAuu6q3q
LBEzpGoO0yHGB0fQF4HKI5bVU/pHF31I+EnBHYsXDgeh+JQWXuBLgRSdnpvb8WsRw9S0USZLwWGT
QLBC+B/tYJrJS1z8YGUBj85BSzAxcVA1xCwv9SpGxs0NpLo/L+BmP/IDDeEcL7kyfqOToUWHBZDP
kq4kS785c/p/mQ8Ve8X5Em5A1y+b14cXUzHtsUMkHSKhIDGR8ZhZf+naW5Gw9ymGXSxFhhEtYVt+
LySm+lZVTYRkdiixen9w4e/dlpV+yjXLBZu99g8WM6wqubXwmpfFzBRPj+iilxtY9DGSylonFFZF
QYMwIbLaisuAVFjLzpPoqytLV372sJ5yb/04mDlL5IW0wFYgFVo/9DP6Sy/gLsg/a5dryKK8ERIu
kdLDMcKIvyqF5dwX0A6o9rHbjt4zFOpIM+p0VLt6ziGC1NZKYQwHm7GaZxQvGwBM/XdTMh6R+vbD
hOwts2/jMooMVPTq748wMwdnnSGjMf0qzWbSHUeIMrs5tgMgerNZtcxSxLRPeeLzSrIxjr+0Zcs1
0b6kPUOJRD213QB/F4TnSjvQSW4haITGQqhVPm+vl/W28PHgzbvdps1bG2r/VI2mef3IGI+d6kbU
w9to1Serw3wbZc2ZaxdZmvmuz9sdndoOm8vmCSvhXIty2v3FTdvahfHhD2UoHTtXyly2ftTCWJWz
xx16VsZ7T6RoIvweTHrk1y62gP60i6q44BstGT+33DdvPxk7VlKh2CNKIml938W1TweleHMM7Pe0
CJdWXUKSFuGWrZugkuPM3sBv1bf2LmdIpQUy05CpTDR9/iIf8z0VBlItA8Do4QsbqyYPfNS9cnHt
J04ej54pXNavkLMyXXWi5+1L+NjODJEPjkoy4pnArd+T8JjR8ApRXBBMjmL8qujYfWysDrINV+iE
yxrKkCDyNboLNLL16rJowFmY/fsel2ZMNo8+Jhr8gVLYsNLsOASyb07I5HNqSQAoHGaACrwA9muM
bWAnICc0VZVuGOF0kUZXNbyplHOakXOQ2hxj4EhKVjU168jSIghryZQnAHFtgxB14WdQjObalOME
wazXOk0uABwSrBPoJyVcuVs8OKcyRreA+QTz3SEfWucbr9QK2Uoqp+/f1a5t2mY/7FS8nhpOVJFW
zX8CTCqTUrIgvoplpXJyO3bg496pnBDUR/CqhvOXfnGTyDdTyB0DvZJVBBkj4vv/OTRh/Ep5AsyR
dsJafZHVdSZUkgy0QVioxEabknC4pySSglUuBKoiKGsxrIPVU4uF0+uUO8+AeJuFVPiWYACHPXIn
3cSnHfThCeWdIj5Z22uJkcWmVMjTVDSw8jliesaul9+bfr82sWWeGaI4k8vrf42YeLDmASZwk7sc
yojFcn4s2KAMzWuHIww4TrvQOkiPgH63gzvM+oh2df/gaTtP1fixV4m4xH6whgaKQpgeI7FY0jjS
IWHJbRxOQOIt6C3AhPbSAPvZzZmAwr7IAvTqfLu9wwHqq0uc5ncZJEbiIICJoaXABJzS2yIhWwbc
mqfV6tS5jLbemzk+QCuL0hb+be8rLsXBB+YmkLyUSWIRqLrfj9Po7WsQbViSqV/VYLJagsc12LSc
DdiVNxzM31uFQPdNsmXTmFpeQ/OeMFBPtS0qJ3AxR/RYq+7BGuPX7YRLX11tbaRjXlpl0sfGk9Q3
jyDjGjysv5Ff1hpCTjWJA5Dsy6mwBH6b0EzwAsQ2oGyhhGZRdfe1KesVqx2KXEFGEPeDepBgin4B
TiDcdOgiAE+suGHAlJ8Gdz3lvwLdiSpv3LR82mTya5ASVmulNThXZwyxf8D8QMWWcJDMY6WalTx3
rYOLvBbGR5yBTWKvhi8iz3AL+Pof9JQ+xxt1OwyQ3OeJi1qLP/THLakjs6AYYXKY+wFMzunueRxo
T5oG5JAOqV2V1bR9dwV5d5dP+MDd7ill8+mQszDyTg2TD+UXxk57B4wyOSKntI+KcfTZF2/UMcEU
ZWcE+naJVqwdl7pUZll3q4ZsaM/n3/PfHaGYPJE97bPosq3K5YTKuhNeY8MghpYw0jEX2lXoH3Km
luhiVr27zRdUtlC5/YnCz0fqGlrsXXVY0UqhRzfLnjvM+3fJZFO7oNZcjurmODDkoutx4ADfKjqO
X0KYDsqqT2QLa/DXGoRXuB3X3F8mQ2mp8Hu1skLGN8083Gs6bdTZA+4+TVNTGF+0XlIap0ljrKys
MrpoRnqY2YNU0yPO0wm+jvP+mBp5rimBcccPrXSdFEngSOM4LJmPFkBqnaWBi4ooQd6vakiuWH6L
VoR7wRQ+at4e+k6Wuly2rfECpkzv+adku6NOMG4VMCKDmGHGoUzaDv2ue6t+7hefwF4LZRNPL+BM
ZMWQXQOJKzcnnZOcjkTOtFUdjWgg4WBcuWnCCmxtkOENVHKyzs8bH4hlln71uXdxqDVS57IWycXg
gDGbhkuVro2Cc0OXB2amtkck/MZvMRsDdXFaRcNtjsoPY/lSYkx60smJxqkZMRtTDQmFfipa2Aa4
vQFUGr8po1auz9dznUIw1TBdMWt1phoc9H5GyHnB4H46eSFihCdlrXMo3f9QXOumxSy6C5ffsROA
RigLvMSuikFWIgyq+zv7vs/SRYNvYlRnWqlDauVM4pnUi6fzrsVjN7Aade9lQxcQZLsMeoIk2F4f
62cJrWnTwWiH4a6gMyQIjZj5Jt2GgBv/xJK7tb94gRpmemSyDsb122VRgc7jI2ysWha/8zNFWLgh
4jXMYNFX4qn5u2XEvSeCK4f9Gq7bDq7X2W2mVpO6lbU8geBkUjxWqPwkzTnfmKsFa0SCbDFVcf6D
BRkKscPAZVQ7i1JPmrcFH5RfSv7RaXAM7r+XUpLi1t02d9h1sh7lLLVef9GnziUf7bHNXxOY2n54
Y5HyhHlHYp+fHMHU27ObSo9OcVKneNLYaagANhRYz53akYLnceLdKBLD5jwoUE2OeDGp4x4h8n4h
jZeKCocsI8X1qTlJbBHziKqgMINHUZzSlL5XAyyNOfJJ91XEIUqwuBlSQm+/ENfkGTNo7Eg7s0cL
TiuERUoKS+uVVcyx2N1G8jmcrV2lseug2sLNKgdsOKWGDYTSJkgiLzxdx3K6lZSDMzIBo8owGplq
5jBD+YGIp45zqsqW9EBaHO5VmIduUZgPZm0epdVjar/4PoSu3rDiSdqH4iLzLp6pJY8aG+VKjuhg
6NOEaR7Hoi43Bfr5+q0AxN7JxjqRyY7Kq357sjhuB+sz6YoRnVdcvAyW1+oHOuAIJT3CLxM66yIH
CPJ2sfoYGrJhTWiRSc/uGkLjCdR05WJ78BEEr491APiIX347MNulECzHTun3zuqZqh7IsxquH4Yj
Epexr2VaSY3hFabzKaqT+BvHC8HhT/hUm5HpN9+UAOBmVWtu6XPMFIfSUs/WRx31T5NyTwuJ4VbM
D3bwGsFEn94vyo31VKuGOG4mpnIkLBLQ4Qcs8vZ7jwslLm4ZWG/IIlXTtnl/7vJeT45vONhDzX3A
mXiArzW1jhKhKTE4YRoU4BHF1RAWhyqnbMMEtPwvuamCZpt5FajO1gdvek9TEkBHlGxGrgojQC6W
8GBWcuTl3yBMFySkaUx3GJEcwpvOtDF7jrC+JzTPh/hbI/eYWn+aqsBAP5ANHz68p7Ccw3wzZelU
DWubfDtio/WsTOyyvt1VlbO2ZbOAB0WGq1rCU4wx4/iIoI59ID+JEYUU6kiX9QnBS9kyLrCSbIH7
3nDnB0GL5bwVnHQDOvXIDrpJc7J6f48drT7BMRZezybh9Ta+/s8YYCrXI6Nq5u/+/pm8rMOZzman
gZeDFjif3Hq0WPm8/+eQ3OduL3Vpd3Am3f2lwsg59695QUngM1I7XXjipgNCXcPaDpnPSVsXJzkW
e6AqfQEeT+es3aeFQnz4ZoE6KilOHLOVO4WJSi9sbHFg1ZXUdcbrLbqZS5ncj/ndwmwaDOaB4/8T
8swQiK6FmGA4iaPDCLbf8KX7EgWuoQZmFmZm8H3AGse+AZv+fNJ6tVterl+4a6WPlh6khkb0cFhN
WRbyjetSJd15jsZJhxqFhQPBq1jJ260XoYCWFl6Gt8UxW5XKdq/D7XCE8csXMZAUpIuhnwigRi8I
jJvXe6pxlYQ8VHvByVj2pzH5r9w9Mwn5yOTHQkeBPUZJM595GltXnepIr+TYHfTum3rNOqhyrNck
NvBMjvgTHJ4ixdjz+T4lGEi3ST10YuCF4PS7E/9Mc7iafDFslJW6ASaZk25b3XqlejYHipRVfnkw
oTjBt/jOkduiHv3hncAfYY6TsLiPB1xyv+/+IvRuboy8WFwZ6XoQcCQkABecbg7bxApKXES9V9hz
12HY8lNN7kMjOe7quK0pEgVH7F4naaOeOF6iUm82YqqaQiNcFF+PmA7dK8ckKUlQMrc47i4O4g9k
U3E0Ip8HWU63OTbKGgR0zZyfB0NPyWHtLAnkscaUhQIp1vq69jriPOx43xSXxTDGIXzuTyXLDWvA
oTl7+W+VbOgULVcIVdoRjnLAJASLiSImBu3iuTheq+s+pY+Zr2g0TTz4EcoweZ8bHdkjNrCN+6Re
hTeHyphR+8bgk4Mk6ahnkcxP2Za8AzhXLsWA2oFQrcAzN1pBONIGcEdljvfzyWpTG9spgq+ogzN3
bwY0snZywDWCXvW8vmt6uA6+WI8LnMrOf+hjRCB3A9s/+gCxLk7ffazi6fE6qp5q7yjqb9kBf0MR
p7NeHu2fvmkuKym2OLE3e+CldUalhdf1RsUG16ca2UcmGamKGmRjs6z+3qds2E1drm7sFRw+pDN7
+5DQmZx6bFwQClC4WRJfXibDo+p3v4wmelvO6EZBQsIKIU5xKmGpxjCFZgy3swQT4ihCPtQNTUFL
iQPj9V/FPm8u4Oc+WUw0QOrv9p0dXRgHl8zZcnca1RgO7SQdO3P224RxK2fS5zTKB9uavY1OsvPm
lyhGhkF8IhXwISoA8GJARG74yzNQZo4j7pmqhDlZcL6vKCp9xSzQhEcirkl/cFEktM76Rxf5XXO9
p8m9lGTSHaP6tPZoGSnzxs4Hy8BjnKXTPlm/ws/PSCF+Yn3p6HkP0Qh4Jb0hM90yQdeJeuXhH7XF
jQ2FMXpkU7raAzWRJX6CE7GP/z9TfvoXVs0SUUNwuB8QtT7aK25f8iJS6k5zBvsZp5wmysWRBGFv
Sr4WLXh0f1e0A0l0RBqtyrRopruA9GQhhW62RYxH8z+7oJ7xs6jSfbxsDIV07/YBzvCXF/EsWPIW
m4+Ya4UA0uRBp72tn6gQoLnZxzvpTksEuAF2Las+p4OgnqIaXgtaeGVEJI9E/YnlS1xVxO3phh+n
01hGM+hulMpq39aFr8iYqQ2mglqw1SB3BGGVe4LvpoQMnNraNL7a0o8y8WVWnbp8C1OyrFqJPYYE
AQlcBojs+z95rpD6ZDfl5H0vywACQ0y7176ZWHlhIqOR3sbl0k0yP4576eIU9Fkp8h57ueDjU78Q
J+7xbP3sVxwVqHmv9TiwGJQLEVsaKhbAYJ5whPAqJmSsvyAXmFvZobWh93q+tmAWwoOMi9IZ8Jm2
EQmnikApTuEl8ziE6r/nyLZ6pEQe7sfqrMnBJHgML01iIoY42KGm6JjJHO7GZariae8Ba4A5CnAd
ygYPWVelhDUs2/0trE1TF5m18p9VQyKyRSkjmGRs3rRVnr085cKuL/xSJjdJl4oP80bDin9/NN6M
NoI6KeFWfCbrAo+Gw/XfvIsttbbRJKcGkR3bptFlJcbecMcDO6wLS4SOHD2R48uk7b5SSye/1Jrs
hqNpQUGQ4Kz8MsF4r8fH8fUwyhRqDQymDnsvZ2IuYq7uB189dgxO6hVtwLjjv1HDWQARQBojvsYw
LW6C/c1mjPWqKIxbNpr0/C+2fGYM6mZV1FAh9SSoPx9rp7qzQnnztWUQ8d5NZapqK8enZhPJLIZW
EDaUakgmeeqn9aNcrkoonM8595P9ZeaNnV78BZKctedBiuFESjoPGVhqcTfRRY+SL2FMXj5OSHRA
Z/m29ruI+5Fvgo4UJnyjh5Q4uYnx1NJ/GYV+LfeEVU7XdkuNpobh/G+cUMgFybV5I+dB/St68bCO
IxGyhYQXChbgOtEgDQfkGkqhgB3jRuj46styapWiLSzpJFXGq8Lj4X+rYhtEzpF93iFKTMUuHY0t
WsLnf8rMLG8EZ9QwnN4ZNA7v81x5heSXwQKY1YyWzkyCQ5PfVM/z6X5QKDU7huF2vxGNiBGoGm/R
jZOHx9ppJDKxYYpIr1zTmL9OQk+b13SkBaILrCTYgVFibVvVm7yjfhR3a3GBpatDdPXYRT8xbAHR
FN8IIE05k/0vlEZqq6NY3JuFSkSPF6zU5NQJ5GtR5VUdvukGtl+LiyIWBHW3yRDYfWoxGsW75CFS
5ucRRClaaNuAPziOrreDaRWG/RKFTiugqvAE3ZtQaKBdWofeQFjoTiSGE0CKTNpEmXLuJPLPxwiT
j74UFa5i58PV6Gf5SCoOOs0c4KD1s9NdfEtbL0U3NQNVnbuZVzpkY1dzJksaTPiZ3C3XFSIouyAt
QJH5IkIfXEFOQBmSuo/ZBuULyvxJn6jqd2gKSjjqj+kjKn3YdUapGBor2SdNEY5u2sU9KZyP1ivu
KeRnm2IM2A+dr7UAJHc/ei7e+TnZs6COZCqq9N7lxo0G72fh5Vz9nXQaftzfayZZ8fCh8OACsr+c
qZ/7NYSjEZzcd7WcUesF+X2CE/upDV47Gl1FWG33SkUWffPD/VSCaezo9XtvkjiVMO43gmubZi1/
uS6F6+PxLPu0+aIlcPcbY39lDVoV2WHZKYtRGtl2oMhYZgCbHpkJ7MdJtlhmXl/PShvCBsATKqdK
K5gMWBDgxzfAoBmp4EN1Shozl3du+rIdDg6EKapfWiIZdjnRv7C/t3i8gxuMa9h0i0S1Q8HcW5Y6
3LIJ7leDdrrylFkZPv1ZVXoJxXdd2m/+aLU7IRjQ6pmi0saFLubtt1xhDFEoEp0w/Tk/UqUFNEaH
ha1wuUOwHmrK2yEY2XmnNqnF7KJbwmdliWaVGMmZ5ddzW53tXcW0T2u+SOtRUjH+kNO+9u8az1eF
A0QAtGV6N3U/6NwUFQyUWJ3xnyIxov0YCPwGh90bcJHem3X/ycO3bVCx7dGFJDKR0VRy2w+59/Zg
Fny32uj6FMuFaIOF3s4BlRR8K69PQXfTxRWg+/68gJ9mak1tIQA6EnDGV4dTZN5k6oOPfLju/lfK
FYeUc3K5dKp8dQG6l29ytyz0+t3sWhy/nKTQbyz/1WmWTbtQUVtgU5M91OhHK/gX9MBiSl/dsHQR
Zgsk+omErsAyu3y0U5a4wrJ2DN2+ZGcnVpd+R3ekKVnzUGWWdjEsyr1ATiJNvLmGfY7N//bWSE46
E/4Ke5FyAsv/4g0U80xJVTmJYx8DbjwYNN33oycCXIHcy5pQ0747boQjiXHkGSMLpwNPsCp+961m
MaK5R6IS3dKXxyOLWRApMIHneUlUOLEIL5OWg/L33+XCv/lQlfbZIQaotdWbntOwMke4Eft4PnN1
xKqA7C4+ox4/45lWShAvHk7CI/grp4Qsek3s3PQLjR+JBWVfAToSh3KMoaezspEo646LyGqh9SBQ
/JZZmX4w2DeEztZCtTz7wguRlX6LeWAl9wG1bs4zksEGItbX20sa5ekHkyqapVr/tfCgcn/nai5N
X+U162E8fH9eFdQtK5sHePSzmaZZI2AqOX6pdXaFb6gfzKzRBjrJubJpI2mQ36qcbt7mJ4NO80m8
bU2JQNTRzV2GGyOQQXVl2mLhfhTTibb8ogatrdRYwpoUawPifjByzocmn9yG6Y3YCmpZZh/OpfEX
l6Jy0KiElGC63mZIcW2CggT3x3cSDByVVnu6ce5lgMHC1P4vqsd1SZHEOFsonK9Kcx3duCOqzDBf
aJL44vpiEV8iy9jADThLfw/+d2oimzPU6XoHVwVODpswkQZZXYnlcJsOIJzLnhK8q7f8kTaKfqt3
6VA++efofUj5LVRrkvslXwylcE4NRhhBl2wafJW0Y7yskgER/zeIAWxfeZwPr/1MKWAYa7ctUqq1
kd3V/vnqNYo0FtdWZv5OV7wwNJrTbwOAkNgvhtzlnJxoOezqcqxfGfHTdKib622V30BMwtXzOCNf
jOsYkK70Sht5lXGNvxqYV/JGCcvHLQTjoAoVaP2MG/EvMbMhblgAI2DSKXjY21IWPLp52k2oKS6l
x5AW/sFHl2mGQLiPVk2XAuVur62JVE1a3Sd2V90xLbuXrlMoK7QNp6kUVHmXEuzdZkj6BnXCX03A
S5Vak0iLwgcK/iUKVpH91vUWgGQ7McQMUVRXOlIQ8fYrrZLpfBgVo4ctdLOR++uf2CcCGhP7aqE7
bvae3/LtcpP5ha11LC2sjoufrXdZo2+Qp3uxq1ORwMmBDFkkP+AR/br/zLwt/covEBjz34Cy3j+y
VOayKKhoWcL7BluyNAQjoGd8aWNjye0gsEcv3JWYlNMPj+njnw2MS4KQm/YXwz+FsZZ/p20gursh
V4Zz6FLwZ5ZS2+puaZdkroKSPc1utXdAGOzbimcY+HDS3lPb5ejM4MJDw0q9X7FIjFHbtYqn1S1x
7BW9FyyIk5XDVW36DwwjvmtS23YYX4OURrxQMe7Lcxfy/+cohuM1pQYVluMXEQCSNsJbvH8nafC0
9QQ5WObcwv8T4cxfKkOIQ2LVhBm4lg0T+pwT4EgPJQxzvu244P7ky+JudMyR2LQRbaE+EL9zJ1mx
ctrwjHLClF7f8E7jhqzqUFmS5KvCj6WvmKWy/LP6IRB5bTNiEZc0HJQq7RMDhJ5rBLTzVUFl19N6
wieVlIhCkgGjaxr15/rI4kbzniVnKIjy7okQ4QJ+ElMj8dTALgi3eADs7+jZ2dWWSmOIzbbqQ2JG
dzdoziCunTtiDhsYH8+knma/uAbTm32jFcLcOG5QDxuxyMrlUPyEi8GhdZkgs7MjkgGib9NRLeao
myyw9Zml889C/UvpBxCbXRAMBBY04nc6ul/nZjQTcLcVhCUjjpCQF1GIxdd3uL+9C64Ij2s3/bKo
cnpUiqjccAuhSXqa/olvC58Bxd5PbVXBKhpdjMJdpunp7APewh7LkKToLE01u9ORMErhlljT1La9
cCV+JnYVAHgfaa/JX0wWBZkXB88NqJQJb4NtuY7+Mc9fQpK4zB+dxShGC/zq7V7EseIVKJ/cBNZ+
0/+1mks0G9BNJmEhnviEJTHQ+XaIs92hHF8gzgEC7W5EUhuOZFvbzpR3ZC7/MyOKayW9OthimeVW
SOvrbyJsjpHGWasHLGSOoKIqPYh9jWtgkhea/If3l2lrzy9VIsBqKytALRS4apxB0drPAcHdzcmE
js4eoX1h5567V2hK6HWV+oLAsjlRxcISIGD/A2FA8KbX0flF9r5jkOJlLQo6pZT2PjL7RV3tMsM6
OKZWx+7jvoB7++4Fnk+ChgXn+XK6f0WenGICuwCXNt1SNlUN8ZReAhDc5QR2Nh8SbLjl5GJZHrtw
hTWxPtbONtktwVn5etRPXrE4HFaOy86kRYL/oW78PlOIL7bAxJzjYfBynEigWpf+txtB+kjF5dPO
hhC0sZDSmSutUUYsXiIUMBTB3NvxI05+ViZWrywcf218UkC0aMQyo4U2zOj2Na7okqJYngp+pGQZ
In0Xi9ERK/VSdzDBo0BjCtoGK47LS0CIm1GFWKVhwPqVVbXWE6QKFXrKOf12EUdnjj4chVBZsPWK
7EXmrrJ0ghATH0WeAWKjIDK5IsSB6yDKKfaO1NdAuzOTJ3B+h3lPLB9/t3agT75izADvDP4TgFe4
mV2hy3hPrsmfpdofjOJzkectzoFBorIA8uH5lzm9RNrdZr0gwMq/UGlcHpmnYvk7cE1h5p7JVL7d
2VmDytaOSeCCtwr0XmSpvfU+by3v4NKJjZew8V3H3SP8OTy9SBMT1wxLiycfmUT5eDh6HYjwzCIa
7KyMqWUhkymp03N2w4U1BOs+NK3EaTdXpAn6FcZVpDU3Qg9Njf+S/C1RcPp3i9rPafl1qYFX2PpA
T86Pn0Ic7wbN/tGfyIK5roJ/DuYbfp17RnpbMZzY3oWFNjQnsExMdNetl5uvQ8is9Lmf1UNrqXzZ
5juxsBo+q3fcAxCrQYpUapSoxsIhwkI0e90yK6ZApZCfuul2rnjkf1no5ze+KYYDTWdNcBYzZSV+
4PjGsfkLRqnbHHyMZ4jlS63DsPz4BN5VtTzYLHgMxTEqOGc/Nd4yrivXh1lAosf/GGtLSL4lBT3r
Wfsv2XPw8iLnKCnXjen7poCM9HfpyaXhUaLR+ysA5DVB+zC929T0HO8+eVECXVJ9wuSQKvSkLo9e
1zakxxWu2JWWFu1c+SBh5a+eO/9SL2IHrpdlxt8FW2WebAUUGxmX4qqC2nkArewDpUmouIkVJ6rJ
YXKNeN3jMonAQ/RTVQspD3u8WwSlzBZHCXN+De569MQERGz5Dy3DH95Qt01nZKm8oJhNRfudCeJS
YgTmNxoOtF/zJnQpU3CYgRml1xcd0XYMZBBlzsH2UvMBFUcR+P8kCioAO9fvJUvvWghqoNR6UXaW
AdKdoTOMylzx9lp0OsY4DwJ0r+78PGKnNP6LZMPHBHgVB5N1+vY9griNVHLnOBxcEI1Or4+pVYFF
TQysbqdWBAXI4UqT8yZpxnRE375McNdGMdeF169SgBxm1mlB9IPe2NSX7iy8VQqARfzOxlegoaf/
PiRxYWgnx+NHL/RIFWDRkEuakCftWxFFL9PiHoGdPwhuRlTkX2c3/GnSDldSbflnuGc4wJFuE8Q1
J0J7N3ffn1iPKEYKKHHJC9wmXk1HHUFGcyXr7LmYItaSzZdfz7SguCqUQ6juZ5pc1b/RnBXRZWw5
VhamX43s7IHp0P+tf5wWXSCRmVl/uMt111yR/7yEl+hAJNTNtdudS8TCdRuH+3k4Tx7KjgQ8sHU9
uXdW8GQZ2ETdYihAs0W077lLr3uvEXDSQv0ugPAfzJWLjjFLCee5m/WsQoswmYmos2ZDsSuKbb1E
TY3ZZPKbr8WsJ7X99xE/QnMo2xjDHtD6Ip6Hvd0Imr8y7SspqVh9XNY8nwdZVlTNoPDIeaaS4FdU
TFeU6fiTpbEL9SwovDzUajtVZVBv8PrLG/AmquBUwoNni3XHe7fPW9ogmbw3WY+lyfQt3XgCnPEI
u0cGd1lxKiaxQoaTc13Gh3rMKEBrX2x83ZvebKD1jPyvJ0NnIgmAR8r6WWdaAPYWl6DWAQVXhNZM
2xt3gyssrGOMfS18EtuX/XHSdGmFrEOMmFthLosOVzr3aMEqsgm7ZO+yJWZf3W0TUsBma3BJLygM
v2cuc+HzY5VbBsVIoGTTkPthNxb9qgAidlsG8jiB98n7QLbee6qSqRHjUpdG1NmYQfMa+lfpwZGB
TBcpaTK2iHZXd9xJuhFyMM4yhozwnxX6A0exshW/97B02X5ITmRMH0ptKNTK0y7Tm/YVIpPGW8r1
NMSyIVtxOzKp/9P6zi+rbaLwFXPSJoina2PUElTV14kUPfyUSYvF+5eGECwA/JuIn0nsvIVbtTpu
v6ECQlbD6Q7OJaFvZRCL9yHziG9vsQC3je1/Y12468L1XEQx+540Wg/X7VkXcfGXPxI+rKG2oPn2
EWE2oWGwfW449HH2crwr3X1uE6ZB5DUN+895P9oxQc5MSJGBM7QjxIHMM3divGDd2wab3vKjosGQ
pVb0gvIdP2vf2LrC3+0d75CVAqIGLHkvXDbzlshWbVLLSyfPZB+ptNzmnHJqCv4YYBFeiq+BfoFI
BZXV6y5YA3UqHTahSKZ2Tbls+FU3p09+n2wUpmmpLf8dk6g33bM2st+Ce4vg9p1guXCXZqy7fpWt
eWcCyFxkBeLDl773P0LKyTOxv8HpSQfpU8gDY+mUrnuMHbMy87Kw07hZlRgv3YrXZExk87r4ffrn
/4wUMUMf+NfurCxbHDSkkO2uJM4SULUR14U0DKwJIvSpmueTxmKVEDOolJRGnEdqsDGQkanKEtwa
sgRX3aDcnFyIaI0r8f0itbxNqfrl2/zTVwnC1tW1ZDkktDUeeWKvwpuZzgenSzKKCV1NlctqMRTL
cuA5xUUMp7HgaNKAXXrt9HBAVaeTwP2ZJkfqZSLHSd9J8wYKWeJbANCc4SBPaxrOMVx21LeLLTb1
iZmXKy4BPDVGwSMohVVirBUFcOihKZTUkGXMmQltteBzV88E4jjm4eAhzzX3oNPtf9fmqthFfZLI
YaHVjBclq3PYxedrO84rKf6MSdy9W4NiLPico59VggtnOYw6fvMxEQKW4Jms1Q5SRUijU90VfV5u
xQ9WiFZZDL19r/N9KROmIbAIc+hsGG9521+nXmLoAcWn3OH7kjYPxzJdb0BH8/wZ6SXkLopc+dLi
FlkGaSV36Phs+hnlheYgMOXcrpPkfcGbHFT+UTMcaTBXd0XMJgT6ytfQns2IRUMjPDPAwBxLNq/N
L+CehvBriLfDCB843TovHM5HGMCmHE9tGIaig/FHVumWuXkYQzGXX/rbYBf1tDonVc0wVOkWU2Q/
CkS3JleWflHG9CFjKTosnqh0SgTZnuQqwHUJAjGmPJuA8ONW9m5mlahy7BpueQOdYnj+AjJ1KSER
9th7v9bN5jlgndp3jSuGmnMPizIfiMIqauHhRtrxTqQteTfMqaMsQIqAwzCy5NPGpOSyFX97qn7q
eZgQwlwihjztVizUjUG+dUe1VsZ+xBtQ0YY3O/aprmIlkGcnqXDZA6cRA9jJu3/8JQBRZeEd7dmu
O1X0iB3vrs1aCQfghaQL0hDR+oe2w3WSeD/8QdMnXw0vZvqJeFUYAZoacUoFZuRO2uPnBLFCWrfC
3Vr5kbasQXvDZRz1lNOBEs3lvfEffqfLJMwb9HGsSoQ9qNmA9D+pupZgc4e5S2HfR70qntWXo32M
etXjuOQQnGWqagNO27RCnW/ZguqR4hogITPGVgTJvDPEMVLhTnAE+SpErhOhF1gXmjP573CJX544
Myw+QK7fF+vT65+ofDSoxTbkFR1q0JmXCMTTA1/rgk5+QoQt9vYRJtzri72mhWfdnc9v/P8hSTN3
DtZEEHTyHoebjfIPacYUixJIcg995kiPmYpthpLgzqZqrtFIGdYtFa5nfySdh1T5eAQ4UqFvBT+2
Uj5JvE/0caTFFaPgIdemTVhdkKSGUWU3Fk+WISdyLT0zI6fdOSAuCyLhr4Y0PNMZeOA/cJOiDD/P
Rt5yMft0IL5RAYSQz+gnm1N+HdxaCK/UpjbuUiy+Rccs2orAzOvsnztmqP7K0SSKgXb6NUGTekty
eITuRE/wZV5OAGhoPOHBAJXK/0lbsV00EwxwKy1TslKlYgpeFzSjWkhHu/uzNzRv0p/Csw0VV/pu
Z2A5zIg69cgp3YZb1KEPkoFee7oOca7J/uEgVv6HM/YiFAQXFnQ8XRQPpIMU2hBZC0yCLGs/HRBG
PuQZgzEcJwnvvjBzsMh28Ejm1ZouagimGuQw8ZdhxAdGBEqel6A03isn656hNlR9ZNjcVERr/mh0
8ws/YreHPrf52PCmb9p+J6UXnFsT8qddNK0QtQpnwkpFO3SRzAOhk3L/Q5WP0y/Ed9t1KPeploNU
/aGTlNk3eqyjho5Ibp/U4g7VKT2ZKx6zogQM68MdpSmUkYvdiKDE0gBYmLmT+rG03XwtbAKjPL5v
+zHj+mOdo8sWxB/wc6sHQFDD6WgZzwuqxvGF0Os/uYz7XP5uBMkJ7ya3w7uleOi6bev1fL/Ttehy
hfbA+3uinNEX1BMcvAzI+LJiSFXv6dDxvLZ/wqeuBI9azTsvmRky+f58UiHqmAZgQgkeGp9i7Inh
VEZ9pfrXbw9WRSJZRlX3BqJ/rn9g7SEz0yn4D/KZHhBvYxYfUIJVbmava3xoyxw1SOr8kZ//B7SP
7LQm6Cm2iKG1TyIp+EI3NOntZEbwYXLFbwyIdP/rYJDwV4XVVJV9t8bzhzw6kdxS1ThvZrBO8ok7
tCB9OXEu+lPZZF57I3htgmSZ09wiF5t8+ANZHmMgKo7c3Jl+xPgdMaWZuhUTl7r8qUwV/v8qIJ5G
usdtAcrZ3UyeXScphkcPQlAqemD1g9O3vGHtWm0KojvlGMzTmSJegYMCnCfD+9y0E2MSDrhluOgj
q2v1MpNh9pp7csX0xw3DePygALTJ3lXyAT0/eaYJiGg+wm3V+axScPdyEIHuK8ALaIhPKSTMIM+P
Sk4Y8erx0k0pKLXLaKW15pYUfaKpGwCHgTB9t5E4nMge4pCEJIYTuZa58lxd54QmNxoxyfgCPCWu
RMPFaYraiet2pzziIodKpOfFLuWjMkJzFtf4JlaUTTwh0CTBIP1xm0GVZ5jEXJ9ivQiMVaBelnRa
KPBx7l4Cwnob+LI2vmr6qzpBMmmLrkZbNE+zt34RPhIrvKTZCClDDrR7MYkTLd+2pgxRqQifnUQF
+EGu1SJcWAod4wIAucv/D7+/+FZXncH3VmtJva6RDQoxb4jdI/n7NOPl8/fpR94Yt5lRXpn0MkFB
4EK4IHrpD3yK70nyIQ9kfDLFnd/OA1VwQEIo+y/OBTpADJ/S4hJiyOGJ4pYAf6wzQQahR/le/eRh
yahb96+Zez69d4wKEcIQmXvVFQAhyuu6CWxSEw+hslGwzeZGI+VJq7uj23j0fyOk84BojxjINB0H
9Lrhn+Z3+gwAQdrS1ISGJiBK6AtGtQMXxt4cj+UJv04d09r2swYqnWteZyoxj+xxx/htSKGET2uD
zdFOwEVbKvmdTMZbnb4bKCZ6GoRWSmlIUmlY09vwLUq96zwh8s789Rg36UpLCDYVqYNffM9cj0Oi
TOVySILtYgrd3CYSQk/HN2TsBgxYWn1Rgu+e0ASrO+OduQAb3sQcqsDlr2kUQjNPDybf3iS859AA
miF5PxKb9Gh4BwmKSsg5ogvewWPhUHoOK4vLs+lHMiZm+Hz67bQiuAuJ7pcDHaBkxeWeWtDruPRV
8V4UC3fkVIHcKw0FeNTLAV6SBctYpawvsxgJPYxSFSYgafA7V5GNJjDS8JJVZZ5TcQgx+aay42aW
lkFLEEe/qIqS+eVBWMv3vBmm/dMDj0pcZsmQPqfYxEQeJBFq1o96pnEz1/DpM4KUV39DeKQQEYss
n6DJ0BtDY9kNCJWW4yI+iW3tMKz+ZuRD+2UQ8CVJJJgVYulaWYCC7wNnvcLRpcnFrYTJWQxAJ9gh
Xi0KvGEubn5RULtOAgtTxZkuwhU6JKaD7AIROBZfFEuHRHb0Q+i6WzB9qtxOeW9ZX9ZlQrj9QF9e
x9kmmuNAF27TXL0KQgIe0AVpRRSpPLlqgytXEsAkWkfifwYBh5KEbcAFoVm7jCRsBbYRzNqhpmSo
PwgWVq7mYgzePLehkNlR4W8n1pRQxQjAdjKmgqwRLEsu6a0ScLjzx5yXugt2T2r6+myNoa4oJaCk
9La6P+mOXpKFS+wsaVCpkTH0z0OI+bowGiW7J/LQOmSxnK/AeyP6eTcL3PJNtoax+NCgx1gyHIOG
vo3ej2R0+igRw5L0qCMEdnBuJK5McRAj2GHOUlzilyVaUL/GcBx3PP/xAaH/J4EwofcLi0X6lD4T
YM0yy2Ra+s+6jSxHQFnMdaUPlOcYEQELUv01iFdtkS1IxbwO9DAXkhNj4dd7+BTtWlyCLww+iNpH
PqXGucK6PlU8OkTJEizBzYNf0XlFO8oNpwJfyI+nrPQ5Azpqx7WdP2v5/XPloxtQUxzIu3RjgW84
l+cMmslg99dBO4q1Vk4Wz8tGH9eCGLms+F8JYECAIWUkKHjti+BmZzYUAeVNxmDBUEjAL6XPZSyi
I1ydYAUah6Ez4GpVVPzR+NkL1S2S/U7izym+e/OvctKGHqldYMXtCede0NyU1jPg/MBcr84I8a3S
Mxif7pn5P+qKOJzj/1pPS1s1GuEvO97a90EB163HolLsee7Xf9ANlZ/98P8lrn/4ZYEa1UxgH67r
0hjH0tSa+Uhy5JBLtn9MMrw6XfardeBPwhrxt82dNIcUKwV5DDDEkCD+3j/mZgaeXfx3IaCv23n3
otzwcph7pmTeSnPXX410sm1Ovp9TuFtKNc7UPfehLR4V1Lo8xxTdpjrLISZ+IWkKwIoS8z0aMJL7
pCp4Gs95GGwGXb2NQ/5SrWZPIz+OBLePgscqTOTSuMAPBqStLBNCRie28K0Fk8CyUsY3UrsGzJT8
X3VjP6LyazpVMQNmqA4m9ldXLdEE4+AoNMT4eJNIpimM+slyBaa1ttm9MS1AY7zXGNTSLQwfzP9z
36mPNEr+O9hHISB0UPqwhUNLZXsjGIG/JNLMWaUPmWOV8i3aZ80P7n54tOdqhr1dNqLUQQfqBr0l
rEdHfChGQzhJE1Leg3omahCVg/CI/Ae7GwPiPrJzUv9R3IO4tNQipLN5hiZBMiE0Q3Ogi50vf3b5
cy7IBmINQj9yu3rQUhqsBYwlPG2scURfiYNJMMxvPykW4VB760mcNmGBs3dMgQqUAQDVXo/bqZ9z
I5aNKlOWXvSXkx9vrgjyetBHqwxa/CdbxdjKg/yNc7DJeTtlisbasIa2wsvv1jupPgDCxICMKayR
bCX3mBkWOwgp/l4mmc+Kb9NiDMl81JPREMPZJ6WzBamRR+xlhRSpW8FKqlF0LIJGzinFgmh6BFq0
QkMnUHRg8exJbfF7fH2Dr+ji+keCy++Yz6JX37wD9/ekiiO+evBJl9EcKSz/ePtsBkTTG8WZsHs3
lWa65cgYn/FROkgJDDQUg9JiQK0MOFez3TqjIJJw6wHbU6Jg3bpWtlVgJgyW07qiFZ2zJkG6XVdC
3fFzQJFZrKWCM20yRMdm2sOq0EG4LWI2W2rliEvGeonx3QgMDuJMe9ou8yvI7r4rOrHHduQYl6Cz
NcVfe7FUfi46otgmpmIVEEPNaExU3ZARnPbXxBEkuG/w2gxCNDVCncuXfO6qPPI3/YHOJP9AUS3K
OIxQ/fM7ikSFFtU2Gs5m262UaSzPyS56v6sgYmItMbIBGIDe/pDTfxgSWgnuSPZvD2MRzN/1Umk9
tM93BJ/ED2VqxUjlnP7qvH0IYE27PXr94Tc/I+39xPsoW987hOUBz0DicAqN4k36YDGJVoJe3tsw
9WHAiY7Wr9I3DNT/ElTQMICP351JzCBpcjMgpczq4eGvaJIwPx71r6luioWmkL7aVEPkWqL6rZF2
LJQfPcfH38kBzUSzLALBVB1AgQqtVLMn46Wfy9wkNtWVBnhoeoPEbZw/XiAE3vI3kkdA5+uN5iRx
MVP9s8y/H2YMca6Yysek6yi5YHEVgrTYHPuu53r8JlejnhUf7iKG2Z9P80fW1oDvE9zoWxg5YyNL
OriYx2fF81wbEV23XwGvSlC4YAtfeQr6aOROFeBnUQfk09DIwWglk8GR2EGcRFSVMgfh0k/b7NxK
8g35x3oQdD7MLUpBXDJVqwaW4Hd0eWG4I2zwQlQmM3kOPj0yq2OvaF73gfj5QuE1Hmunx2L2yrEr
gyxfmqrlcegS9/2riGFz9txKgpAgB0P0+qHapQvuF1eU1R2ZnGytS01LEey12OELrpiXg4Vo9JYy
mUBUgdl8J7xYtXZ7r6uCfADzxRJuG3mS3DDdHHchIAUhQWpkdzGdSwJL1K3kTsIlOAHbkAocGXEy
7Dy9WilZsbZ8rufMUUP6jFeE7ozfv6O/fdHlS+ZlibwtlvNDp6Wr3OjULFccPhARxOED+kUtWrQ1
DqpvjOkw2dgGfPGFUtwUyCOWa7X7Pjs2HYWOss/H2XUWaRD2tnVzXm3dKnYj6aOYk1zjkhSr4ARF
E5CUeZYaO0T7LuR+YEXC6zcstQLI2J9sJwBiV52h7Q4O5IdMP1PJsAOC6vWZ16h+5FxUjXp5LD7A
imlsiO+jYGpweZWmSQdEx/EPa8MoDx34zSjEXdLxNW3HqLMnglk6PkvGRniqoeLp/UemcgsHCABl
YOQNzFqdOp8r746UGhhYWLvHGdf3jJnJA2Xm4nVuSD2uIQ2q/oBtkblfpm1AZVJkKjDSnjGD1uBH
y4yFg2F61HI7PaBN+EVFg7bgCoqRQP6DE+l8tFgYOLSuGNanHq5o9zc+rD9hDlNk071IEu36LsJW
LiYHd66fLofI08KzqastUXDaUTHxajSfaqSz28+6Ca3lcvmkSatU7Xv0ZrAreWP5Rev9IsP9Iy6o
2rPSWuz8iS/cV/2sIVzIY7RWY2pTnDZOkkn7qPyRE4PBF0LCJ+qBkYcSFNkT8+V1+l0mBbwcFE93
Y58ppgesHxa4IYnHvlqS+F02bihTxTKnEDHxK7IqAbVD1hEaRBrLf2mw3+MMFvvz1mUmvjZqAu8H
CYsRRpAZe/gOuBiE7gJBdGGf9/g9xMV2+Nvo9Zpd84JWyG+69hN5KFPTrzJCq/MdggkDJ1+peFMo
a8ibiudopcOgwEgEm2ag9w+ZxoXCR05wAWYgWd2ka0pPJFmGJ+1cz2x3LKKmpbwHSoTgMQ+H+/kO
zdIUl/EowMV0IKH1u3fPEe65di/0NtFnIznd3FwN+D2sYjHsYYCAfNCXXDfk8z2r+CcyV+uokNGE
5A4R2IlBDZldRQJw2gzmT9gxxrayumoBF9r/8oNh0Smi3TDzDzd2Ew7RPMxcxDKphkPrxZwacbjr
aG+04OJP+ejh9E1eWVHoUhtAUTr2sGnObAV13Y5HA0I6KsPCklA54pddZtKsnpaX8G+/CCp6SmEs
YxtwiMwArelw4k5woLTpaf/gNCKjexGSFWDHAz1nAPKUNlNczcmp+lAzmiAEDOpc7Apgf5wuYTcc
xZ3W24HALrUQ9vs3e+he9BBlBShh3XRs/mEi+3HzERuDgQ7rvlSb3mVL9HOiAYPeObIIbfD7BIiz
w2b/OfwPqChKKzgl9w+mdccdeHCmNw0whv6WVrrxTag6mp82sM3gTL5WEKExOUwXNuKiyq0uc0AH
kkdAIjAUcJxVFqCsvKDbQj0Qw91k94VYYzYG1+AnmF2olcosDU4Y78eIxqW5fG2BTSq9oMKpDoda
3NF/4gCoP7aOnOnISYTISEWaFwOEWjWrVOE42D2nF/XySSXXDIGSiejjUCcTZyBJYPVNeg17CJOq
YViUl9yAvRHkAuIulwV5eLemGSf1U6E03pPLdBFPUVbPFF2JbuwpigFrCUK3JxIlLJLx0m5/kJps
0UxDOmmCZsftxzf9g1rSEjeyIpfsvWYqAb+Ijaa6OKN3b59isDfXkRNCkhnnX9aKPW8Q/Rqo9VJb
EqMqRHm4olF7h79mRBV8uqtdHZLwh3+8RhsFYtqjzLo7Y0tnty83ZFgekHKPhEiz0YQsIzcDf5ab
r6bG2cz7hvvc556hvjNENrJ28TIskSQQPXPhyeyf+/3vN5+jw+imgf4h+0ASlITemCSLvhuBK1LJ
s5lG0xgyHZUkIaL7DjkRv8bIHNFM/yzgbButz+whHwwbtRcfPv7LgOih1CJDh79hcLvJosgDkcdL
pHxzZUpuiv6xAE6EbHRd9y3Z/pN5vEwyBiJ/9rNPOPDKUxb9RPrJEvSKwXKAZhkFVnfxFLpeaRu8
/lskAeyoyrjWfJDXzW4VECLpSydElAKKzF2GEyG5OA+tghG6xzB3oXDzniZYTstwNNCKMHh4h7SV
/ilrq7fpDbXloy5OeOBCfC3VP0FT7z57gurLinMMYzpH/2YrH/Acvfe6NWMw2OJzd60eQ3tD6baQ
CSQ3OTXGQL73f0fTHk5BcahJRn47KXbd0yq6olVL+gYcrjzcB/A6eN459tpeRMnplqJQLZP18vTH
NPc519/6TVr2xrk5hBRf7gQoR/W2tgKN6rKrYggJgYyjY6aaXk/uTHLy4biyKxc1N4NJQXatJWI5
q/GWKzEUX6x3i5iZA8+EKhpO2G8dwuBH+D8D18JUX6YScKW45ke06iykgCimrpWbkKGJsZv747Z/
zMiV1Na4zfP+NefJ83muL1RopYif+vOiLsO6nNfL67RCTMMA1MGauvtAiL6MZTJPR0oFCrux5VFL
iAyf2U1b9fNd8T5q0nvVhTZA4mhHJWMuFrPiWbshabR7KQnto6QIAUHwhs8HpW/CiIocrOP9l+Ii
ZV/ctRHW8bPVsDaqXQn865lgwVpOwx3iKpZS+/sHCD46BrEbDtmCICMbIYg2yo4swDpKgtT69GP6
8yFBO1X0EQKHb1+xA8wt95ZJxGGZ/75BMt64kumymh1Xi0Dzdg/RWpz6qWbDZK2Pq3NvstI8Prnw
UXI57FwT6LCbcV3LuHq0m/CQoiFlOOWLooJYxN3jD2hsOVqJkKosvk+yJhl6W0LL09lNcoqcR3Pv
q+R6FXCHIcSXVMwBv0wKlfRewQv/gPTB6cHCFSHoqJ7Iy54QF/s7pLSTRgtNqTypVOn/bNOuSN8T
eJz1FozbJmtQo6E93nJrOdiE2GpeEvgH4MFP6I70hpTWo54bkXpE+dx0ArVYhXBSHZDGRmEYkUGP
70Bdc75cY3EAm2cQRDT7GYPZ/KxAuP286od9BS7uCT+yPsOPE+WRsckUeCucE1aKOqF562hRFwmZ
EDru68Mfeki+ig4cuuUGXJ5+o1yBfRGLSY1Y42z5c2dgt1nAdwvZYwJ9oiS+gO+2EwrF7OZWxJhy
ZamI7My11DsvjrPT3YOtGt8+OJRT86QLwR9gizIvvpbMDVA0iTkWPkyfCeilSz+fbLyO4kFfTKp4
pAExsGbMCTmTOq4b4/S6ipt8i8VNYli67aVJyOSayiTy3LlIlhF4lFkVAaHlI/Z/OXr0idbYLJvG
BQk0Yz62176AukKSnDBdooVZYVy1DLZT6FUC7oHDFS37YGo4ECrUx3wqbiN8vlDyEiVcHEbTNCFR
oWa9cHlmbmJsFFfodz2kwKnwpbQBaVPZzWHBRDtrHqvZyztJdwmHNygn9oY9DtniCry1AShF4EZ1
7B6GFeQzNjx59pCJf8fuOEixLDe9bVSv2jYjmG8E46Pr79ouO5z7Y4THQ09t2T/AoFWBHLdTuPms
9+oTQhGTQL2E3qr/mbnJD/BwIdH/Y3tmKha1X7fvHYo6FdWsBnAf3fBiT+fYJ9PmQvVw8GoDPqpS
VgcbhLuH8f6VVg7x+HT/P+IKphkSo5qL3CXHTckS4y1NdwczQJwXFOo18zV6TusbkM6IwrIGzNI3
bsIkVDWV8pZNJRbSWn6vv2JUX5FamoJy1H39zuxuBnmxi+9LobZzrR0ZkCzfzhr0jm/J9fkhbII9
HatMGsc4qnISD+AxvfN8ujna0DK8G8idRy/1qZg2TmAkp7jc+7seGps2NjbWyuUEa2cHpu7Jki05
RLjrLG8K0QrXLTSmQNNVgbHUOggNSZx6DMh4mYbAX4q57Ee4ODXPaawnGHGMURaSQETvGpVrqfJj
lvCt7GO1niR0hfPbJJtRHHHfLs3CAMDOASqgNsWpWow9q5yKrZkxqxxFOpvNRxqCVaS7yrws5Ikp
5fsYgFZ+TiTKscgAzlaR6I188qsaQl0BkbOVSEWEmvZha1m++3+dcvS6st6Rod07amUgjAT/f/Lm
lQ9YEZWRr273zoDKxOqtRiwayAtRlD/J4U1K+5eMRni8GSHvo20G4RKOoK4UiiHuh9itYqAfFwQA
420wUVC9ZQ0fvYLAHPf7ix+qR4E/XRI9e9CyAqR81dryPNCZZTwEM8Ca8QrZARgs+mI8YHrUkWv8
CLUZHJooj9s70g1vNHAoCBoIuqWBh1vMcoo5tufb+4i3ESAkTahlTaGXrwuLEkUITj1wIU9dndHm
v0YQpsn71NJ0/2FnFMLF4SpGM2RkHM1Z2eEMmmuoMeeG0WEKPoriS2baMFCZ9DSGXXiN4qYHYsas
HqsHw2D9QK3DHlgx5FQkZloMRw4zg10CU7gDw3/hsRBf7RgaETR0IGXobCFcsreTwOVQZBM3qU9Y
4OybE01yTjIXmll7GBGEVByF60tBgmR6vQiBc3YluijmL3XTCuYLZ570oZf7Csgxqo5t61mQCK5/
62ocw9WUWlA1egVA0qPpoKD4Ux4RyPPxnDKAOVWpAgEKQ2gB1KNqOo/eAIqcaYU4e8CylxShrqYE
yvh/5edpdG8AGGc7JDB6hk3TcyrT27/wADUU7Rb/IAz41Qb1KPfBH/IQiSk9ltVZq0QJ2FNB8CwL
J72xhr6ZSuAxfaU1CjoG867UEkguOlwJenuCpoIougLCAsbqGpjETplwUKGtAfdnd0ccCzXFXYdY
sRNYqgI7lzVZTjfMeSDTaB6V4mzemEUe4EH4L+w3HZSRGLrf7kVky95zZBfv1zFHGqN0T3f0tLuQ
t8pufVkBc8HiFvKdQFE9upAdB0KxLS020/xnJdBcehB5mSrD+0lgiHtynD2D/0IeX4J73QC+TO+v
eppgeVVtDQxjCKCQnK671LUYi1XQJ61Jkqnw4dD5Az04oHrmfzHwAVOj3+oVS9cV1P3Vi6iBOLXS
GqcIrW532FyO4sJjQwxw4BENT2mGC5NttujR2p1+cqt8rxIl02tT9ghOKLrFEONODNRAa/8Xrk9F
Rp7q0i2SutS39GXcnZqAIL9i8DRgHTEL3uFg1Yol+bpNi612VDllkqrbnm2iQyTwvGzr2t7P6VCs
4NkfXKGqVHlPKMaeKqIGd2aqOqdALvs2hu9G8XyR1jJWP5XcizrnAl1+2T0F/mSKPE5gP3n9MXlO
vOkztnYW07mXPSBDR8TAz02HbsFtQhOXO5mEht0rdEmNFLCO4Ri42gFCWLB8ITMzOFe3kiozPor3
hOGrUsQAnTc/fmxeuSOiZlOU71v8OgFhwf4lPyFIpx59WwBolPxeuGweXdFxqxg6J7P+PiCYs3on
WwrHByNvPQ6L8YgcNC3I7bp+ZQF8b+/Uqxry2JG1xgypO9RLjBoS+MeTC0QOKaIWZJigWauuKOYt
svXh4aWSnBEJmTagP+asCMFG1ZIcZrrfnVgcCKxuLdSjKEBnjGUvdg/osdRDuzVQ0jwaAS+iwJJP
vVkeWp6bToX8wzXvrCSX889yuaClPsrgZYjPs2rskhXsBVtcZR9pkfINZ5Zc8qAbQwYuI5E98Omr
pwy+L+PdG8b5cZU69Dar6mP0b25QxzeJ/FfXjgJ21NUpmKyq1FVGn2O5Dryne5mF2z2LDnRow2qD
R4DBAl60EpJ9lkGHY6y0FD4cPRDmvaQPKlzwYD4EMOAr717c4Z2IbHBnT0PDEqtRvEDLb36T8pn2
nvoKb6UnTeBDSDrixd8h/lvmiKSvcZVrWSud0DNsLUZ+t/JkuufhqW1dObnOJ1Yb5WVZWx7nGMQY
wp1Lhxp6Ag/dq4XpotQkeMJwfTJwHgYQhkpdCUy70WHeuFMp/G88sOF/6a4WvQ7RjisvCn9U4lKV
wLg76MlOXOQTpdzGVKJMQLZ8iWtVCNr6qaP+vb8SR70uHzVBK7kFeTKzAn0XJNH8QUlHYNYaH0zq
fE/dFag9bi/YFIDxV5t4NMkeUhv3kJZL1qoMi5NtIxmqXjRu13zy3X8iYspWo5RQL63WV8GELfvi
ZuMoKyhveYKCJ6awc9pmhkYW6qJDIUkmHyaFEy6EUwu/648BI+lTxt+TFXQ+azRi3+SGbIkKpbtE
YCp2xWuDJCNSqf/VdRu3aKaPg13hWByYszvMMX/AM/K90YaBB2nXY7KA3jFzQPDW9PYPAhNSTdMc
ucnWhbV5VURlo81UjlSMhZzguqY+sl2oTHYQfvcfqgPH7jY+ZawxY4UfvYbuNfUZU5eYooDu5GMK
8C53CrgqiBo8WSncX6nZ9yyum2cVUlscRyS4eIORasujpSgXcjRVurn5dfPtmYQik6FkOY9Sk2Y9
CHxXQIp9AAOxL3gNTYsW3KY2aEsnY1C3sTGhcFgRoveKyIMn9RFFUr8uV6q4IyQ6iSa6bziY7idk
0g4WwM7FwGO3hE/euum26yK7RmoSENWjnN0mpA9UGMDqCDpUzljQ49zVPqVh1OAa+m5XR0zO0rLP
UDxGC9GDN1wHeG2fk+d2YpDZukyWCa82hYfW980otfqYHRWQfUanWX6ubkt5/rTs9v+BlaMsC+H4
tPjzFVuyNKw5SjNii5Q5HrtMC4YZZr09AJ+uS8uEBcbD3vY4bFAVi3gLf/0yekg0q2MK1hYvGbTX
fMbI6B4PWdhBcBnQAKyyibPJu6RGB7rrzb1yssKjT1CSjWEVI5hjtJgn0EEE/aLVV45APBRNWizd
zdU3aYC1s2MfD3Tz3Qfp5f+18QNBrWuZn4tt2WP7Cb5xV2KXSAJzV/wJqgrPODSI2TIxkHUWf1u2
Y/J2dQIesy0F6hgGOVRUWZ2jL8T4jiL3m5JQzO0LYZpFd6ByJgX23WmZp/KB61KsxVgirNasw9eO
F3vm5GuaShufV+YGK4usMUJizQ611fNHgoikMGd0v2i2TaATsVtp06Pw3zxGjVAXyCVq9/ROZ/Go
+pUnNK4jR6lRKUnYcD4p0kvCcx3oe4oGADNKjo+/mLV0QRhn0jjxJ1fu/rJ+CaoJDOdyWEc3RSj8
raEQkLZiGaycUkqyDZBtkIIYB//2+3FA3qI6diaCuomNAzYNrNmW9jV65VEmf7nVVBy4ODPQyEhv
5BL5ptRH3uRo6gi/FMe40IiYNa5n4LmkEehucYBVj/I3Lxoxr62h9vC5lRhXVVPO7Va3vOeTnL4U
c4Lf1vpkVnT8kfpHItlWa3oNKy+RaqALAdt4zGtXgcML/Sasy2HbOBwAOAyK8fkiIL047Q1Dv6jq
EVegAXyDpEwUuaaMe9DNlYnxDyPuOntItE4rQlfQQFm7FaO6Xzk692JuM88udO3YavlSDtF87T0Z
SJHiY0Ir4Nlr3D7affxz1iwXwY7juEpYHh0vSpqdnc0EkQX+dnSnWfZOWKfpFQw1BtQgZH7Cj1yS
GdE/bUwXUfBPNuh8HGk+6JqBa/eK2FGP9Zpb6gwnz3ZOzmx88OmDJbpE/xHqQVArieyR3HEwITAD
Izq5unrn07jISfyIlikC6lcoltDW7qkss49lYoL9UIr5K8Zz3Dcf3Hk5vQ1KHrr6yhkE3w9irZRE
8swATD4Sj9JcpB2SGl3tYq95bS9N84/sNSf0HWe3iHHf6ZqwW81OFpAJfliBm0MwAoRYJ+4VBEwk
irZMpciyELVK4WMDSXUYfvx7uNotDgrUBgpu+ot8rl9A1iFN15od3OmMqgd/1KG8jJXRJED4JOQ3
CFRk4TVkYLd7uN4KA9vbfPOFF4iBLdUgFm5sDI7D+mDc22HRCbn4oh3Da6gkeW00N1mdOG/CzAKM
HeKx6hwrgeW2kKmdQn4Xgle/VQjLHxhemkfR/KpjwD1vmtivTtgiKKEhCUdgrhpkjGlHg8ERtU/L
itvs2SaYhj3ChSqPZLUWJLRX5Fv4nN4VxTudUnwtfucisEbbUC+sS8DdiHQomABmjHGDmsXW6b+9
bK5dcsBIJR1tamRQKMjDAv4ZSwg04E3/UcdGMBBLM6eX6TRVy3mqz7yMmNIbP+zPv7h+SN6CeZ7U
/qJzdNttFj9VYt9BXHu9S/5Fn54D+4MQK9GA/uYIb3rBZj7LnTdCC9MCBZB/exk4M8irVniEnoCn
x26Nl8QfvhAFoCDg3J2WQmaQGDR1XcZlI34Uh09iQWqjnlPIcPEEFwETPWRKtPxv7KJVlgEMYlJT
jef94jxba0Ww4IBM6K19cAMbsHL9U4vyg4edKESf6/qg+2VuyMoSRQR8YlrwsBY786x6MOlUR9L4
omkTH9tPUqgWHAht/SQkT40w/d3+ai7j9NTKSdXrZZsS/WzZiBkwpuewh1FKCeHqW5fX4wpTw/Ej
HJu/s9WeqtKlkh+vIME40PSvDbLlttEMt/Tm6YQ2wIYJORKC7sO5Mfy1I2MQKiuFKUGc3KW8mV6s
m0F2fTlEmXvacikz5IhehRsM3lkhcdRj4W2yOZkY3iw/AGtFMz9ARIce6Fn2MQIK+Y0fyI5R8oeW
7u4Os7ZdzvaWGG/niVb1LkmQt3WDcF6mq7HWMR54JHug0eNXYA4YxPetcZsxywINw0Ji41Pn3kzf
oOB4GhwsW34SEvq1NV0PC6rGd5gUyBSm/RPV7rgPywz9Lwkz9O60QzTJUwULpPzqEJyj9exP3zGz
8NbXkSVB4XekI73uRPvaqIj1chle/v5/ID2vp01pbPOxMFOjbGK9y7+TiSaRZA7rs3lgdY4jNyD9
7HU6VaRsM47GpPEq0Nco/e6u5W6aCK9K07YNMLH4wkl5dKQkS5p0w9B0GufqcP9jQPRYpOKwTIyw
hJev57tR3eK8zEa9qfqPZ4PuRuIvBLeJ5My6nSQ9GuSvG+o3M2PUdUWELk8zrboNXXK36ELqPVx1
kixC7fVA5oEA6cij2iVkHmXiXxFhDE2vGJgmCFJQuv/ckh5kH2NUsDiLFTKVV2EZsRWQU2dIM8DW
ijeBZPNVfaM6z1wI6AxNznhWyLrDus43o8+oHoa6LhnU2iwcyGU9inP0Zl9canvwgLuzYrhVv5++
gYPbQlcSGXsvQiFP34vF0SZTqrmxH9B9ZT91nxFip+Hn4h21ANdls01f0Snrv8W7B0vxMlMXJpx6
ep9yMFtFwLxNbXj9aAnCCnsvOP373tRtg/LaM3tvA6LlSiRAF9Je6wHW9W6+4A9zP9Lnp04PeIwU
2aQviJYTzDG71XvIhoOP3t1HseLK0MCE2PUKZuIvBDftxAxYkP+d/BRme2TlwZUL3TM7GbBPrhVA
cI87DVaSxwptwE1qxH4wR1DlBBFjjOZ75bXurO8ZkFmzZhYpF0Y/iBzz07gIHWxoctAHvtt4IDuQ
Ubzy8bhM75gwxVN8dqTQ75vcG7Ja+jafbJpvZIpIzJjUB2Jv22xboj98wGzJjOEhw+hNwdL7vvAp
6ljeWRBj0YB7kGZqz9xN3qzq/P/W/azmo4QtyvOTKRxfgMMJvqr1VqxX3EQwIvJY0xrWQHlDJ4Fi
TSlI4YIweDjkKClDFVL4YvBjb3GFkeZKM2C2thRg+1mGOcMK+FQ9FlScfF79uJDU1UJfyrK7JCT2
djjSfsQNRATNlVs5aesLZMV6d24ayPd3tfnxu8dZ3atsf0Vn4SGSCByvcQ0Wol8DR+6se1Jtv2ew
Lv2Nw09NRvBi8Pd3oZAxpb1wtvY9GW0B0oglHpyFqcgPjR2ExkZyVGG+ATLMbZ00S0JYtXVlBvrS
v4CnGH1Jib7ViatDUD41AGZDZgFR2o69ry2V0bnZ0E4h6gyjTZLeRZh1M197B9o4bfUaG9RyIMyn
/h9OzurhbCC7Au+2sG00Dj912PdAnwknUkDOnK/L2QPleZPcHljtU2n/xzcqaKoaOrr+2lxh/sau
U2psBB5Dq6yFfpj3ZuFTdEbXe2EeiYlOlImpFls3QqPdFBq8VJvHdkGNiH9MHy2DUvKSnky2zzNR
lUpoDb/HNQWPuOwhGWE6RTM7y5+vu1T8JG2nsFwCEZ9JYzzYX0V9g6OTv/FvxxV2EQ8fohGt/BVf
7I4X0Hkh+57Vv7nBbrx0D/fecX8x1YEJQm8NG/BCrBgyZlNUjpfzQrjJrx5O3cSWN+llvQZrpDba
5KJ/dTaPe/BHQ2K0XtSv1OJlEO2nI6b+YDtDSlgqgI7B/aRYGR5grajqlRc/ucQUGqUtz63+1oog
TVmt9dHX8NZnCBWGv7oGEJuOln/uXlNFajdyjx43rcCH/iQ8KJcuJxJIDrRR1zA+pTHB5pHM7lZ4
i76bHEZ2LKzB3uwOJ9nY1Q3l98KiCBX5AwIWVQKQ9+TGeYJdqMwkPPYl3yPd/P+ryTqhT/TOh2X/
gOwlje/gzPp4crORCoE8cIdd4pnw/3FjanKnzpnXkYmq2kIKtAyF68B7iEHe78x87WR+FnbYVqsN
q9AXBR1LgohSxCrQErqgo4LakDTco0RpaswKsVcvDNyU108sl7fWdWlJkha3OczLyNuqceOMaeIE
sNyxL3e3og02CDNt/EAnwo66s2u8aVQJB7C3mYqdQ2ir3+v73g8+w9FitcAP301/A7WtKPqbr396
sPea1vng9CnKvlC6eRPgR1APg/cXvUhE6eK6oKJBGeYXzVS8rqSQUv4J1sAZdpMQWUiYJX/Af1V6
/ELfL/bqXweKoBEjCkriAKgLzeKSwmXKa3okeJbD08sz4VxemWjVbBfClrxY69psYMHCaFqdE4XP
qwqAOvNnNKVsHuaFXB8wWZkybOm+DxOn87lu2aWnetlXouJdHOFz0vcFoHpWqB9xf+iVvpH4inIn
nqQ0iVAwyOe3UC1k57ELf0gH0ByAqNrETkEaNyZbKy7Y1FruYI+aI9g4oXIJILWXIr4QLkwWeW1O
3a17Q3xpAQbWXw8lyWsPTzne9RuG1dIpLUdIP55Q0evCfF0SQ88a7LUMCmQbLwuxRFV93wZXf4nA
y9QFDUdUIFZK2QP3ZpC/YjcnQpugqHVs8YUHPI2O9wOZVC80BnFcS/z2gu30zEjSJBpQpEYP+C65
n5WISvJn+t+C4KsC69te9F/HbU8hGGnyLT3NhLNHoyxTybVpaL7qqegxGzRle/00pRmOwNts7wgO
He6qK4/0h3P5679Qu17w4i2P1MriW56juX4O7HNWFbDlyQe6TxwDeicqS4C+gBobvZ/AOGcGbhoI
zwo2jgY9zRiO75ta9na0xV7IDcFhxDInsWj5bAdUwxMQ78HlzOrlxfcQzXTirVEQukjg/92U2Ww+
a3zjc1r4n/WL2WxjhLO0GsMwSIa3Uzvgj60og7ktlcTAMrJjtqpZMPWXdv6ui5Ac5moGneiw0hv6
zYdZe6t4gaLxwLbOebB4LeF9Oj0AhAMwxE4T40/tdAggGW/gkf4W4JCvyKnwvCxcpxjHL7xRC2wf
PxdvidGhHMQ3VHTLkVy6TjOl8EflBabsENy5ag/ZuhJwLoTpd1xHBmiZqidEYBZZkqNqXNhwGNYW
RDIIhjb7R+/hAL3JTN5cuTC59WWv3dieJQ8++ONO59iR+PyGXupVLkArZZYscD6LIdki8sMgSlyt
hYr98Dg/+uknjKe1WjtsBVNimUtqKaCkX8/TQxywl3sbo4NtqAg4/+Nave8UqlhhE2RKwrH3MiMi
ub+fD1tRaIQzQfSn8jOcHOKlS0y8szaHfgI0GKW5NJ50NKT/4hJ8Qs1iI/PfchH6Sm8pl/Gooqqg
QZfPwReFILHgxV8bZl490fnsoka08YHjWWnV6qAmSpncsoDkZ7M8bOC+27GSmmArLfEtL9wi7znR
unYw3/v1jip61RgNPw3lz1J0/NqPKamQJMjld7Q90xVjmiWmYk81uuRAmhEd4T+z7WERfo7YtIKa
GztXIRtJ2ZP3AOFqGgYZaQzQQQUghyGtxkehkYKOvAx5AxSg1EX6smUbD+k/A61KFsOrzqOYhyFU
3V+cHeTMDFbQmd6PXOnFEEFL3Q5+Pyybwxw19fuAj4rt0xPU0TXWWJsfIZBFO9Pos256vPhIgP3T
vNqLcoyjoY0a29CA7DTN4obblfBRaVdsJmuQGSTqmYyo+YGfaA3b0sghYZ4I3MyphOXGgvQYNHT4
TYQLxWkNyuIMV9Q+JkdKDblQE+6tH4HhRtJtxNb46MuywS9Zw+IGk/7EuXWTg3tOLy5yasEdp7GT
IbTab1z1zL9w7EtW7TG82Kau/1xZzJ4Q7hZqZMrKSs4MAOew7zauIb0Pg+aW2YcwuTRvGC+eXXnG
S32N9F4OAPhAZVcjgdjglWBdfUdkVsKklGR6aNKxjfKN1nE17EfBi7u10ggducMmYcp6OKF+ZUzf
aTq6ccvdfnQXF/u3UWFDnvchMx4S7/W0R1pw/lo6BqTmWUMUNL3lTDTfL9EJi3BxsnEkYGP+AHAq
bMPHx4I8wNBpYZUKxG1gCLKY+gNprPoYvRla1FjDdGQ6vUpbx/csCxj6mdq0+6OUPygddv32oHrj
NLRElwfvydmKVux2LahTXXYzV/oIasv4X74nUQG7jBd86z4qlXAfgCb/zKQNqMbaVjTGlfAct7mC
7aS6mfb9stinAR1aWtbneRucxWQD7fwXOP8IFzaOPyMZ9SKy6lo+qSsHZEGFgSOCXdWSHaMbZoIW
LRRqz9/8y62F/4s1zJbif0oY1AKGzqpNl/HaZw6HPM5psoBW4qW1fNVaOIPBLgF+nxieHxFZ63EI
L6eErdCGG9y/89tksdS9fy9you507eGE1xI397dlhF4ZyDTR1Y1Lda1rQzOdCFrGHDm+O2a+mrBk
LiyAWxgfftdZQ3hIGNA1xZE6UzKDq/Rs64VXw1CW143guq+KoCbyuIJrt5ldaWBsr2HKUGHpw8gE
V1+S20TwrBGaUOf2zqMxqv5IMnTVkNzDCIB0IDCkxqgSTLW3IjeVLDsKSH2RGFwh4ZGLIoWtVdtz
6bPl7V3JaQkABS9RFoqsikMFIkLV9Y4X1WfsPr1QHSKpZuT+WLChTxlhLw21DJyOUX81I+yEI46U
JGdVZUaneiiNvSaOOeCefhhRf3//RrmZWFej7vEPqHW0Y4MaCdiEW7z5Erb8ChCGQG90pTlWa3QE
hnPEITHYDao4aijtuWjQlBMMF3RO63FAcGYNrKc1PVg0VXnOU6YReqrCjCqYWuvz6d2iSTGFK8Eu
4OOvTb0gVfIIdAXhg/nqcqxy1Biffn4407vJE/XFDRU4NaJSspfvloPDLtWvOfBmkBgJtuUk6S6z
cZN9qLhkI93EokGi/lbV/BzjDTfovsgYoJtkSi3dQrmiXfSmvrPxAKdAIunwYI/7xO2YyyadG7tZ
+C4UV3QnxIEnPQ8nrhkcC8TcJo+uygPQ+bo9IcXj6ernle85Z7MWu0GKh1RvCvLG9iIbTF4ExTbw
/r4Lr3qqYWxGwaOrx6XNSgcSW4O60BIFjwe3+rg7i+/HIweCE3GSyBydMaFRyhdgbSxoEzTSq5eA
xHtZBxXGmM1/SLEomfShl5w68+iKYmEuEGirv83+TunR1Mp/Wc0q4KIyzeUZy7rsdOmuDsc0uwGZ
KkRwJqvlMK2N9gTaLpN7U1+BMysW9O6kBRbzXd1bZ83WsJXf85o2teKj7anNXTWQ5f8Z9PjCNPot
xYG5I3E4UbCaeUkfruHUVXanKJxsri+i5z7lNCRY9GvWWfGm2NhLEugDm8dXRHJb84bJynw2CC8Y
qtpKOPQLSXUK54r3IZFXwaPkfvZbTYqBcSRxLK0dJoylsNCveLmiC9XS+lkNlF0Ucz9MYpVPBA7e
iYI8zn/OtUX8XdwP1/cIku9lxKImgAXNvz4y0UsKar1vF6O6Rj3vXuafzPyAvLn49Rxv5Tfuyvrb
/2LPeti8WAR52LGAGvAKT0N49KlHX6U2yJHZbVOh1HCWgI3mxYzGxa8Tz0ee4SHktbJLnMl+qrsh
NjAUsWlJeMLWNcUhY7GgA2jaY1gtApedvXNYtBkK0lMFrJKL7qiUSyswtF7xZeH3W2rC+n10YR5H
AXFS3IFlGN9aElsRPGXBpUhxMnj7TVzDcWay3EbHznnXg3JTTanSNySyDNubk3WpU5i7U6Clz7D3
Nvgp9LTJwaRs087814NtKHLmnscM8J43ntzcaRDMilvV29X1R+m4N/jxTr1abYsHoKwXNuirv8lm
+U9xPA8dcze4HleRSiEt1Uc0MD/JU7vsBqoaZsdqYVozC6MUrcV9/QNOwGpO8HormrQOC2SSoK2I
KCCouca+UHLEX7aN72w/ZdKnq8ziduCxeNguAKdAzmnPTSW6ERzcmwo+60Xj4kMFUi/zNBnLro0A
cL3f1rOgqNjzyLQI6owZgTMHvtp1Y5+jDkpE98xv489a+CgZWnIK5fI+CAS3JwBFI3JOT/9UZbh8
Wmct6Ojzimhvx1QKC7y24rhU3hwVDTr51U2LX7X3RK/A2+v0YBSodDBmtUykxirmSdgVXCvjY/X6
0FFh38Y5OKv0vafwuM3w6Bl3Rzorb39lhsGhAVqwd92sHxCPXGx2iirYdCknOw+J59/VgdojMGmv
D8FCBEDmRS2hjtGITlw77uVcIifgbmFDNqF+Un02S+M3JWy4rR7x+stTg8cMLPNzY72mtgpyClzk
OBvt9JMSw6WpBqIIgidmZIJWAZFbrqNARPUlmmFXDhmQKYIFfv6eCMInfuj0DTDwDGOEjTuA0fwJ
vHzv/TEMkfn7r4GeXnntAOHfgTeXxnxwHNZw2CxAfldHkbMNPitcDDUtGLrUMu5HOraiffUKUvFY
xbyFF7JD+3jInAWgpjmaMuQPpdc7VxI661sm3OFVt3NzDoMGCABPekcka+cvSria4c024RpilF9o
vciZA2ESQW8eY/CGebJD4F7JsE2iuALb7sc8I/u0MgqSYBr0etQAEJdxcEIlAo/VKwlfadG0N85t
ZkkZ3I+kxRq5rp0FAG7eqU198wvW3fQTdveNJM0at6zQyqzQDOf1qkpqDVuM47+4uTlpJ+KgS0xx
rbgt5BNOgkl+c8fwJKY1pBU4el9MVm0IBnMJ1VrmoJmEIH+TuxFOUOSARvmCKI9lgF2fPYoDr4iY
Gzg5M+bne8EylFyH3+V3oF1jvn6V9ToRp69YrxDbrrXwlvn8sc0a59SL3MUD1X9YTCpnCQAUYT/H
l1UP7L1yqCz5bR/Pm7ciH0wuSrY1KRI+QNzQOtuVtMODRXmlQhSpvjsRIZQOrj7jpFuIX6Z4M8Y/
AALXvhva7rw8FsOhTBHREHnDwSxWEwC8+6xcr7dgCwU4S61bBohGato63HAN65aIQKjuCl7v5s+X
Pi7akilF8bWFKAwV5gY3w8oqHs6+hlq1/E392uoQA3aN8SigZqZW8y/BOsTerPCmdffDmWGXTECK
9Cfj5Vrg7DK76Pk7r4xq2jtXg8WB5eTZ2XTpHcMbDH+efzRNCDV9KGi1ecMiTXTHQ6RbRfbPVk4Q
56O/IKi7+4VbVKtks65oIM1prxmM6Hw7vyJg4dlq5aEdMexehWh19WJ6wm7lOnAEOmhGa8xukdEc
O9iSVJ/xikTwBAZUdJFO4TrAkrNEABud2Jhs/4TFTe4WlO70hTr6IZFxgF4SRoJE3QFVXG7AoBnM
t/cZd0GlWmj1tM3gUkA54HRgjYHusCGZHwGMMvVG8UbaroeujZZjZqmRuIMJMWPOmMp1trqMNhmB
oxX+YwEjVWy41T4rhMPsG1KChG7qfCTH/+MaLX38EZAAePTaZrvZoQaRfpigTEs9KuiaJ5o0Tjf3
JwWWr4APIpJ2kR06QfuUx6s1ri89WZZ4nrMZdGENeIWusJ+r2xaZvS+PnhktYTuJ3yL7WzMS9+Ya
HU7cqTIKdqDFJcxKBhWR4T7ixxnQ/YbI5HiXuCfOcZfBkQljrr7Gm6bM2yXfNeZm6VTn/h+u/C/Y
ETwXJwyWW8EZy4AaSZRmgLKZ/EHrihDFlMI9gyYHgAxAEP4o975oQbsq68a+hl4WPYdIuA7mZYoi
K5rgLjdvVGHFLkiuG65wm1kzGRknd4nFMYs6yWUX/WqZTVbqp4FrPdFxMqh8Dus5p2eh/2bmIDpl
WmWkDP8cyVXeBhTZmVITc2Yu8HJ11ImGBXvts+vj02zT2UkgMxs1T3p5UWLvoInB5pv80ipXrxle
BQavlpuxVSx1I82HlUqS9hpJzdz9Qplo9BQVJ28ICx9q12ZPpllPu9l2deexN2r73jRwjlfOLCnj
dkzomD2Lyd+OdlF6fCTlzm6CP6/OS5WKVMR5UPR3mXYAPMynUwUM1CSz/000zvTzpSPcF2tRckex
SW3+/nk6eDNS0JfXxcBojkHH5fI/rk+MvgZqX1IqEBf0amOh8HGML3vQjkQYG4aOIcthx2G/JUxx
QwDmpL2U794g7PKjDGUu0hToliF2kRqre8gQxM3SH6tjRFW6BNg/HM7JY8PXAn4k7AUgCXqWCp3r
CbEqGC3R0Hdk03LSB9YfTxZ9wwVSSCivDZPAchz3740TV1M9SX62h5DHP1GEdru9YeTr0Y1EYkH5
pQ2Lws6XYJ/cqYRMEpaoeFyKhViStoRTVIBfKcXg/Tm0nO4F/jI01q/hhuh1fx6SzOW5s9WBxEj7
TzZr0Y6vVIX8PZbif6tcTt7SCR4nxZsujVqaA1qaBKM+cdzyodXhodBNLeAlRH78RbJisGmBlerI
rATh3MfAyDwO49d6X3j28Bim5XPT3AQ6Zn67xBAowEhlUhFLkfMSp10AU2x7IEGQKjnzgQQSMZd6
IAtfNuFzOv46YNjMMe5Rckss6uWUN4hDneEd94do4wsOXw7MOP3oc2LNN60VgYOL9/qLaB+3/CfK
A/Abi2TyPyL2tegBkKrl8DjjvfTGIv0cYq9HeRgdmHm8+8xpHj4ibrLa10HHKn0niuZjrl4BAS5P
wwWu0HSIBylJZXXUCCjiJYTUzllh0jDBn91EA5LroV5NZpRPrnehVmrXCeCKdbaeQoGbkwuPdyv1
5u/ixY3KNoNcnX46IHZIFtdxj/Vscqe89HLiZNCkgSym7+u3jKv+ZEqQrynBMJQoqaQQY1r843xm
0bRwCoHKUKHOh4s3HUc7VFNH/ClETKxAWLV8/IdB25avfO18CdrsclueaD+BcXb5JmiohjpKhgWJ
3O9Z9nmJG08+7vXMVpzx0G20ug2qVqlmZ1QOlNI97UyKZ62LPCZpcfeB0DJhY2U3DjGh4hH5nUub
Nw3r9A6l4jS68CaIQinaSMSfyyrmMyNe84DJwB9qXPa4Ww5P5X0f3isKAq4svbYki+dyou9A33Op
679xor6jA5uSI2AWpF/8bFpV520LoNE12eVELqncFjpfaRgVdwMXCWEspzWzvIX/JZqku1eOn5kA
B10L5vLpChP2lbWa41qU+ZJDAwqQzzmeG7dnZBUeixaHReP9Vwen/phV34QX+Hg1cbQD4zuo1qrO
HWdw8bPmIAa4M4vF9kfpeyhpvTeTstrrLQgJrSYfI8nVp+4jZMPzqg+PnQVdKmK7nXj9Jb1aKa0q
65Sc+EPc/kYS6w07vc8YDsXn99XHuqGHcYS/MFpjsfpyKAw/PT2fTUeHcCKhgGJjm+uAXFkfh3LD
ka+pj42KNIFqVA9u2iXBSFq09D/mBotvLb+m0EhyvVrUqRTqoG+eW6F/d1OMsHu36ZovpH2FITMD
GHmIlwXkmnUStw5LSTrfcpNHOEc/78tW8ITFvckD1zxXbT4dVpw0/KKddLooA7spnGGR/gEnDbeB
vydOdpOA5hrn+EJ57tWgUw+WYGJPt95Rne3poJltIRO4a4Y9jmZ2ykZ3EmHb59mfNeTeiI9k8Ccp
k7+Hde58J49GO5kWSHgxY9FBxbpZbPVa/UTvkflcV+f0ELxXYG44fP8mjDIEysmnxsC03+wCU/FM
nUS0LegC3FW4o2+m+8ZIajOdTyqmB7ddAU7JQz/RhTCmTGMPWRN/dxu5/XAkPFm/cUAmZDrrXZl5
e8678kRbr1sPFfkWv9Pw+azCdhn9nRmd68XGKUpuDKfL9er8/v38g2SR4UrBihAF6Lj0NZv4nD9f
oJMr2g1unEyprHvGN4HlCqvMkAkrkKR7BCh94zwZeDb7aswUcpcIimuW/6l1c7lbVRuvMnMD6x3X
lYmi29yL7Ygicjon+3m915vX4RObDloHFME8JQAYGyPat7+C3MlSQcxWgk5cImykh6TGIocdXBUk
CHdqEo/1BbJgI9rL8lYUKOHeHNCpS/foq3Xmkzp95JffgRBdIKy2j7kj6M0ZR8OMA1NKsI9HYaMF
htR7jMolxBliXRpnoA8GG3Xh721ZwKu/7FSI3ZGmka0Au/azUtZH9X/lt4RgMrMAcvvnoir5q5zI
XVXynLlQsw1uVntDe9uk0/xcZKiKgcmrffbBKloxNReIn5T9vNIiVevJ8x+IGlp92omIx5Hr7KfJ
H8iiRPeyNx3JqDqR/OTBV+KJtqxEDzUvKz4FUVyVigHwLohSUbuHevnZ/wFz+CMpsi+oBsA2+Qaw
M2ZdaB57w3z/7FS7Wny8PbdYr8ev22CDy/wCigP+vJ6FHB6EagJrBfZz/DYkstYsCloe8SHDcyuJ
bPKuoBBA0imw+BDjRxDxnAaOdQ5m4k+1Lxbj1Gghbph6hxOfSMG3MXjSKwOkoehT5hf+U5sDZJ7E
w1icJPyhocCMsDFsaYDVePIVuEZYU7QJsWqGHZwLXCUbUftHyRAwu+PsQKmv73l+XKoI2MzKg9+u
zk22o6lO3j1q95i5DUj97BjFDmRyEBcE3tmOuO/M2DRvcmABp8gxki/AnXdzWJ7wN5QWq4Ecg32Q
buNChwgU5QLBW5PRW97KoYOc38wnj0+rQLvwUAOj1sQY4AUHDnW0HFSkXFEhRe1XMwqU31nNl+J/
SaTaNKo/IUWAN3eTKcYCIMbIsTw2bsYhy2g/i9xk3Rm0kplmzYWa6Nlo54nRHm855f4PpYEzl1Ib
73/OetzWcERV4uBejI74xGXtDTJmvdemTsAAIG7UACZAWHWSTPfxYqLaR7mQnjJ/+lCGN7RmUZZi
D53PvC3tTUNTgRulImMBH5x2wabGvjeIk27Zb0nkfRBFPWXs4KqHgbAQSpW+RQ+mIZsFdH68Cwuq
PSSK8bqbuyp+qAJGBRNV1vS9N0hj/ROQ0DRKpO/PJBZbNcogPAD/rBTH8+rUM8OWtnlCQczHng8T
YqyyftJhgy67jPy1AubxhfvxgMQ2fwL7VVLaGjDAFn+ei9Jn00CjD2rcxXm54U2wMEeAsBXusFsb
dqQCoJlqVwQuIYkBnobodvvOYSZF88ItN+OsR2XtyojfihOCQDiZrJxxkbh+G5QKygeWZs+UkUJ9
xIHY4eOYJ+2Fri/7rIU/pzPsqrPIIXEqQim3iHTlLLesY6xT6ARrw5UGzEdlQ93SyGJiZ7hGbhWA
gmXaEVAfyfmUzAtcs9Fw25IWvGinTI0YlHNUUMOowYuTguqqwWVCk2x9n8Gbt577WilEgeBH1HRu
arPtrM/BPvoqHkCnchqbDTz+mhYA3xEWm9V/SBXsO/tV8bP/uWsithQ+L/sDLinE1lLEvcP0QZhP
kr6ALs/1cXbAh1zkkW76rG3aNoJmnG39SLNacRgkXYv50k7PVhtuPQPEzc0b9Dzo/t3NgMci6mbw
ojlPfpYDyJAZ45GhM8VwfMJMsMgAnrg+A3eot1gyuMFBN2FxN3CV5ZJsA8tp9G3IcUBowGUq9XVa
mHd8RG0aN1IWhtvxZTbBkHnBV28/CS22FpnHYK1LWYE+3j7JY9w58ZUf6wdh4RPi363rlVdubabZ
SATI4AENqzJol/e7glcMJ2GXmv1uU9wHaX65FJve2HP2soRIaIz2Siw8uiT8Iimm9FW+XGtUJpU0
nh9+t+xx8ChR94CCgZGgIn7iThDOBOaQsQC6v5NjkR6S3xUAiLubLBkCSlVt3VWYjCebffE/kbad
tqO4MbYG9cu48fghZskyagEf3HiLlxW2ZGqmGJ2xldzmF3cNXF4mUKE8A1k2+fDJbB/6XMrgQCXP
79rlqkimZy4m7q/CDZvgkLeESAL+LRzXWSSfHEFkCkCYJCbd4ERHqfADS+EdHRghSnXOic2qLVOj
P4Fecqo5PHxKXPxpHKdooLYXA38XfiJXkl2/laXKNEKpf7bTT1DpWFl8dolL6NIkiJc+fsNL2TvK
JuHw2nyHduyXh9fNyJMtpl+sNqI92g+wIitpB+2u3AYBZbNWxyDOldSLZX+rMQ52fv0X/x8c1S3K
1VsqXPXrEIaUFDm1nhzRpVohDe41nSHXc1G2DnAemFCqM4mrchi/RYuJnF0vKI2lePg/yw4Z8wR9
aSP2et+/dQkxw5raoyyPQasMWhuyHwvv0NZpfiOiLIIwukfBX8tUEeQ+ms9+VW6dP87w8W7qOf3Z
l6Dlx6Gljp9C8LisIGnwty/Rc9wj0JLPkgVSntDIs0fmLbSoksZrON6JJVcvYWKRMDjTNdWGbnis
WpTNrCeilQoUH08TXEi+lMOtDXMzGOw4znFQjlr6Lvpr0qsrt15mezNVKA6rU3xlGeC3XLRgvs5W
BNnB8SEuGPG20P0NW7s6QiOMzlAmmquMOlxxYfmrC68wqDC71MyBhHz9UBBE0zupIoyUSr5K/OyS
i9CuHQ3FQnPqxNTesqZvNeRMiFlgE6JP44JG4nkG6lbdRgVgYTHbt1CLy9/yWTqYsKcJJP3va8/t
rkXnHOZNfUksC5QgBC8BXV0sF5vRaDgEwSQaNT4aDrcr4W5kcJFhBAo2GTPNyst0Y4tL8Vy+iQD6
2fe6cwaTMn4zXuNfhADCjkaQ++B+F1iMjSfw28jr7yIBktDcD8noNAKUsvNUja3vx478j0bnndUT
G2+IxyoTm75OUQy4EMlccsuH0PI+QaZJxAsZrtHFNp/rgUd0Sp3lmcUQQTpMYZWlm8xl8dpGSNU2
S4SYJjP54ybWb/Gou2jtxO9SNmIEIBvHT1EkI4/PiyCrDW9n4UNFt0+VwejOWxZD4dBqQzqkdOdJ
MeKkD9OxfjMx7UcsL6BgOaWi61jIpfYxOCQTTWEGnH4T4WAudM4fxfY/pvepohvqKMelFxldZoLB
+JG09KlIQWpCxMYH9a72zv80dJdkNeDE0Ns+whwILKmxAEepiRqQfzefUxPiMBfKv/JdG11tLvZ+
I5txS8WfoetZnaVXgmgQvO9zsgvRfe2GcoJaiqsMr6H10ZQ1GnIR37z3ATMdCsMhsc0mIRdBKAvI
cIfgHRln/RGBkrGMsR2tQDCWctzBmj/aB+xcBshuuKrRFi28HDFIbxg87ls7/FcI3rhUH7nc41YC
CK8L4J5pM3ZqUhs7pIBtp2o01nY+WglntBdSc6xUd0lwDenTkl8Df+vVfQfodyHDmDXMEAt8A/vC
vbofW4FO+Y/HZiF/PfejcAuozlkqpPeenj9a4/P2Z89yKwAbjARoft+PSe0aEwgs8fb6P/FMqSsH
4W9AmrHYIqLwhCybheGpsNLQwUyow7qloRJI3XkX+UQFyIob1XuOxSWkoAG7TOX9DnWZ/rHr6KxY
DR6sS5F9FUySuFWriCu4p8qeaUTr2+bnQenkZs8/fkSUe3rnVDtuylxqkyyWMaHyivkxNn64T+Vp
KXYNiXz9OSHzumC77dqcn1s52MumY/E63kaGft9wcb43FF7rRu9XuhRdDyN/nU6j5V4C7ho5e7k4
OEYFULLTeg0fD84KRKXFW17dqBBvvMUtYW/p9iVYB8SKpLZlDdooVoxmQ+0ve5CVhlVfeg8OphsX
grsZVPOQYJNbAzUG9GeznjP/KsCywWS00DilUJKqoXSuIv3H+whqTg5aP6oRqgmlIocJxc8xiDUT
m8+hcc9FkDkLTh98iw3A2JBizDH4QMpylqm3JzzWxWDuS1LQF/JwXOXXq9nZTrVtWK2WNaHnMVsS
Zf1xWnMG69tSyUEmRFsNrzsepFD9akKjdXzxJxVJ+6CI5yeVpu2yj2yrlJU4uZE2IgEOurIfoEn4
TlJFSNMQrVHYVRU+jpJU7HmQOSnqvjh/GARJROFj/VFZ7HZLEakild2kZQQGLv4EUuNjnXBHLYpq
3rulVtSTfbmhqfC6ZVlGKVB3nlULj4ZvDw1RC+8uO/p5P99tsQgPtP0Yl3QDUzek7rVnFwbHUb/X
HbWw1cT3NJQ5TbzntdjeW3bWz0pc1ymaw+3Bdq4kppnB/nP8z4N+V3w37JV3vBHcgi8VZ5hkDBVO
FE2O5EoTejvUJLgyZ6QYKTiGqa5TCraiZPn7B7scD70bvzf9VyFzHcSLOA/msiUKXhTe1MoljFkr
fxvYZQnXK+DUw+wKiagxofDPzT4xBPCNgs/48PE5MyN3NvkV7eyhcQpjHAFDl0t0g6Z1SaIvNQiQ
3knWDU7ittdQ2Rc6Wul7/Hh82QmWz3BQgFMZx0HeFKG2NjLi9cYM+I9W5nmOxzrHwg35wF80DE10
sT8K6SlG8bHNEel+DyT5HCRsJvUvtVJGhFDzvNo5Gx2i23RIi3GwwXBPj5xs9bwV+TfuU1c1b0Sz
T/b1+wDDTUQ2eNEdVTRl4yFC1b77UOUHmnXAodzTSc+pCaWiXgq8Wecx3sg1pLrkrkPfbUzgOHB9
cjaYOILiWagKDhf0zSlPs5XR+oPCFVjOL0xinVX2hIy9dPbi+TSqlVBktynnOtjN4GwLA9CV9Qdp
91DLq/BMc6p3NU250KH8t9+z2HsTfz3pbeaznd9mCL9BccnWe8gCDuSaVVFY0TnG+0n0eePsDpjq
n3qZoQCebahr008kKHwmr+1+SPKzwrCphNWx06y5+fwtNnBCA2tAz1dKivIGJjuAtxAF3PaB99GM
b9tyN8FF61IZ6GDsw1+rYQBmyFY7FgdTKzWGu0qIqK1jJULt363hZh4CMtfWhobrCLVTiDPx0TtW
t4BmEdw6q/2kqeyQRQB7wfa78VQ7IHcLsQ4z0U4gH0MfADPPOlaP39CTVFlOhhMdshV93b20K+eC
vM0t4QXU/jS1GbcxbcvRlhyENG2IeFGN3ECYUNXR+hEM73dHhjkWLdzBGnT+zmzJi+dlQvyWXKYz
dwmecwKtzmKpIp2bTyINIf9VPTG8dcfNLhrU3h8UOuy8gg3bG+LkkQgTmHq3RYGgZnsAWaVs46wZ
uuU43KxeMiPeNldRpVPJ4UnEhiJlzamMynVAj+dAislTadql8vCGcC9cGcD/8WUltzriCK/XcTWz
UjOsF5V2dnXORJgU/nOSkJufokP+iRi/AvMC7hBhmiAPVihqW5tK/c+ij0+sSEWxfJ5Sy/XRt/P9
0w8be16AhlW3B+FEISOg9fkVdtLbZy5X6+dv/y6dvm/We9E9/UVfoE5QhPF2miKYrQfpLA61I0ke
ZNBwr0Edc/u8Wdud3yjurakxnfKbNVpg7QuIgwpPCV2Gqeg02eFFHgODIbQNAvMAjlHVqKN+7lu+
QNt/cyukRxXZLDmy4GP0Z/W1vNeYeXSja6ccsCj5FebvEBDIJnlgOSe7g/aQ12T6+rCobt7LruOe
5pWeJDEQz+OqvrBjag6PDEFmo9Rm7LRhJ4MsdTQhweEcmbJoYIQLRBVExNX4d1/0Wrk+CoxhGqWY
im3VEGX8NTAGrUu/eVYTlkunCuhBhEMv78rhadph7P8sVPcB1qW2XUyuIiCH0D0Zcfd59wY6Q7or
tOTmOO2WfqqBoocFXigX+abNtE4UuDR1WAnxizOgmrGJ2ksF9VTh+dLU0WTN1TsNVXIcZlcutrt9
XVrYH3MmZoNubQtfK6KUAcztAZ5xKYVNEJsYvwZW5eNCQkyx/ID16DQoiSlcveqdHl8OFiRdKG5x
sgJvKDwMOCrBxPsYuf7oevpSSw+mn9EnW7W2n4UE6DlNygMftpR+vKN5/pGVwum3TG4qS8ZZogxS
A90ES0mSVDCcNF0OMwSuPGNY/xtmFa6RHjC4ChsQFKjp+DhisVpPwRKNuSEaB6oCwTN/jOj81lOl
ZbtgxZiMVUeAB6bJKfeDiPh66o7YO3zr/iN+ssQqw5BEJbyCCDAiEl6vbghzNVI2jcaoGHaVxYon
rmTJUxLH6Zux7bKo7BFlIY0kvYbs86Q5WVkFutkIAZl0sYGzAiw2lM8DoAGe+8PwBeczJflHZXP6
6cPbuB/Ea1rWKrwIa2Xkl2PHCNQxeZ4eRHsWaTduRftE4sKY6eNiq9jZHhPsJyIyOterez/PWCQu
3QPu4mtSVZVbqYWyBDzrJFsEPYspr0HLg5+bgG23U15LotkqSWsZ/TV4K6tHyfMHC5xeu372t9sc
/z1JJQJfMSYoJeE29MCZ3vfsFAAlvsYtxzKfgXenhreKYKTibX05sMf6dtranDTG9qJ/gRKXXkM0
ibBe06YuS3FJe0fZ2dfuDcKT31twsuSODWrZ78qRXxScre/yCtmFTC3FkJ7O8eFSE1+Vwk/QZBXx
PhQYvkq10Z8kk1gXpRKWIv9OyI6ua9YlBKEq88dMtQn8i4spgS7n1ygkNmkpBBF9aHWH9ncLmDmP
ecgVZflbONXuSoY4XuITW1/qxBkEiT6EdrvEV4L0QEFpIwFxTUtxmplVRI7cl1cDpJzi1uRdVEeZ
/HEk3rcfYkQojZxOKO5ZuJdezG3YV4rfDF9+Sp1dcKLf2AJgrRELfMJeCArykipwVebkLOK9r9SX
UybOe+qWq5WLv8K2EHLuHAhG83YbfS6R9f3rar/bE8MWDjuaHAzK/FfNlxxFdu1Ph1Qp+cmcyMae
x9uxB3unys8EIvyhsZ272NOsaQhiZ0yYrmeCmN4J8WeHLdUpf3Gz+2zWiTFu3ahaEaZ07N+V6uJz
nOmQKTKwwlFiBxQ3jq0WzeqiW4iLW4890A1QeSHossoR4Hy7doMz9E2gmHvozF/V4wmVJ5cEpFdm
LaFAkv0UT27cq5JRI9G/FMDqS94DFrqzb7VtlW1eASDfeQLtFSrKUrOJMCz2ClEhV79g1lrPOXTI
kvNTot32ynIR5sDoYP7kGhQz/qa0uDtnH8/H0NMI9Gcc88kjacrs1iu7VWlTFPoqUUzjQmAxW5IX
vcdFc/9nzSvzJd2jNca2LRjS0zmLc/4KicOK9+O/4cEozY6cl5kf/g6N2MuZExfjlbBvJgKs4cBT
vUd2RQcFCZqx9p/rMAa5uVmqRQ0FFvHzQCHYAzPmyGLpwtM4CsdBzhxidYl9nb8zOP78jdageEpp
EZl65oMstz/BECfYZrAqAnWmdpfGumIsWsqxnjRdLT5NRjWSvL0w5QxAc7T1DhDTRYhQI7CI9+Lt
NKO4NRoo/7UKEdKqNehecTwew2c/ZWSwsIPTxDDJ+N6ynVTJ30mSnUT0uGkoOdF6flbB5E+DvDSN
rRIcsxHhGwBs9fIeUGoG+uAhojKaahy3tA7/3EhGlQK5Hu8B/7t6cMIE0/DMscT07l0Ae+djSoaf
2cf8Vl5vjqhFpXWkUCYiEL+zPzK8cGcCUC5/Y4KObLu+vgs/o/zuEnGcyMMq2LrutHrAA3Tof3H4
mLJq2FfFVVDk1OHBmApDldR2f/8R+ggMxWj/fjhJT3sPAJcppsS1DuGT6AniCKFDixDMBOmjzF8C
MWLeOHJBmhvuu1CFiJcj2E5egCtmtMzlO13FcnN9oQZOYnuxvjsfWNWItQ/6oggtTYRT7gh51rBN
BEItys/VETnWcXaYBfUbwuqeyB2aWflHJz/MuDjkHnl9FiN7H6Pe41Ch1Nlas8uKPtgISXjT+0FH
7h/Hu+vh+snja5FqrSnH52rv9aoiby1+W8EqThYInVmTrSC7UZcoZr8yBNurz17D3ihs+tFUXEjX
w/mGdIrzdkZF7xcD6gIIzuvKyZB4rcSGkBHjC7CCeRPsuaErBBNNVDA7DVLWmtzWVlcGUZnFuDza
prwr0UW7eex+8si8nOiLY//eELLJxd+U+1vjLA3kVOoJ9xWIxKhDvDASoK27RshCyGMIZ5Ih/hCx
iZSDDmoexJ7315gN7sOdbl7W4a4sEudUNNBZ531Rj7c0aGfpEi7a+Lr3jOyShpz/2Djf92b/u68Z
qHBXK14Npbd+9G/gNYDKlkz8UZhZLwwMrv9y7uxnn/bZEfRuV49U0zbPObSwCHTlWljOH5cxJXcf
nIN2cQy/K+lQeGiNTJJOtaqY6clLDZaHZuFVRtXuLAjX437xds/diBfed4oQvbdzD4ARDMGNUicS
rFn32d95oTvocnmxCrQN6Dx8+1AR7J1wyKGxkv2XefQSnAdT+mtVBiay//GoVQwKO4lAdyrnKexc
1AaJ50rqzlyb6eXLFE3jvU9osBaTxFe2ptomFXpHwu/9LnCis8UvTISrw0xFpRePKNeX1sSep8rG
FQ0OoaGo1AUhIdZV9WBfGVvR4UKJcFf3LTBMm/pVcuRMwkoMlzAKbbJ3z0Ou9FSpKTfZts/YgZ1q
tLBRk+5VD2/uc48FOPvmyxJ1MlaP3tF8DcNR2n9JRDqX82cw2LuE4ok7O9ySoQBcW1TDAKJM+MXc
zgEBV8nZNTnFFfZfOSL4LAIdb3KEfhIcZH8/VyLxor5ublv9ml1XAp97/VQw69n0V2Bjs0BqojGw
3vJ4LoDfjA2cMv9rtY/QpCgmetSMlSB4oDAGCJI9BRd0vmrjL0YDn6paNQs6FYEIM7dFiNg8tfc4
0a168xNRyvGX+1emBLD1bG44qD7epLfvwkE5qKYH/3LQdpQbYFDEWswojVILojQRFJxNhLATIr2F
o2gOUxVT0kA2LIfnlPnJcmwkz8qmD+JcZAXR5uRCj/nfuu1MaE5ykO4hEFey8BNW6v+96OJpu5/p
FhwbylKa9j8hcje5pssaReS96uyL8p3XyeARH80BdACeFDDq3YcWWWBUpLYlQf1bsSW6iTJJmU3v
IDtbJvfCS4w4Fbk+sK1JPQAKX5KGrnwcJ+JzFE0ZpxdRozww7CdBpDzt/Tafng07tlEh2+yWQkCy
6+zfgRugldI7tSyTf/GVJThjlpKESssvw8HS5BdUnqnDPYQHTczTbtgcwEQRhKsiSQVJWWYw0SQb
VKBCv1ahZGMDZf01OdjvLWXCiBDlzJMCHrmewphV2gU13Wu33fHHckpLmRmo8OM6P4lQ9WYYM478
A4bZKNf61HUOpuTpTY6GhKJtBO2xdfhu3d8MkKu6lyPB9h4aZWYGxeSdAo0zsiaXC4SqhbJ8aEBm
8ENzzOVZwA4Jh5s2lVtK0GhK2BxeUbuDND3dzZRQuS+la6Lt8x5UUpmkGCP/rr6PjBqjPSG00C5n
HlOxxFxI1J0H3zryaYwLuVCQEIiiRuD1TRCRK/53F/qE66ybwqG/FIj1Fl6ZbXWzxvovWVgHYGmS
YGXRR7eTyyDsaAmPp6PkuQML3pPn3W32LZfPvoF1+LLyIMJAAWbQFozE0rF6jlnSjQmMAJLQlCbR
6TpFg3yKoFjsr3sSroYWmEOWABdQw8FDI1quwxp+4yjcS8nDx00NzTEJyn+g2rOHoTV1zhuve8+c
6EzO83ymyBA7pNctFwOug8LJfZ9z6MopiOcjCwbFs8Tzo6uRec+sqVHpjkYHB3/0Ukm6p+nYTTX/
LyA80Bl1no4C6RqZALQxsqwf+RLZj697dGRTdnsSHDEvxkwrsiVvqTt0jElX2xljiN4xU9hAI9IC
b5bu+dI/OgEwK36mVD5FcGtXBPmcjVDS8HeHuAAEzNryLs8DoNU1gU/aBHWZ95yw1UffoRGcsjir
O2mTxCDT/NSkMcwAWPbCshQT22WhdTOt8bbtlXCsw9hwLQ92rsnbXprrdqk8XbTYcHcBw8wTYzm0
J6WGXBiJMmFPfjRsX98uCvn7Y2jxev9VVaXJC5H3s3J/+qrHWqJIBxou/KrRgQzoL4cK02CxDP3p
4Qr16UkVYpHa26M5juvA+BLT5Owu3zt1AqWw8eYp0RQsjaztnSIBcEx+c0EP6fEsJtjM4O5UsjTl
1TDaksxtBdwE6+rm2AvWl7RhXhTxxaKAvZfQ+6hSzJsH0mFKFZiqw72agKVeb/oi1iqXICYuiX3k
w+ry0X6ObRSuFl6SBNnwHJrA7crCRgKbRmCZFW/bNkrUqJ9+/1LFLFWYpeeQBdlLpE2HVn41IOtQ
SjrP1PweGc9R+3R+M5sYsxHn6JvW0dKh6empOQ6vDElQuWJ579cw6sIMxBnnPc6kHVMEBWP+V2si
ejDJCvdjbEBXNFcqHFxp6GnJzW61bw/iVMA4FH9FukluLX0hMrKgKFceDIkfzwFqYLvbwGpLXmcu
FDIf6Kb6EQDbfntD20lChWMujr33nlyXXW5d0LvAytFm5dIJbk9UYNYn0L4vHox0pqscn86zmOK8
tNAjo5aCwpsfnYW9woaK7PYtmfuu+X5LhPG8fxd3AGKQQMQSSd72P/h9eE6qL3qTPcVy+khUipGI
u1OMAlJmZDhN1eA6XTd0QRq5BG3WUoRNWeQyJvYMtwkoDmjuIcNUYioC/0ZZVf6qaUkEOa32iJhb
HIsWgEAyI+RQdDBuR3hvyljR0zHb0efezT17mZryoZK7Wn18zXaTUbTivNtExobwGfhq+rJQnnO3
09gmJ6732zdnB5BPu+v+Nsgn3zgKcs7TqQd2PF0fuutgO/yDhL/LYi2X6lhNgHIudUmrmRocm4hj
Z3Vqi1h3v0qP3VC6ymPqDJetlfr3TKd23S2gEcdHaTtZMiAqQxN54Roefjo/h/n153SsS26sc2TM
WpEcUipeQ7JOBH539jwZIFSom6v40FQiCzu7r51gjFm5uxW5s8DZLkD2mAAcDNWC1ZxXsVtJcNgu
M3J7aiBfiB15YbLqY6NTKhguTDsVSwmVGz5FvyxMWyj5b23bFgwlYOJmBArVfmi0z/Y/VQA2nGwa
iEre0GE7Jn60VuhUwlIB/ijW+eTJnira2fUpmt890vUE/6p87BRBW9b6lTLbO2Cm0aahfnp/vXHW
v85E//qzc3z2mQs7J838tnmJtYWcTwctoj5j5czF4zR8PYIv49UN43RtpFk6cOLXSzwUWiHsJAK4
B+ZQ7sfZbUUEn7mMf9Lr+9Y3GfNekdClfAqCCZR+mbsNzbtX8w4URTCdHZdKKgmmHnIBB0BjRy+2
KpmEE4HmuURDrqLhuHH+vY0F6Zy9Ut6bwBpOxYvZ4ZvXfpdtlTlhLR474ZGgpklGPJffzCAZ1VQJ
U4LJ2SFoc0LZpg6AehNYLPCu27z59zLQpy2ITHh6zSezWbPYvk71noG+snnK7M+jNqg1BQZtQvnX
UapEEb6Q8Vy5b0//kWIF6EChIbmqCJw0bQRPEX+gd0+Qmmu3NjD6Mv1fV0kiEZz0v9oo1igtc6d4
A9FK0PqbZMwSDe2LhEoVH4h20ifA7AtNJhBMTFV12YDc0JbNSr+f4c8T6zrtXZVBjfMIoIaj0A6I
46/RtbIqoSHPPCd1yrK8Y7wfRvXDgbFaJV5NaTcOvFXOFGM54Iw1QO8qQT2OKs2lx+972NfeqYCk
HGSUAoDd5zlkAZLCM3tl+jn/UP83N3XsYUuUXRt5EOIW7qe7+QyY0FBDBNsfzTXLczjnymyz2K86
kqpE60OGk1/IqfeuzzVTZuFG+pl65DPKOcOpbOEu8VKgvqC6Td1wfTyX5pqpt5NNbdDakJEx4vDV
DiEv6dBirGv7LwBBdzhrtdEb9uLKDVN29OzfXygXVnFJVdXDkK+4MmcF8CYgHlIUYc+87r3zutCf
E6PNZ2dvDvK18lHRv1XUCTBASLrnBm+c8P1aNYeX/BFhkGHFzSBV8Hzc+E6ZUX7qt2OVRSulxxTV
Jdi2uK1QuFNFznRQ7lN3GHkXq9Dk6ArjtGz34SclV/pkvyKtYLDSpLlrAtylvvMdRiaAjp79enuO
dWr3MLUwHfO336XJJKCjdkZ7cmCXgNn2AgRdAt42+TiGoPyhwh6HLmjnC7psSB8QUHQ45oFKERr+
KAGkDr/nIM+ETlNhRYNfN0inBgTpTrc5fLsydnJ0TetfbQRru2cLkXHE58kr0C0O8a9ujpsx6t6G
KFuYG+A9xCbD8tTYBRrI5KoBkNtC9eVPjyPUDz8RFnp/gZf3jCv0/66LiV5XkTtAF3tbzR+DlCIO
dy0hzge9wjzzHSDyxOf8+JoKNaNaUm/7u9+rXpwRgKTi6U4n6yBv6/P/tGCavYtpHt5Nezaz+oX4
XtJeN6527OxKg87DqhFoh9izw5MS5AbPL+QN1bE2p9B+I4RDJWFUACWL2XsBQmFZ6+rPY1O7hEie
fDW3wRL+os7legRvOKVAkW++UkOKqsNyJCKTy2zMO90ep6ypLkzVlae8MutZwk3g2xzTtw75kdnw
l8UxThDQxwZ9mab3eUi0SXk1al46l4qJWQ9wk/SttlUasFx26cmKNoopa8CCCTzovBF00TrQHJvA
4FuxFUBgFsb1dMt8tn+DD7hv5G4VVRzh2lJZHR5hFuB5BVu01rxXeEGwtFdq4/uiwg3ZZ8iG6/Dh
EDoX6IP9hG4Jt/RQ/yIGyJkhQulqqhSy9Stg7esIi8x5+FPzC9tPaHEudRDPUtpxHQvq+F73mToX
RdLjTRp3swk1d+aoZg7nKWFxJprBNNhwJM4wtWBffJwlH+wgkwNHdCZu8ncAMi25SqkFqpRD5z40
HnhWM46FHALXoZOX87uVVzFcefPFcRYPXK3mnkTxHol++xpmI7k3mvM6aRvU24YrI0oGJfP5Ej7X
juzLC0g7Kc3i9Yc4Xggc6iLi3Py584jX7Z1bAfJ8z5qm9tmJiK9bTPgNQ87CG0WRsQcIFnwoCFzE
v50xCEhE5CGcz7/5mgLXuBSW9D9Eyqr3Slvv08NH3lknt4LxXMij/qu2zi0ymF54ikBTjbPXHOQz
iEs5YeHVGx4jjSYQZb1l3GXM1oZkzQ427suGAwPCjG3/FWWoeXP1eX3+98d6dGm4SWoS1IKK0s+q
shhrQpFUfEMC4qN6+F0xA/UueHYuCQyusRDTPskVg1fIkehwo+zx7OP87gRCaVXLzzaiYX8u0CBI
lZuGMwmg9D1FYPQ80RqxKDTuF2ZYE8/Grz+ruuA9eqe436g1htOTRrBx+cX/InyFIUM0NNjiDXOk
DzmWmwQKdkoCioH8xoqmJ3LZ5wi74tUoL4/u2C6nEqXB2aUjnmjYQbkb6b4Su0Fv1YCVrIp+kJNS
/OhSwKZZiKB0BhBlxt/zRR0rJ5UGduMGYsGTRy9rhKohuTIruCS6h+kY1HaO2QT+ZApPAHFmLzgk
/UpUVq9/ZhiR8SbbzNAr6KgJ0mW06zyp2CCBrlGC1vudNTt/4IGd3+z5fMbLUw9HL1+hfvhgvrVI
HFLhajLocHIQ95f1D5M+OjK/IsRozaNv5SkUJzHjsy9K8xKWaG3YlBazCyRyrRHcgOY4kJVsM2W1
9Dm3WJSn/0ueKjqmoNQ97ZVXmVkSyALGS6bVQ4w5ql/StFWQYxlKagNbR/7tu/JzWMw9CqgljoCf
exZAVOEnhYLc6VK6V+ZpD/hVR0qE78i+2sn3GvHXdPUnDUbByWVVgtWrB7uAzUx9Hocl97OSNZ5g
5IVKFcrT02hMr2rRJwSK7V0F7CgWKj7fV0SeItm5omnL5D9CjaHmsJJSJfrU1fgX0uiqaICm01O7
vT/vqwoFgen2e2Deu9A8EDJOtFrdGcb+VCtiM+plZ3dzR3SdsTCXGaBHH663S/Ctniv/sbBY3oWN
gx9QalVAOj4gYRqnmvIxV3Djn1Dndr1vse5ct2xZWvyo08/uhmxboSanqXRb+7b2AKlHWEl5N9Rz
tXQVEvUHkERLF5uqR7QY9AwOAVBRVe8hbxgqJCAHrXZO3b3S2V0s4RJn3rQBakF7TbNPpqMPjOhg
kHFBtGFQfgofdDSKNy6jWh9YF8g8uQ21QLdl0I83ZSNpP9KeTYocFJ4Jydckn1uacV4eauwYW+JD
T9fltkuw9X/5cT2n2g0+ug9N84bu8zMsmI3nrRBZ3MHJcLsYiTFHkC7YUaPkMZyPqgHu0soXcoYG
QgXMWJF8lwgTPtcbXLooB37Tfg3pK2cnOxtocPdFP0AjzRd9CZwEoESbvHCRXv/dJ7VMzBwf9WLA
10bUCd3kh6Fdad9iK39QgqllrLzsxkI/EMLjOgIBJ0/qLH4Fwr49ZnvR0HzNLUzAo2BbAjhCQtWr
Uf6DPYbaF4zrPL9E8FfyTshd2tLycyGslNzCb7e6sOM/Y9F2OnqlzMvhvCm06eFE9ZcvUxF/uXMo
snedf1/Qbx/UeAYJG+ZWpgBbrtzNzUquJ03tm0gbpKuHndLNv4vAQbj2V1yFNH1efc23ibiqTUMz
xOtd0mElitBLbXCW3qgacUtL43UssVVP3nXDigbp178GKiiBopuhKqfrJ5DrSUOOAXGfl7L86uOF
ct7zgIA7BQ5lyt/OFGSNl1W+oCCQGHbtqyLPdakVTWtEVjiXPxl1JGaZI3uoLNjytk0qGO78YYdR
K4/xVM9AlJGLL/HHZAZH/8NR9MppQG5ros30z3WwflCloQesSFV/9nbgpEUcWIChswei6jTgoPW3
+Dc/bIipEx89TcSIeXuKjeuVESVfGvLGXxRb5Nq+vEC+R4F2vAMnFfmDOtUJa537/K24CFxnI8iu
e5YsUQcM2m6uR8v3C5h4XBOpbLnLP77zTrXt68+rq5vam+xAMKctsVB3biTGKwOs2F7Vj6KWqvRD
fvgkCoUOWVe+WN4viYlGVNGBdaUmcJQ6dh9gkmaHFSr6CLDCZ0bO7hu9dB3D3dR5JTlnYFALO3GH
MPg9KyUGtNGV/MTHNHFHYQhCXfsensIw2JBwOUH0FnWXFem6b7SlckicIxHJWgJPysysDTZDtuQG
C8jAKOSpripQOloOPkiocwUCCVlJyzQWtx0GU6/4zwvzfOQ2GRf4kEyisNdjuH8Mg/kZXWYnnrRn
B8U/yJhnRGNy20nvxeL7GrKKpfPluJN7tQHTXuNwsqSiLf6PNf49UIeEYiumF6k3djXMqEwaawVl
yaek2Le/Jd1DlwBIlXDb9GoHvO5ySqyVOh6S5pz0jFVc+4zyqLzGgawvot+8A1RxQVcoFtudfXmV
eXcZYmXcBqqkeey6prl7qGnFESRrovOR+JRjYfnMoOaKJQdpHne3OFaBzmjUDLZQRpNXmviFM1tE
RF3QXeUztXdx6YUWrx3dggX1F7xedVcG8IAf5tL5Drhbe2eqbXDPPibZuziw4kyAoITC5IJUqa+l
vq6u91AF4VcK6AOrPB/k1wx/h56OQos2KiZ+8IC9P6owlRR/8JIUurd63Omtsd4I01xgoL5UqGfn
M+c+9uV48eEOplfeSFuwUUWghp0NLo7Y5lxZEIPsBBWOMEByWbtVkDZC/hVAKPuoiPaXdsOjZ6G5
inYpVttXjJ55/5yr0PCkXwtGS3/qHUCC63zAIbAgqrUGgNYmYbGjG5T2kDneKuSRtB54CQJq1z6L
xNoMLvcgt+BJXjb6sBtK7Y71tQwXjRH8x+4UgIiGSDT4Cqtacsn/8X1LYMS74pRG+2wsR5Ynzndh
JZDOfATLN9GLRs64/WxPgI6KWaMvTC3O0zLIhOw9EgLcNywKQBg1Ib2PI6PHeOXlBomCQ1F5v/jR
IafgErHx+n0ZAg0Ymo7J71qPbicmX9JZxJHAKohEyQmjTK/5LQl1JWrNuW8ntGVBRqnQsHQmExts
O+YRpdQBV+aIk0twZhk9TOaKH2aHI5kTKY5uT8oNs50VJb4xEQpS/DarFGXLIeIT3AK+Mq8vMTJ/
p4JytWBeuZgOHy9DFKelsXOjq1uxtMraaEmU4xDa0LhpKv070Md4HC+owkfkrppAknY7zw04JE+E
mL3XwfIyMc4wNeVzaCBvsEI8H4/dO0PThB11Oo9mNQnxU/4yosWV4UDO+unzB8NOk864ruMuADET
Eqr5fXA/CrLBxiF16hrG4n6oHpz/WgAjrhfN4BlgD+/MPZGY57X86PBfRuA+N6xAMYsoC/Ea8eNa
JufNk9RyP5Vr8d0GYsMZJqDPnCo6kaOsKJD2ca+NqGRUWs6CooB7/CPf6C7oi3ILJsJcbZ3fK/sC
yMT8Bhktc07uSNkYt1ZJoHYjG9YTrBoQlYcBgIM+oicjqit8YTOH/tEwbTFEdpZQIM6zl5+7pnZn
Fpc9lYlEeDXSOGgQdT5y2/odPZtM8+LDd0HyaXBqHQ9YyaZTZhSlbxoZ6Jr6CprYH9Ze8yoaGKEn
cdwMiQ+XUS1PElNkusmEXvPphAs36udAT1mD9Zmd1eqh4Q0Ip37vePaxNiW+1titTEjXj9x//sCM
DSoLgGupfT/6D+wQm3TJgnFSytugKp4n3qb350HlYaAlzKJfAOJOh4praVuYO6wd6493gEgUzaBA
nIpBliiH+WZ2rIAsl0rLapbuCNBg8H9687NKLfbvj1wEjZSS3wWUSk/8S+aiQ46SNnl6HLaaHPvj
bnTzEo9WMlr04WT25KxtrkKfrzsNx20SLJH9QfvwgxMpixkuYLDm9q2A6CVmr62kFVX/wB7KcfpQ
IoV6fv5ZRznLNfQCjAXYN9gd8dHqWfNU9xRKquMnb6Ca5B+PwO+Fbj3abTzi8hmv2JcLcAvk+mhx
XR8/NTtGmPVOjsnO8YwVrpGgF2MwumA0yslYYPHjKqCj2tLgwrvQ/cMyNYUmZuYmWQ+ykVLLjY6z
9zCvn73uAXQSV9HcJ1m7L/PBh0AjBgQi/wXv+UEkshUtAqtBFlko1WKQnyEz8UxZl08AlbWW6Qud
xSAPTmlVX5MXbNtM7thdFsT7dr/NHJcS50bpz+C+vSUHsEgUMfeVh6NcrR5GM/UunJipAvQnyqF2
M1gYEGhSrKeR9D+uYCgbeJgo/3BIBn9cnvaVBeWl0f5c3sv0cjZ1fNNarg4RZnC3gUfUSa3iJcsn
8QqyMmmgolfdX7o5RCLEofj7ueFsV0sUo2n3+uriHWUyu6T7YxzzUC/jkIm5c6bNhsd9+Cabbk4f
k/qeoMhfuMJVVOrP+oxYrf9YctsdEfMhnhLfNkBE/Y7iwgtNsmrokeR3ir2YPWVL+2hF/GQnz7OU
Rekb59/0jGqgQibLPvRFVbHMZR81MHntgHQfp4oe+5yL/j55zNO6HGcfiNCKuDZQBfeukebnl50c
U7cEm2eeWwn+5y0I0yeZOFIkJp7TlhDRB0y7YuP2JYLznv9eftC5j+8WCeDg/5DX7Y6PqiKIRgYR
e1UNMQubk8/fOscjsp42zgr6J4TUDBmLnLNLnWCP8pUQbxRTaoTtz5oXLv5w0IMuwAWPVOL89QTw
zdgkMHZwV1TjOqdDFVNN94UiYF1/gEiAbcEbwEiBRB8eyZNNH0aGBGlmw9cmIad6PfxNBva0EtMz
h+xuUqYBFXNRXqaHW/Gox9LU8pBN7FkJjEqd2dKq6BQjTpwx94VDhPMrCJzbo94P+G5ikeJdZ+Ux
sJjGxtTgHTp4feswWXP+2QnPgZBqPlYipoP4TAymWE1/qNzYGOpJHMkxeAwGjHV4OYUG0AuK0zOJ
wvfuzaxClYRZDqf3bnKhUA+fNnkmp3PH4DTROLEcPtto+yLYVyWfrTC7Dz9I3cKWxsJER/jrZRoX
lqP/wy+tl2AHkCYsnjzt2FT7el9DOFoeqdj/sgl6GMMlaJOWqpnEtWJvxvr3SYoRP/YRngc8+50Z
JG+ibIjg8dr2y5/SR3nR3XcXIfEzA5bkqNZoVb65yGXPCBumQcSR7uzzv9La06IBP1zTQFkAgG2/
ktlYU0A1XovefTIbYMsmi5ss6CtTJ4ECmHXDHMt2l6Vh4U9K2E8I7F8MAT+M99+pe5+jziSib4Bv
MHLueUGNqf7KV6KW5TajiQM2nzYghqouQQkQ+/wEyXcvQEJdDmwAo68XZyLx04nHYayvGG8lNY72
gpVBPCMghB1K9b1DNp2cLJGkk+Ry0Pz3M03D235pF6iUWTqH48YUDa4fR8ir20/8HOVazZgc+XO7
T0ZAimWst/tV/UmU+VwAYE/mJvqEEPJTPBLbBroxhGsYVwV3FF1B8/2nEEjJRFJ91j5A9Syjb8+Y
kUcHdZU33DldWNHlSGyiwTrBD7q1JLKgEn3M5HHaMM5Vt288+7x0Rasy1v3emKnc+YRFnDW93YBC
MgwDqfPmgEgF6is0mY94A0VMfoJ0MNdokv7lX3ny4Zw15+sAHuTzsXJJy+PLL9LCGKRec2IdlmfO
NXbuhnbop0xPXA+9+fFg1nM1AXrf3Qp6DYcXRC7jdYNgY+fajd4FsQwb1aGJSE+Zc73/e67ubyam
MpFAuT0uT35vjnmAu3QJpOaHRbeCLwn9w9G4otRE7AWKaJ3ijL+AXTadFOSgiwIc1hOzNavVi1Cx
lJSVHqQmFjmFog6mqe7rOb34PmspyW7MNTe7q2UxcPcI8dZ6mBe1STrtEWqasZfTcTF2RHXbPhDU
4o7xpzMpQi6FAy4z+3HNGiD/3uiFBa6eRXF9XeavTERZDT30hJL9BnOthCVKx1+mcWmmFUti+r0o
yU6q9jZJUBnHqmtsD94DhLrPoMogzWqEIuSSE4snpHMwbhmtrZx3Ztd0V2bwOM78eg5SXx9AuKW2
x9u0M3gz7VPj3UrMe8R6NG6P0nTksHbO4RWsNE01N0SJiY1HotEM9yO8Q11cEatPdUjfOrT6vA5T
w/VVBBej3fq7heSvcyVrXVU2HLGBWYpuoVBh18z7eJCFsfww/IFapM06pJKdLpa9CJowaamavgJN
hX+W5vgYDnhBd3LeX7McXzOHGecGUFOAKEABdhHGS2DQ/7utYyKK4WoDzlUY4UsL3uyEer5lKjZe
wsjM12LrFSAb9nCkxnQ1hdAAfuC2l+8thxIY98WKNopotm5wJLy8RCzhTT9Uj5NB06bAwli6+t35
ods1voxPwxly8nhu7Htr7DUUDPdscQG3Xek63McQ8ZYd7oLOvqKd/rWzrNxaZH/O4LDhD6LfYEcH
n9wOIdKD4FRF7lVgvZe9N2yfbpurccLMcwCzIiEWGtQSrhzKIONIu7oHnvEpyy44MvNZpV8m99Nv
yCKiZ8vG+Z7huggOYAapEqzlDLPjBj/NfdVhMZZVWl1Qt0cp//e2n6Xr1dncJ977+jEe1jP55AIP
mUf1TYKi1hIZr1OlXUTX77qw7AvUel4UPYdxk0ApHrcIOYOHDSjGjkiC3R45XNG2N2X3pB7HTRhi
EnpMvAlDGtt54iQ2Ge1X6qd7Af5o58YUFFJQQRcJYrCtH7keQEdlznalMAVPeU2JwLUbxQ52oHgN
ySL5z591BZgIewXXAB0AqhfdiS4m5WhByEk7bTUAurADke5NnBhYboRYUEJLmY1j6dqZGmybgqT2
/pFMeqzE3KcTpjuXwJvGLE2dngaMZ/zgWmGlzAlidklyvr5OEhgADUJ05RH7zO1S1+Wd6f4VyXXx
F2hb1m+JM0CnMYs9AhX0fEh5f4QNgFoGOqnjidxTs/JAoisWfceBDFZqVoOIAPjiD4O/x52cOGBC
+I6whYOLQNL0UWNIBRahJJ/mYw5ffErdOaPrl/QZZ16W9tNQ5JJe/w+EbJcq6uh/LYdsLkHrvgBP
YJI0BB3YdNyc9uOx0v1miBD86JbfLLmghIcVgCKowlVxp8uEc9LpUdxrpdDrzqS81PyOvui3xWs6
0jXfY/U+r//fTs2+PkqTGnXy9TWhPQo2HYdJ5u12/OiHbfiu9UefmWR3sfBsnn7s6d8/tDqToWEp
lCgwlxQfMoU66MkQFvlPXj1jGCDR5MRYye1x6ZOAN/BVExlvjCV6W1jkXJYLjcve8s5C0XIDr4w7
GuBDx/BYEmnuUwNYfJ5reRoLgb/apVnSkYLEk6eqzDRPI+Xp2gcEylUSqjjZqS4u1lDaLw1abLmK
vjU2+YiHaxuiB5Xs1ucyp9Re0EnDaApLKDvvJt4HJ5MhnP8rQheboCShGFLfGgDL+19sx6AKX6BK
WAt9RsJODjjbF68ybC7wHLN91Ov2is96uoMc3KfCExrQiQiR5pMlEHRo4vW50jllfPoai8RcauBH
hQL84pA7it0IJpgivBMaAaFzAgKfKdr6amgCmqkDpOIsCHJuQSZUNHBIBjFHpSPjYgRq+o55iBDB
AUU5peJVUjTWil0cnf43Q0/5jnVBWhD6Yb5kqLhxQCNQp25vjO1mwK/e4tvK4EuZ3/r3H3k2Dckm
LoMZl/SJjgT+3rFCfszP0VIf6KmoyfrwW0AGGYJsWe8N8oC1zkhYSJxW9eiacti/bmjO/YxXdOFe
yFDA7dPcQwAvrEr5IwwXRy0S2P0VU5iU1T3m1BVIePKTBl/a21TifKm7iaeYf1RdXnKrEUlXu06N
7alJB7HUdcg6UVnJCC+Wi0HlEm0on5x4+EIB0mZvaAhsdnemA0tsPY/01r4qrjZk29aGyEqmZs/C
Xpbt1mJDVLr4FbfxNf+tx9FF67Z6J+FEvDAZ7OQjiIEEIymv0fzboeHNvlyB0Z+0No1qMt/lf3GU
6GiwdEeWvzSHL7pVdY/dhzwQ3YhSmY6+XttZeN/HNhW5A1aRTJ5II5fnRWrThzH1BryKP4j1AxAc
S8O6j6e4pt7PHe7TBiZbrWAC8SScIs7ViEDX1ZjPLlScS8+Z59Ahqon+YxXwDxH4dMlTSIJT5Hl+
c2ad88KysKoDvN18HtBhEOlJUWvl+VKpGHCgfe4YZqvzpoe7zE/5+l24HHhAJtx/Gb9HW6DqwJpU
TYa5I0KSRG8S94N5kHmFcnDwKS3pOjlFVd3RgZ+NJaCBjS3Z8EES9RCCWxAyVZLG30ngYnKxBV18
aMQkZvt85vHNZv6LoX4GpvHM4lTEj0ho4Gk8AsgJgzvtsa2nU8IVGnOX93uDjyo4LuIlm3YQc0eT
HJj8F6LpSD+cbiv4dFDCUwcL9dDclS96n2UBi9W4VH8Qco3Ocj1XRD2Ow/+LHyUCO7GIMDH/5jzf
JqeXQukEmgf0bi7dmFrTYugFxJCbcHZjwt1HTtrMdQV7vG5YBuuFO/2+pIxVpkz5a+w5++n/xezp
TiW20SbO9aZG9XpFucQjc1nTUWLw0jy9ee4/ZTmWFrTyF71X65+SnCtsmrFdLDzEEJBhPrkZT20l
RSy2VlxCiDmPrJKdRdPAUSiLybQdndHVBQnvd0hpyJuQrXkKCgFk7SU+utzqrzZqlBNjhq5ogN4E
zQAc2exo+X88/dRMLdcd1Vj8+i2Ychq89TjwzVzv0fxVZNroiX0QSNm52jUvb5EVfU2mFf9tgirS
2D090q37Vp+dauFw/1+8GkeW89Yqe8uUKrzZK0EO8veplGWLIeL729qFufY+9w9uxlMAyk1sB5NG
63vItYTthG/R4rdi09QGcinv2/SJx3wx21yOOvNlqksj3mo1QEpLow+8osqe3GHJodbRIOTVzvx0
tblXzmoRTwFj3y25agPAtLG/KeX3RIRKBGErtO3zgTXi6Wl437QRWeg9dhSAQdAJR/ci0njWq7gv
0oOM/b9aUUZbrVq/zCyZ5ltgDrZp9gjHXOiFF1TFJ2FMv0PvoWzA2F+Q/bL7tPDCEMKiavZDNk9v
uDgZi6Bbv+dv1AVlpHy8CReur4ngtqBYNfa8f6l2Hc1aKaun7y4HS1fDSw61A0L86z07xj31QiwS
IVZwBrTa63uSBC2runUhKKUDMnLC504DA4FvUYiJuC+3yUMmeu55sUWajg549cZxWnv5k3Pabjnu
jfd3MSEW5boGE+bsxj2DZLld3UL2nZQhqMm5aAvh9JZ0xCjoWjpo+XXtfXP0ZHH+hgggJ5HT0pNs
Uheh6/pdR7jVmio9jCSx+9BM0VhHCt/WxjRPhkv+GDscvxfrHcZ/AhuUA1hBhwd9h1eMlg7fWpuc
Cewl8+eb/08dNzqEqKESTzjFRrmjDnX761GhrwYcn6ykmOJJJyqap1qv3bryLpg6So3jtyUvMAcd
uYFd6R7fxHxGd88ZyWj0zr3JAluU/SJRZxHYsoS7a1wjjShRTl+kWTRopAhPk6y73HGQcRBinZ4l
7x+9LUc08WDjTgdOtTT92nvPSHq1W4vzW5TFZ/i5F0kZCBn/1dB5lWelL/TVr76Uc9HkB3YhWF5G
I++rNq1Ls+iRgrv48EUTbthPYfmj598kJqGb2zetWQ/O1LI8HORRUfjhMCO0sdgm9fQ/H3mAUD/k
EsCAkls/61bPkkw0FJJII5Rx6ZD51n5jUwHOtxRmO5Ds7EzaDRPvROcnvfBFznpMDXCMqPVF1Q8N
7kz1tPgAYZgWQ9wTNUN4dZ9T0c9EMdToxkrhFIy970D2e29nOV2/iXv06aeuRlPtH8FxDdGwNhYA
cZoB0AVKxXWPb8gIeTt2vDlqKbDSbqCIlxxsSEC0g8JHwgz58nvl5Nt5UhzePDe0IXYaLQGIwlsP
8vHjmWnRh452GzcQXhcpgw+gGT255SzKNxElP/7JHl66LiMUdnYrbT3Dqf8xr896vJ+kNQakSegD
VFeu9h0CjtuRk7OxATurLV0ULW8fgwN+pEJvjqyGoS1zcyPZLCSmN75IZmLjFo6KeeolqAkS1mX8
YvMlIgKcHFvV7rKy0f1316nL8fq0CGBUgPSSW+PDoCHgEZVx//v7teptuUOhcxa0+e3jM+To5gdS
/gD0aV12tC0yN3ipTJ+ih96SWbtntEy0p+DkPxSFI7btN6IzvNoyocDMVTQZXCJ6VfMUSnMWYV7U
M8zxPZ9ffRLacxx32+gCfHi7Tn/J0HefnVyOdzCwuAxbHr8OKlIVKKrUp1IXgbZObpsHDCzPfuo9
736aYHMK+/d1vK0NDoiJ1JWACqUADsRBNPsIbr1mffUrWJx9SxaiBVyHaC0XP+zQisFE1IKwXc1g
zYyTS+cq0ptG+tFrIQK/14CCffeC/Qyhx8nevMhVoUX839MZRyFnhRE1IXppjy30Xr7QWJvROAnR
52Frz8Dk17nYW3OXIs1ouA7R49uZxt8cZv/jwyzcTZ28e08JEJKtlh3bty/ggGz8OMp7bBG+puIX
4nZZvGKjfPC+1e1qZ44EdRGdRu8Mvf94GnuFhGdhSOLMTr+iIc6pMvoK7nSZ53G26J6ZEe+uMzEs
mtke4qQyyJ/iLy7hpILnm5//O+rWeMzqyNG8qTDmz9x2v6zP/RsTjv/Cm9mD+P7OHkeLdtc0gJlS
T8lWnkaVYoczdNtY2bm3ZsMl2Y0XvnyRrdY1I4o2DudbS7RckzqzDozKu/azbLC0Dgwvzx2KfH8E
C2z280gGXsHKFJnHnNnKQl2jAPqVVH0UxdFyunIyr8x8r+ZTMudwfuDqQnFDiRwLXL0k0eg0h1yN
KfMr/YQEs3F6/8CAaAE/UwvGiRM0+0V5v0HhqgXZt+g+hgi2ax3e8+2AljmMPECe+5abImB3A6Ik
DiEFzERLBeb2dQJF9dQmRAWspmAhHMng1EjZz/fEvB1KtrKxl3doynoI7vTC7vIB/paDFsY9/Ow7
Xn12am9cRGetrdbMEgXcTMB0rnAZx3McTbWk39f4zssClAz77GwK9/QDFxyZpJIkXu3yK3pCzWm5
bVljtpbpwcUMNMe8Xrne1yO2lO4Ok9NACgOkU4eUGgxJcQvd714TMRDFSWpJDTj81ezUGF20BspF
8DOfv2aY9KXUktur/DSV2al7CiNUJosdnQULfurBD5sSofkwwKE3VYFFbon1mOmupsghzp6cV+L0
YSKczlhlzN5ChcACu3fuRCfwqaU5le0h0Oo4jfpPXhtaddBz579BfzNDvqFs2TlNaIKhO0ch+LPX
3eVcBnCLoOdWOUT0QzA4AAzqXfggkCUyKp9d7bAaxuDp71vG94f/drBA2YD2x4CDnHcyVvxsLKSy
qn+IABFudERgO9+iBDGuBhLXP19lKjN8pg2e9swH1RU81PeRMu1D5Ge4Trg0ZlyERZlAjVBT7fX2
hAxcdoDQ0C1F1kiTo+vGfjALEl+HJ/ob1+HtAfjr8C+lqvWm5KtwcBQSkVdVOMJx5TeWuVaI9Whc
4qKr4ipbOokFXrPFL2MdQcGNlSh0tLNUiUfiOn50sRoyiCt1ovSh/VL0mdpqPmAsK3ise3UFRgXF
QzTun11eGiz+9hxE3L+OND7m1deLbav7eTDPyzumsOhxU3DhgkBYykZIqr4bndWxWhBIiTdmQQDP
IrZkJ95wwvHAEDWkdZNFA/pKZQYe2OxLz6wmTZQLz4uE7CHZ//qnhPnD8S0YayRrh4HJ6+UV+nFJ
suvw+VvuVOCUE2mnA/nl2F9Hr/Tsv8cioLKpHxDyja78UAu/MwjQbEkbfG4uSRKObOomb2Wp4qwz
8MWOC14LCRBdDHugXi15Nwb2GdxoWJO9OSLoaErMW9Ga/WV3Tz5rf5Id2vc6FmLP0ieWf0kyf4lT
PAS/bwllzYbrWQ44u8yKBThL7emMd/ZHp07fO9pxhSh2VkfQN4S/nqnxoTNLLwbv5galNmztoTEQ
VTg3cyYQGDE9EaNSEIFq2E0UJvetEwSWn89KSYWhWlAVb5WA8MQa1BaKkTVU7iuc1qnP2gl4FgdU
xsS2kUyuHcIrv0cJgXJgF2xWCahbcRG1MxaWHEw4jHwpYz7sNbpVxfUhQC+Yqeu4ijBGxpgwLTOd
nZSsIXLA6Jy1w5ybBTqLkypZ3x7cy29b4nCzcU71gpRwVmGzgVcfy5X6PZv8lu2vrHfXtySAK82n
nWnxfBnDOWjRWDgrnauq9NiduxCyB8u8jkItCFoo47DQkLFVNjkiOLGFpgSKa4KDnR8LRe/IofvQ
7BA/283XnsTl8DzCifUZzFclbGiIi5AxTf5o8ToxrqQ6I5wYDeOUqjLvqZq7bVp2dca6VD9QN8wK
IOXFDpNzUxhZyQt0f3XrhVdmjlglrq5xTN0xg2wj/PLTKuzWqXZApXaA6VNHRK5sZutkc685FUbr
B7BzbX5lykKKFMnw0QmB9E7hD3lUIaJTekfNZESTiAxGOpWX4UKGEL3MYfg7YzlEFwzruVUR3rEF
eYLqmemVkPEwRowS45We53pPxbbFCkyrW9xVpp/tdfXRnXhXfLZlba9ZpSCUrS4CkDcdQLANcRg2
n7sVlaR8BmNvhzp8/eA8kzVzZXOwqvH105M0TFt1YdM5PuFVy+sB9TWddjEvBvsNxb1XcPxA1GJ4
Ao1bySVyrQlgy94ClaT3u1aL5C9a/FkqSSWNJcNYTe44zZfHDsDFSQrFyeJe1E4JD/3DspCvBR+E
qH2rR9T4UJcEmFAe6AomyRBEBeNXEWf/vVIlnx92qLzDhg3eS0LyYpDKuV/CqH/cD4L/diZ/p7/s
49BkfzdAEYAMxZCAaTZDlb7Q2ryxCrHUK15q/vD5HCiyhlBsUTMPSTWGXygU1KDYnhXiNNlDcPfm
FWNvvV7bHruIB7AcZmbezssl5Q05DPMVgE+d3kFpDDAFXJxfpDG2UEcjOsooEBqeFGMuwVDJg25q
Y31h3ugSKwugCx8Ymz1sLG9jQCnNhIpE5WQcgau7f8vEpeu/+wlE7sun01fqor/QjIB2/6+aEsH9
nnVuAaHp4bM2AP7YdiD28pHNI+qQqVFS2uMcA0N7zfQoJoH45BQTGj6Oia73Ymv+xQFB0uoV1KMs
34HcoAbIDPdBV6dqxZBDhyktDuMINSU0S5Z1FYiL6k7E4roHmUAZ7HqIOZO+Fmn+QHg8Mn+CVqo3
cof2zFoajP7GUGNBXl7Go+VjUJFbJaYFChjFccw7WJcwzHv+YAJP4YS4fBhu274DnYe+GuEGELkF
QsWJDR+Zv+91xE1pVpYdde29Uif3EWRbxbyaDTgz0uuxM/u5hPY5CaivS4nVpiMMcqgUtQhjQl/p
QtXQpi88i4s0qhPdCLJutlbRDZA/GIpwPEw76x2qwCoGqTSOEonkeOYkyveS88X85y+cVi496feF
nM8ZR4I5DA9vCo/B0W55Mejrog31LQmbDEzSvgPXfg0j8SYWgPe7u5Jdg3EOdsYEV83u5htI0NGQ
tMRDmW75omnrPVW/ZWpMCdTq7pvLDWipGEo+uueUtJZ5nqlsAoH+zeLiw019DN5w5N+ODxr3sD4m
VdyG/Owc1xcSZiwx2kHMLI+V2YXRd5uoLnfY1u/mCZJDZBRfGAN6msae/UyCH3l22ZMImbAjy9o0
sXid+e9kOm5HDEhKnRCwD5KwHE5veGVWQwe0+cV4l0PC/kLYrrCy1bNqsWPuLqnIYUhD4jiyHFAO
FYSc3iFcR5+XXydRfNasLzih0rOUHNjJXSKtwhv0FL9VaPtbTeD8PuI4CR0ftZp2b5+oTEHQJuet
0vQ0WeDjOTJlgDiotuH0CPtpJq1Bsa25+OxaAqOLAj7qgTuJ+mMG9xglgu6polrAYUWXVGjD027u
ORcpVwj3za2iFSSyIfZfUNMkSrcJP3ZlyISOnU2qBvdqUSLnxphVyBRI04LHSSjgg6w+t75lHjto
ChivNQLyGi3/mNZpA24G2PVkabSL+gbEXPKpS7PPSapI2ZZIW2kTPZ0N8h57Jhjiwi+7eMU0n+Ko
IPM2/T0q+9ngKYlGT7mmyJ6R5erIfgJPTZAFHpC/7zPwavG1kqdVCPECHWxuPxEqqxXkhNoPeD6D
hozs9cLXQSOPqmLaIEccYdVM2kQaeFr/4nOqvWaYFL6k/mX2duNWkcqp1szNPU/Qadjv0hPxiIUR
fM/pKf9Do9ePwiDaafAfSKaFLIouFe/kwXf18Hc80A16Py00i/ybLRc5O+6pwEc3fLTmekKQUbCv
GChxB1x/ho0d2yl6UJXUHx5py/2QZHuOcehx1o8V9GJ2LTvBEV6fVBoFHTYQIheeflBjDmnKfmkh
fWFJf/9ciBadAgCAfnPmP0pTb/ijjQrYexm8vz1gRhoPGll5wvNtzHJ7Ehvux2vU3yuUSy8Fgb/z
O/uIxQjMuSN7uGrQjcMgGyf2CPGwDIHIXEM2d+d4dpJfVOfmWTXh2Yt/cpKSJqOiD9vTbVdGW2sn
X6noikxIff+8yUUjJ7QzL9sJHgG1EzZ2D4llMM4q6W9T6zysX5Wu+iV398bNSSfzWwl0MHdUIjlk
U/pQ18keJ+D9Bmlug894cbqtVgkGqhPRCYjqMYl4Lx77n5bQdZ2SIFtubpek2vKIua44wPcUPzjW
Selw4ryYHRPQnkvSX9LNSEeVz5Eejk9QBIfVDuRceVbQRisNWQQP6VD9qhLZV0h/G6Bu9fAmMF4F
LvomvSilmS8EbhpU7762Ak9m16cLZBzdiAvSm5GYAeZ43sVzlBEM4jaBuqTCESTlAtbL3cKT7D2O
AkU9JfdA3csGCmguTryWDxjif4Hqz5tNn/8zUUG6bFfMJ8ffKCwRPUz7DCvEBEEu97ejFnrHuG/O
K+r58rFRnwus6xs61oOuWqjSbB2tLr8MVxcM4bqjXViqRTkwPV5rgK7ADpAs6cAjJBAwoDWi3YyZ
TqDP9ku3sWuX6gq03VyX0gauApXYe7AJ2Mpwnw7HbH8FpN4G+Ij6KjEp2OXlbsEe40PiVE/zI6Ch
yhzdy1ujc27s8Zp9wptiFDPHIb1dcZ4m+4EBS4T90029joWk9xuDXr3MaQ5wz1xCRRdxr0WX88va
6ut0Vw0ncBYBHK9nO8tKFKK3/0OLaY29kAKiEDfswObpzOmJZoQgO9he7LOdpd+1tK4RXT91ILHV
jsyiHz+pmEUJPfktqd2TGSs9I6j1/04DLmHlwPi1oSoCZ+K5X0yuVj+KsztKs6k1vjXcXDnyrHNo
YusF66ftoWOl8jqzkvVzJLC+OAHxUtrFNW/zRc6h26hyanjipOOfRYOfIL4zFJlkpQJfgnuPBfSY
/15V9JjzAAn9XC7lZUQSNfBCiaanZ8i29oLFNJ764eb59stp9NCYHBnBsJZ7i+N4I2Xgdr38kv5X
bA+4gSNMzb2CZKcXKpoF9EuY7sGTdAsTwG2TqKtYwP+YSyPAEFgZsW8L4vcmxinIcblaDQk3m4ME
l3HCv7zvvLUgUL0zfbe5+57S0ULyMopPm2pNEWEudAel0pvLTFF1m2dajlxmOB9gzeQnZdgFMIEO
IIxYaDD8KMhjLI9IqEPdnurHlIYVvF8gcZJeWE4EZ4SyoIEtelxniqwsXHiVfn1CGuz/gGwSnU0D
5en2ocHsAVca8Lag0k688yZu0pH0ojZkx+DwbkwlBh81E05Fr/7VYUaVbt4imh137t++CIdaB1Bx
V9J5qCjxRm+q4nFAYW8/shMqHt5xUy9j9m7wuoEx6O1TTRVFPzwQAxmveqzlQbVL4gJf3r8Uc7hn
fT6boiG5me4v4ntabayCS4EDBcZH7/tOfs81kouBxuwQXD4O/UshFfbFV0AjS2cXopnkG11FhiCV
qLFMTDK5l1rSn0kDP7k/vj18hisf0KoW3mZ8Kfxg0HIc88D5ZmW0krVC3jdY5W9INMUEA1K9YmsH
00HMnuM65ABeMUsQ41zpzgHydSWf4dMiP/jBHnbAJsi9vdtVSfSQvRP2KW79HNzu2688qJnCiKO5
DtRDwzErgGwN5THQ39/r0X500hGfLVK08ySwAlSs/WLDOGVI7lxWH5XRxApicqnHjLiGOxFAKGtW
eTDwhO3LOz+J5Nbf5kszMfI5hp+72oeMKiirbFovsB/wbf3RRK9fKG3eoWI9tcd8h/Jik+8sF59I
86BI6i5HGlUuAJDH13HdTRsQCyK+0BPDwsBECrMUC+VSbrkdcysgWdWXIL3Yg+i+bCjUixLroSEj
HZI2YDEgZIKISiI7o6KEbiYZHbuOwleqFd8BQvmd2bTnKPdDjDL/LE3q/SwnRQhYcHhoGtLKGoXy
xi+rh4qS+QvUuopRjd5QYHq7uQFXVizUAB3FikR5KG5aZSRc7ctE5hmRuJZaFswvYW9LnB/d4q4+
sgFLG//kmEjqRyAAz/4dEW5BPGPSTPvYPgHXh+js5MZDuZjLXwPV33NbQuYD6ZZ1zC8HXeGwsKyE
O9F7V6iB9g9dxSVBjKu2U+JK00QaGH979zSIWKM/SwTmXnCE7mW4VaJ+W9uBhIRwfqKZavfShnEi
gz71L0Oo0Z+CfhZVSUgGi6BpohwJfwdh7nI5pVCsEheBQ7eTCJ9a/7ByL91YYhazt61cB7jxzP6u
HAxPCbqthyWfhc465tB0X/afuQviiAok41Z/hhdj3ZsQ9ia/rC8NEhUsP54jiTZEW2c/pmRGHQiS
vRWcPNDmkuzGxMe2GSKmjy5BKv6D+uibLle4TdOuLCaZxqtyflNJqX56oFBYsAI1gG//leEWNrpY
kwc506MSLMuFJ8MqzVUViv4tSG0Ah431/IZxWH8Vagn0DJlMgBli9/LYTSatRxG8ecU2StzTGseC
eg2+E1RQ1bAH0i0iqalHlFi/4dC0QtW2Rye9TqP6YoVzzLB8zb5tsi3Wkrdjr3Oko0rvn9IYE9LA
6D+3nk5R68DOD7G9vLoA3BPiCzRYPMR4xLXKiVL4PTSlULIIC8Pqd5SKDv+SzvQoRXOwVcCRydpR
JCjQP1nxMCgahYo5nA8rfg11pfYnUMbvdt1qxVM/1Nlw9jE+NDUqQC5L8sohHaawMkXbiopveB6K
gdcgu6MTRXSGzJKFiIlvjY1rqMW+NTa3oudcbDh6Bg5meBgypbmFhTd8NK3DFlH+PTr53B+v5Z2Z
FvzBSGDhRVdmi+CR+mIonWLVg/vHcjNvt4vfvwhVMj32w84s54Y9DMsSFqYTcLw6FdEVlxhZ6Ck9
FSUMry8Tzw6GXK25/Ikt89uvD6qr3ghGvy9hbViPEExZSJ0/sYm6qnTq9ppFr4YZeFs9RY0jJy/h
2mS5M4hWEF/r0AJ6N/N9W2oCR4yABjTRFgUFRNtiYmaR5wcsJupcn217xoJ8MUxiF6fhHE+JqsBz
frwDsB1yDu7S+T3VGPnnkM/6ZjFE64nloq5p0RsQbNzltAaVYNuiQ76Y8z9dAdKaNXwY+plDBQyD
bIw+7pvTJ+68PRvVPAyHAi8L0cGERqB2qQSUDbhdhQe0zhDqY2UbKR+vSoxUvLDFakPKNSkKBhcz
WjmzQ1RocKydMPTdh3vka1eCAI5ApSGWPdNRyrD0++N7DtUSju1cqzMuvvWFZjqMOR8HSyQicX2A
TZeuOEkJgLh2AdZllQWm2IN1r8xstIOOs4zhglzGRZdVY/469uglw1URgBx2AOy/dlA9q2+LtbTw
2M/S7lsZu25uQ09IBaiZaKhKQS156dMc9JXHtEcf49JQ16XGNt++VVuTldXC4slct5OTvs6ayoLg
VPEAnx5bPzF8NrAgYoJm0GyaarndHTIdm0pVNkc9l/0qpC4jl7plP8BqcaVg7XyQZeXpp1dJbIXx
R6bW+MOu0E2hNkr+Io01TFJBleR2HBSoGtrge4a3XvxGJU/yUqn8Z4Zw9aS97UiEEWHEx5GCgxRQ
/K3xvZsDpoeS9HbwNXYyx/z53FJiTLL/ptKbI1/uNy3gCEkTqa4xRGwLFBh+m003d1n2UBxHDt6H
E2EzmwqpQ8BSH4K83eUd8XE4Tq7onxQ+2OzZxHUVCmosJ01woQ6dHKhTswJAf3ob6EivYskToF2q
2qDOcQLWC01M8LFfi1iP7KA8EtEe7uJAAaMJdSjwzUQ1iBi2ZaY4YOK8ivIRTFEx2V42D+APgm2F
Am34bVIXLzNiWF7wxoN8Qwpp5p3aqrDVud3FxjLP8vxO7jK/Fpq3VY7+yMr+XeRmD+RXWnVX4dsH
+25Frir8yEqHxzB+TPits/G0A7a/HZGJS5OsIphockgpCZFjF5iZlAiPHjQ2AHCbws343LoNqJpj
hi7DVC7JFFETR6dvgFLEEzfdoU4cYT3UqT/oV3jabTzws0+nb+gv2r21rA3W0A5zqM3lRxy8WJOL
tEsDEDvkkzx/zJlxZs4hhiQqm8Yfwtm7TJY4Tl4FdjkyE+iCR2j8lbXmh8/mVgeBXtVSZptQgy9G
q6HHhppVNKlgl2jbULbuSJ2oK5qxGJ/d3vXi2XFo/hU+Yv9AkJ81quq/cs4ieLOTmB+GKfixVdlQ
dTiQYmYw0iKqwwVqkM7YZIhbSNTPzDfVYzGLkMPU2QP7Bntsw8WFpUhZO00bGC7a9DUSQRj4Bw8t
FVSvQmD28Fr8cbJz6+Ih1yQLIiQV5qA6JZXI70Rv2wxlRpJBNLC1gic+uZYAxyK91AupoBDtME50
7ATAifhMKBOoEsMFK49juCwd1YhqYljXaLqcaEpbSuFg9uCLK7G8UMY1JsdOBybRW+EzUKBhIWWy
gq2qtPcte21yhxhrje+LXc9qs0hH/cjuXpKvUo2AFnWbdnzt3aJ47RcISZ91YpS10lD8u0Eqvv9J
JZkFXXOJKkClbgvAglpHcJvAsQ+HjaCMyFaATwn9HPKLjoThcGwQxWUvrmhLhW9QmVnlGXaC07MO
gHO5EeDKA3coYhdabTCKH8/FCNXEm1BpipZ7lBbRMpvuOG5KU/86SfLK5tdCx7gdZRZudyre3yHI
jM2HE0RznQwhse3PCZG57YZ9QCySUHf3rRsraCWkT5V6UbV98kTUJMmfwYdcu+wTsp6XYfF3rcGE
61CSN3ZUk4CkTotQynv/tQir5hgN7/wl/DRklLZ9U3prfPX3ZO5TcSgJuq8WK+CF4MFfYfyGTYGB
0Li5Vv97V12sBujnFIIvo+beeByKsz5Pmz2LpzNgPLvrEc82ccSOC9fqEboEfvIu5U1zydfgpCQH
5ZeYk5lQERVivwZQu6SGznhfE3DbBlIGFMbABXQ8LWF2j7OEV1IfnIKKp8pRtgA++1HAtWNg/yO9
vMEVnXWYrR8/x5HV6UCe4Iq1r7v9oKxSiMNFFb+lQ5DUWqWKZ5L62+WDArgLcTfsiAnHIj68JA5b
S3CGIWcjPGWYT9eWcUkfZ8F1FpPfJnWs+z5HiOVFGmBXd6peOg2eDTIcj/+ZF2HzAoBdLcu+5EFJ
lM2fXWL7Bgdjbf7F06dsELmpw1TD0p9G9+OjRZqQBofHoB27hJTmQZIBJlmn9dqMxGDMCSG8Fi1B
gpFNRRUegM2Lbr9oNQhNESharhHxvMlmvTNyS1lSAXS599pMR1tdGrbN6gpPRQPERlkLc6GcCtKz
YVQ5+vOt3waMYa9jVZ1t1V/NVo1vVW3Si25siaYyhvwqpJ7ydD5u9fMyk/+RD1hmLkPHG+iDfbQR
uRBlfGrph9/FXc3icxYgZ1eAVlf5GusXHN56JXGB/Nb/FQBJw+Lq2EnPAnTdhkXUaiuOq0kB81/o
aSP3IT6/pTRXXCMjjdAyml9uPh8Xqysgae3Pxs9CpjVe2waznUdoL7zn0OSQe2t1Xp0IWpbxMEmr
16JWiD0HQRiYRBsOjzzTXlbZeGDKH8W3dYcaJhKC/t/FdAI58gbxIrUkjKgd6QzhgWKoNnCT72zy
gvHYYfNOWv9BlefJoXMmMiWsfF/KR+splON3Dhj39K1wN9etG50fL5MMTY0Cfmibym/w65eTYpTV
VGY1tN/Knk1E+lnlQemJF7N0CxQsKhGca8/NxqjNd65fsB9IbkTkVJ0kPkwhgWmTlbUxw8oZULE4
EZN1syMxZdWPDlRXWqhqKGXzWjNFRi31NbFfg521f3n2xCok/xlGgJySeA4VGpnIXlYMwU5By9r8
FbHh6glnzgUt1bOrqt9IBh0myeQeuL9z1D7Urw/84wWc3sM7fU/OaP9AbwHgzKCN9vdJEkvt7bE2
gOBapCIYeUv4bqrIOis4AIxiqwmeJP8UEJW0vfB/5dvvN9FO6eKkbDvrY5YscVhVgoUh089ivv7X
c90SGUx57z/zfzLIOyYSZg9jv2oRPVosqmoytoyhxt3kcqQlgaavPxaL37SrKtWuM/cGyH72jvV6
+RReqvnCnlIh096o+qvOQAnhvWchuJ3o44Mq02VFMpmFxPQ1mGh/lo+SxU3NgAjmw0XVTaEpD0eI
GkdH/vDjdrp06Pplm/8Wzjk6mR9OtUphB+5ZWgJNlhHDK7/3OghpBq/Lv723v1MEN5Mag+lnItpS
95+oATGfZuBgWNfhERlHLsK1Kzo1gVi3Das3fD57lzAF6FWiEKOTMNpS464Wzj4f9tEj2ZcVEyHP
F1hPn1tlCypnR/1ytoecV24lb90/2JhDZ/LPg2eUrN878/cn9oMLBky9qFx/5hx7ZqVNRRPF1eGU
V7vhaRYlZJFJQROKwU1G6WoWzHrYEVXk82zNSd5/Hotn05YpTPSUsPJ3/0ubgecL7D8W6KgwRrsC
GolJMnksvZfGEXuHanbG+WsLwug8SDZXRZQOSAJfcxRrdVZP1hNbQhvLyZoEWXdaQJTOvA/XVujw
hioDUHaev4YQmFWzXwOOdkzPdXwRehIggqWVL/13zKcXyYqj9+r5359gMr6PYClU17FM9o3u17MJ
E3+xm9lRX+tdV0VX2EGGNGsanIG3eOxIKs7K3wPphG+j8DKRML6a8NQ8Ybi4tQuDu/OCAQLObX73
Q7xGrxBu4hCuTg6Y0rNfeZz2JDPOKxLl1CVx/ZP3bHTDGOJExFZD/9oHHBCqum2hpjjo8cVxnVHL
e/LKAc+lWksCC14IVqcTpwHp7ldNcfkrp2cjjNK9ZT29loiRWtcA9KsddDudUEfmlFXKjhmofeoE
VL0Gud+83+cHEV/Aifo83apfivoquwr4nZqNdCrY9IZGltezQudf6PV7f55XUUNX4JN4QWrOWz2h
6eKgORT5bwiGJZqKY+VjWXcHAQif6x6QWqIa1LEMFQSF0lmCoQm5M2Cf2oOXWCghug7uG2/2B+lw
KyseebKMlga9qLtGogezcxevdEHpw/RkkxeRSKtegAo6qLsk5+WzM845hxDEhoigtoLI3UgUtiqS
2a4hYIhBxC2wHUvTm1zV6CU3ITvb6JE6X2hfWEZwljv44WQDP9CCMTOG6fZ8uShAQCQdSYJJw+CW
I1BDA1Ib11v6WdneTcxAzdlLnWt+5bCPH2K7P093T/vRYuMsJ0fa9/7k1BGs/gv26pmm1Wm8Pc4R
Ensna0lwRIgnFpBoO20VzDKcp8DCYrc5eId5U/BFsqE7uEqpaOxi6J7Vxg4fPtHf+TaChW7qy7LT
QGeV1SPmH18rA0LYEtoUUgTM0r7al2frLaa43LiPsEjbLqj2vhqhMM4W4lhVIGWXD/ZlQGbQzPeU
AkO32eK2s/fOr8dwvDVfUK2k9ew837+dtOqZRbql19hVy7SPsDfAjKCHHwNNH3+3Ccjf2pncF7GV
tAWub1ePERsE0QewkdxjxXL57lm2dJBw3leT+teZU7DfPx6+1D+lAal4gEVEAsOjd2udpgL6G2ud
1swg8dBJ7nsekoXd3JmAeyjTN25gwQh+0KPQoZbeBv5taVyVdJn66Y+9JlbF3If/gHE/YItswyEf
pR/G/Qjk1LCvN9HcXtB8+ojClaiiRhXCm1GNfuKmUuHXGsz7N6Adu/GYtzIQR7mFrdjUj226FFrv
mfc95cbrL9xBN9gSOOiBgGWebqvGiv92Daxf/dJQENfRZbAlHPR9mS8OSIIfhD3ludpg/lKCMQav
nY4l8L+n207YUpbQniop7pRCR48NrUv4o6F/9XuBIsUMau7CKO5LMP2ody5Tbpc1Hun5yDdIz5eq
c557ZppGcQAxXoVNAtV6cfFjU56kvXU4Y0Em3IFGqty415GhHPOSPRpmPXwD14p9n45+iSR0Qh2D
oj9QOsbMhz832fFOMiBxEqAxYgRxbR6fs53YDBy4n95swxtlsnhKn5fkNSXVOdINlPfXGpoaHdTA
YdjJJo2HWBB4qWJtcHUxK9eTXjnunrxNu1+YB3OPBwC2AQ8YNlMPGxpfzdqmkPtjwkCqPaId+jtW
IPbcLv52kXZ7Dy6y7kTmJoJKJq/ukXlj+H5hGNXeTgqPZf9+C7mz3crQSJAQHrZ0v23NdfFzZEin
noYjrVbTuHTXtl/w31ecYOJgd7aK4yLE99MSSEn2WJjOX+I4+OsDgPikQEODaEpVMbBn0CHGqgin
f8ePoxraRs3b/+efBXdMRxdKW8JIITHpgDd0KNop1f7KnMb/7Q+NG6bWIj8Q532D3l/2YNeCYnhv
2r1iHsRl9fYr/llidEkdpUCrENhVGL41uQrE7Fxmou/yBwXz5iLmy43WfPo3S2MEybPOs8cWmJy6
D7UsZyhLVU5tunQrTqopujgn+fG+//hOfbterYtqAdYVjWSqAm0oNBO/tfI1n3OBeb5oZk0CkfCF
ZPBT3S6ThaS5c/hk0kn4TX+Eschmdmb68Gho0Ziw8aC3EZBKLl2BMVjbUglqivEMnbNEM297JnyL
uD3H8J7s0/o9MPNQ++b4nmL5NJ5JCMc5YX10fSJW3ziN5/WkY5IAAS8MM7scUxfyjSWgsyXrGZE7
Ph6aw61HQpx5AAaqPl7pU6HzW7L/IAfyPWcz5kb+UM5WARC6lBVmADVZtKbCfNBItdbNW3dMsvfz
UTWK08qEHJV0lZNAt7BPXU9bXzxHCqgIkv9XjhiOFdzKXDfx+clJ3iI4w3MAqvqYuqsyrdhUX/w+
Y6LumHsgFd3FdBADum5KQPtP2rV2pQvqyR3VqUB5ogt9oYKH3HOPVn1OQSvfvVjPMSRqJ5O3uUs5
rMXQgyWTi/xvVcFqPUdS6LyBjFP7eIqqFbQeuA3SDOt5AYoVzjxw3m2eVPpxrrd/EvtVkW4xAlfp
ZNirICY3690AvarTk3chwfWDp/xki26WyV9mW7UGqfpHdW+IIw5P202+JGEp5AthXWBbcxMP7S41
OqsD+9JWpIrLu7wUgqiQTywht22IuYxLuj6S80cTnBGII2shIRU/qx2J+YX+oiHi6VZ8WgTDlkpw
qJSwRRu2n0F7DMgqQalZxqG0n5Ybs1DNsOjZKoDbpuvA6CyuSdUVx4gRDuhlnHvqYHQxfScyrX0y
AZMotlodMbCdsF2bAycBYoQsl3uDnTOdJQoGgLUFYZZ4uY48to6v1zNdtTOjG6Yo1npOlMU3T253
eM2B1Yc0JA6/OlIWaHxlQmgFcHFWOLqpeV73KZs7u6JOLfQDK3Q7U3TMuZw+ngHhxxCcrlu3qLe0
8VjQHJTivSCDIlAA+zFghDq+2VjDj+Y5NMTtX8QrbPLgo+KPgQag9ikvmIJHNovVnx9iXESI5xeM
wavmcjAFOmKyhxKD48aqS3nxmxszrlpBv+gtvdHn/V9m+qk0+Jlxuu8/HEMb82mn8x8zrAbveppa
B7MvxA4MhGNngOPzXB8JXb0tMWKb/dX/kr1+NaX4RLmNRNO7DgCEUaF2XEpXOzE9jWk5tQYQ316Q
dS/0hFgHOU7ujr5da4Aq7qMBQ5k5oQJZicx3pF0BzzxNal6xPCsjQKLa1aVdm7sURMlEPxmH1OWE
EpSEUcsnVgXA/ka5fgHWA1C58Lbvo05kbGVUCYXaKv+KbfUGUSfPA5LQ9AVFzEPcIusvz5BvvrPo
8/nytk7PxvnYercowrMQSr4V7HNzJOU2LDVgxJGOmKba5PcMd3bl7n9aML2Io4+1/viqSIaVTJOV
+DTzoLlbiNzOZ/5uxS/8sNBt2sSigu3us2d9LZQ0sUb6xRrnlFOd/V0hAB79dDVvOorAsCKGiuog
jp33VW/WdDXX6P9WcWLhF8lUyh3ZGfrkRsylE5L/PS35OINIUYp4MdAeWHagnHJb/MGQbR1k3WpI
jZ1/Yu3pqCRo2Vpkl9mps7DKn2B4wWzV2BL160xrzinGxyrOO6862pwr0Kp30/T1O56dybSxqo0e
o33udHerQny6m1WwmOsJGAiIfbYS5GdNeeoazgYoLp6uDQPvWVewzkWGcnGlNRlqXhLTlQPS0phY
9rjAsg/HbdQwN8PvYBZS/bv8C7u/G4FDZ4a7MPB2KyjHx/Hasge1Dxbse4WGFKj8Y2B6wp2rfars
jzTUVWhDskErQ5dbTlnf6ShymtsxwxQt9UVrv3QvtM/ZiacdGUc57JKuAN9RDSic78fxemlrUyYE
F7HZyuc8h9uAZNBwpBrSabIlrRh+r5qdnFD2uyfxvMj76BpCPHe9SLBIjexQSkHtmdcogeCzB0y7
HhSI55FH5vSSAcvnlj6GtAOZwp2vflObGEjMqtHkuJQoLOX2y81PBxRU0zxuZ/tCEt+SbfH2hhHR
IGb7crZvlXpRsoYPq1OYJ+tJzNVDhbRUx9WPtx1FirWfJ1FN6/gkti/yMvTZRW4Kox4IGHNa8a0e
MoLKF2vuuCCqEi2VP0CDX44//1yag9/nSSe5wpkcI2+kDAp4O/XtGNTgGfHjx6OXHgywUYla6UoP
gpK2GwA2sTQ4uUJB0RQAS+1Clf5T/v1v+cfxK/81H0RbEUfltNxGCi3Lsv9R7oxe+YwEKWc7wKUV
GLIk4iZwcdNP1fpeHE20pM2PEfmkrazW37nxeMeL5PfSm6SDEbvoAca4GvPB2tMAwgTO9kEuEYUj
NSrJ/egI4SzG/FPUVp3m8oQ+Ftd1379Dj43LD0OV1CDALwuOAyeAubThM6VhTbZilZAlwgKx0vl2
aRmTGJaZBTCtR638kaBCQrKmLGGLaQS/dumg9cLGaZFoZ5lpcJAxA2jm2oJO1hO6j7j0o7oDIKik
TMJRkeDlRc9dhKVB45sLEYw2ZvIR7+cVQm75i4MWmpdG2clcw1MemU0RBsSPQ2DrBIA+6IsIdOaN
kn5RvfD7SmVFzoncwFZ6mCN8uskhVO2nsMwv9lEqqoBhPobhZSvwNsDdI3bwzISF4Aoiy2gVq3Au
OoxLVbhlsFDiJlaKfdvxwWFQJq27FTGj/ac3s7ESOT04hDqdQkU4vl53vT6AXO1wemN2pQa67Wvt
aGng2tsbQFdWOdER7n94sHz18I8EfyimBar/YmQ2JV8ruaHd6gRur3gT92rRZCcpzwyDj8W0m3Fw
YaISf2rZ9BMm8+qm5UADIZFlhU+q0OQT6H96Sm/lSnQxYT4c8BHIZJgY7yQ4sC7x5fru2oaQGnCI
L9LmLyxjjinL7cvjDNltinP7G26VgXO9PUj9DSqsiRrRrCTMVnOIBetHOx5fsvZzqC0eKJ88uPQj
T/ZWpblZH5ijSgicyC6D+fsJEIe4EfPhIMfpzku+xEWA+0TZXVHrozTKz5rWzgNtulPezGh9pIKO
58cGwDZn6f5726jWMNIDSF4qbqTJh6VQyh6XnMFl9ssUf3QOvOa7AXR+Ecd3UjNeQcLItctEHFRi
/j4Wn3mnPvh0wGnX3ZtyJoBR+ngjulcJC2OimGtaRUt5udfWoTdx/sIXfgoHZellyqYNr5DYu3Im
7Og5jhphJvYIbW1TMj/V4f0ObBGjbhbUhZNScW2sHu4u3BruKwItkq0qPHp4Mxj2VvL/rj3UUQYv
HCeBmma3vv853lFGWoM1ns/+7gxooDwxHTReGQ1xh3Fm6Cjk7MSYuFg1H1Lg5VlJsmU4mfvzCY1t
PxeNdKU5Z0HPnBKEVKGcoR1dq6AAEQKxvLOywBNrwTvH0jAKayFUxwPTycTKKm24qAlbH5T0q/8y
zAQXu/ejKOzrqTmHhlB2jGq9irccara+sF9DUQugQVwydJG30kE4h02qXoLETTHruFXGOVg7aFUU
HzwpFppHTDVYu6HQOjSM+YcfwlF4z9ic0uHoqy6fW9ArT5wcR3M0auPMHpxm2W/cCNdI+k3NSYmW
jxC7m8dvH3zscRtOoCxOs5rclZSY8RrxH/zgmjmLr8KHRhOsSSiF3b51WgpqnLOrTy6TQ9HpNVvA
CbSFXAGDG8pIkWQXJMvhIoa4NvlBV5cYgvvqGtcGakOAzJmsWBY/EQg5AGzfRQbULz4P4ifzYXYa
lMUHBbu91Eu1CFZnrtDgdfJ8mzVbVXG/FXtfqTV0gqZ5eIE3qazIXwysRgKBG0z9xVlRh1z8omf/
Jk9cMRZE8aEoKbAapRO+eghK+kblXp1raH/Ntb7sbtyXTrTkFcdyE4LwQFtp9H4WSgHKejNVxhou
bpP2cLldfTeahMWts5IIXz6JPPadGGyGgiB5Fk4nu6ihyGt61cO8fuBMuynwuFPvs+1IU0t77JTb
WJsHIrwVXNeEzzSapy3LKSjqTkTnJHBv3YEWMQBHcmR+WEDZNXW7jxMKZ+3CrZw49orCstXjGNhY
22D/Sa0dZBtMHuNCxgnIKuTPGzPnuB5Nq3tcM0pCUp/dZiLmObQZRFltCgL2lRgMdCFQABhlwWFZ
kDd84jiJIKC7r+VOAg76EPTI9bIy0zd8Go6MCv5o6Q4uoFvywBbYRhcKiBbOGfFVJ1Ika6VXLyCp
GO6AxQK2wdUDyu6VA3IURfEgAWJR7EA0gDmhwMXoL8uYPS5R0VvHmP+evMUQZ4PCqF85ZRLAW9e0
3So5qDmYwhJjxNTO9kBxta+p0f2GKtkHI9AZQCEpbXNTDqlLz4DspZD2S/w+ypf/1aYQobJILyBj
31nxnnXReX9zuN+JeC6Vm8sPA4tenlafbXz+00vZjG7RljbExDe3F8/DB/MUiEQy6bLB2hxbX5/3
Lkx/UriKNhw1PyIrf58rN6Z2yq5nuw5H1+Hzt4Zg8yAE5aZwkpn3UtfqmlK8o+Lxa+iQSBCOvnKu
r/fJkQfKaKC6EHLxzbwg2eSYwQpeFciXz853U6dgRZwPFtYLZrBSji4ysn3f0KyKCIwhnT98c657
cKOfT5lnepqE22x0nxeywG392q4ryim+eIEi/eQtL6irUe8+q9lxaGv6NARQnOSfcjPkcd++4WvF
ZQ3eMYdYv3Yu3sWbzPftef+8AcPY6mI8vn5GGDWkGHH6uTwa2NtcE1gagXbsChHg33bspFeKMKt2
8X/veiLcnUVNkF3kTNMMejzEZ8oYIncBA2y0aBlyVIjaGwoai94ChiMy99mkXOqpDUYdIC6765cc
FJqIZyytvlrdgkpWKFHgsaz8gj8+sZxDQRR8+bqy6HQrIOaCUI7YnrICRl/IORO6N/qXI1brcOmO
YfahpysEtW6HqGpO3BVQNjjkK42/nVxhVUNUAqP4wFOpSLLUugn9KKAWwYPXPWsqTinL14uNLwoL
66HsyD6VmLQvXc28IfknpSLaIkefISjoU+nReEbl6LDE9JtUdighN08abXFeesXWObTxAjb8oFho
EsvEP80sR8Qx4yk8qpSJLDt2l297yi2TtEdaj9BZ3V3Lk4H5EQSdIy1qHTjp16hhB2CuJgo2kbMe
7UTKW4NtfaofMzJg7dx4XPJB04diAfNLKdHjvhYE4yu8/rAlgjYAfCxkYaf09TAI8CQN/Sf6e7sy
V33Ye6bIpTglyqAJ1jR9c++q7AcmOh75mdhsygAUn+ffvRvV3VyQ3G0JJRPy79/J9Izhl8iw0e46
MqmeK5OBcn9pf+tPI3fZ9HzUCc6h6ekYv2V6TY2VkyAz/LdP3/qRMpXhZpcnfvhPAh9RylV2z9x6
p23/SIPmZ2orEHBkEKpNG6l1bOdJZR44Q2Nfk11fHy512vE8HFCLn7M60hswYCVfz4GCSfwP3bvR
XJ9G1TlewnQLwtpMaM25Cgupz6bx7DpvV5WgY0nh1GpY+j9j37SVGrJHynWNiYhoznetjfOBtdkm
tLUaGawmP2Au6+vX3kB+rZkyIyQ1MVnOD0BwqV27FNZCzqPv9npthG0tGWSex7xOEFLz6LlPC3fX
XVb0Mt05+tsLaILZkqldDwaWU1qhHF9WjRdA+yyhUiU2dbx50tOHUjYHLeO88Ij2WDxEipgGGKT+
KdZQ/SSVXcw1r5S76BSVlnVQYuSYMcgBL2HHID96XO5P2UL/3X4LLFxJegDOVHF5gfYti1THinWG
JuXCfSt6/KIwsKb7iLzHCwGcmbczZuhgJ1oDPrrqbGZyGnEzNjwUdCkMom44t+OLrF8/fN8Rtf43
xprP/+17Z+2LmLp2o+xu/ji8sALGWQ7YK9XR2zbzoomgoFlJy8kVdc702JRrOjtQjwZZdi8I1xrh
PtjJOyClrz1iMPzu2bA1KIDEpKGOMp264N4jn2eqx/uukcnYSRny6jWBKe7IuAUy3PdGlzERSsb9
6LwQNmcdXoqKgUoJILdM9Jf/15z8FZ1ziLu+p3CFTxNUJ0YoIWdY4MgwdykXe4JyQHjji6wOmDiD
mVN17gcCU58NVZrqE916UOAvmletNtZs8esWyMUEjWM6PatyfW3hDmMxX2RgZkhRSnckJuP/IQ5p
z+rq/jCvSg4Jyy/WWbksd/RoYp5mRqwhrrbJBEnizjNOG3eMAuUOrYLg7j7D3djUz18L7TEDLG83
LbLHt5p1JstKVmiC0rW0RAwE5iIkGC8wgGQKDMShKiYsUM1XkAVwYd4g6un//f+3DW62P1M3KyzJ
iV8dB5qpQiPOke/z4E0YGsAJPf4So2dAm1B42uimxXsYehXuYs0NgPD9rcmRiinBHbcUDxBDXzto
KMBhN9PgSUhKXMmhwS/75vRYKz3Z31jkZ0m/rJ5igMK08A3A671levTFxxtaK+Dmw/a+WXLh7sUv
0VZpHCCbRRLDDK24LaWYoQuNiEpJnoJ3v+yAyZMjlluXAwpHW62voHwhOAMz0MYP7WKma0InMDOa
pi1xVJEgoGbbEndBUhqWtvM5oDDSsA7+kbyi9c4buqwgncu8NPsTZCVn98843da5P3SDxOGejgWu
VqRRBhuKvZnI4GL3uyfztbwcmwQf63OOBsB2/AJSDS3+tCKrWFadCgQvqY8vKqiQD6ZLnWAp8Oo3
48l1D5K3acLYAR7ClIanjGb7tNvVDKaYYW4DlDC8o4dMnw0LXaI3vv3Ya+sdb/5QNbeMM+UpxzYz
fSzMIkFVyKPxGd9bKcv9Av7sk9yMW0j6rdybeEVIqY4S7OuhestQZmwNjSc2DyaAghhLc/wlusZb
2Ie1HcskfOl4XjhAsw1LXyDHdwGI39p7bn5ysJe5cS0oB4NOgHn7Ycv1Kew7goMpTvI9ZtwvvTyl
GrBpKExn78bT7Tl06Zo9BET2cL0AdCueWvA8lHPXgKRlghPPGkXdaPRCOYM3W56VcVqG8SszXeVN
hiCpoc+02oyUjQ3AU8yMlnyHK2gjibj7YJM6S36OlrhwLga/xc+vn6VKclLxe2Li62s6w9n3IBPZ
zSeKPaStCSrTtCKAo3G63MHjB16DGRX9T8NhIAGr8c3MVEf5lD01I99rFBoM+FpHGOMTghMlQwf/
/FYFmblBmcuATPByS1/Fr21smfZd/SCFebGc/6WBcVsE+tk/nTQpoyA9CCcQtLA3+cDkZ9PneqTe
UXyGi2PfLthW5rcmNHp0PdBT89sFa/eAHamhvGrEV6nJknY3Rqng9b49ZHI2YkcN98lpmLo9x/Mg
dn72Kl4UAMEeP8W4puoSZaYl/Rs7EId9ur5/nzCSdymDy7xSaDfb8fe7Yv8kgVcEqlPLTfAXK2rS
bkrHAaANyMCW69PHgP3NCn54/OkCi2qs7f08JWn/CtZ/zJW9ROGzwuv360sK3XUXvZjOMgh5VArx
Td2OzqJmHvabmzmJNWzVmHK8C2HNnXk4QXT+EcNVduvaeMrBKuW0PD2f5ggWjdAEeiDgAwZLOZKt
651Hoy7N6wydcB42DCdldeOS3X7arMeLYU15gH1N6mLSST5QOkbmrx1OoaE9FpEnar3Sa/J3R2Y/
TicC2p2Ajl6bDZjH94PuvEd5EYr8MF+/3jhIpj383RgtjcUTVtH7iD/qhp/NTFQ7BeHyGNEt2HIl
2/wCaPsYHcgKftuCr+uQFCAJiErtlDyKLyhJNBZ1ybyJiNm7Yp5/iYBrbPHaRCV4b8N2gLd1uzop
qMRWHBCnNImPSWIqRulayytKZcuiO25t+Kwk7Fe2ke1xhluFB3INsYbSYDxVXpf7kmY8VbmCp8Q0
cdpcQD5iW0I8aotH0HL+3WN8vQtWgDLzEOS0WPfa466xN4lC/H2zweYY05CV5KO7cgYbeEFZKvzX
4QUAeie0Q3Ff0i6EOlPGLerHuignOQY4NYfn8ME3UjGF5hrmh/91iuWYvZu/QYYVsHOFDuTegoKI
Yrz4B71CZ3JEiO9gnXdgDCkI2cBal43vTBD7k7/5AL/4kLdNRlYyYwLSwmr3q7IX7meuXVyZqugz
nCiRM3F7zPmXCIfFUqcfjYACuh4d7w9uAXruiPkjZ6FS3tWO+aZyqmJM2dsvxWhsLzVhnf5h3lE5
0EtKOv59RW415Qe0QqMPpjXd1k/VbH+9APYKtFerG62LYcRxcAgJ9qHxGlu0tyWi46D02T3jjCwu
vO2sMjWEQNKcVQNnV5eslfLzrEsojLZ5e07Q1idqfn3nOfHAJNS785GfK+EZLMnWnh7y0zA7z2Kx
WS2qTM0pcChtOWaFH2s7f5TJyJxK4jrHTeT4uuPW5MSN/EgNc250GtH6FBlFh/l3QLxEoq0Rmb1b
MFryisutyfQ11HJSJgquEkLSCxJqwK+PwXMhLumoaBmwLI3pv+tJPqaP+2+oPeSL/3vUyi5iXZMu
q2YfjA9oj5WunnnV61xsTwJx8DqwlJdCpsPxhcRm3xUUtZ8cmPZFaON1dvCI8UEMZ2WohF1LZ0h4
GXGKKY7U6eyz3YMmCs+CNeP6rprwdQz+edsNqbj9xSvTMsJIpjMYrNkYkRxqBpRLrg0XbAxIeJMV
akRUH8zZsAbf86EZ0S4xjw5IXbviC1W6tSRX9yGE+dY06biFsQlls9KR1WRJtD/K2p/Vi0bUbbsd
bwgP0SIOWjtWsLr/MCpUwOGo62FN2IseLAXtO/wYe6pVTl1LMrz35TYUz3pMhT6q2edDH/47pGrB
4DGhsiHXiahNnDyscK7GmSXMpxJnfHBfEQM/OjjoHWIbMyDTjEdM3ZXvH2bf42FXG5xTh1kRSgql
EZPv5G38OwKHqUwlnPQ8cvyf6W7AQ2asQm8b+G4ja2PvrC3aWHo3IFAS2vZBXA6l6zWBOanWu1xG
AZACIA0Ak9bcc7ZAPWAucrkLcnsx7QZDh3iEvEO81Cj6CNpP1IzGliNZGpkHaRRcoQYPJ9wC1A4+
YtYhn1tfI7aQuvhMVsqusZwLd6jDF+tUKjepu3CAImGNqsBP8nAamsZ71IqKk5f1dc6DgbCMlSiw
ZlvSCwR7R9khkTxXqdJGb7s+UaOyyoprYCk2GZWuG8Ti76CZKDVsljeYvXSjV97TO/S3oXEaOYtr
OvrzOARubiSKCDq6j9Z10eVm3/HZSUqgn0kdNEmUjmW+znlsKU8JOe+C8DRYnSAquC8rd6YeI+Yf
StaD1f9Kp6I6mZYT0dFZ4ahmnyI8RN88HEbl7xqfh18p5Tqi8URXhII7RI8wXHWlKp+jvn6p1Fa4
qDmQQOoawrXHf92vmcOfIblgEYoYxLFq8OiMeY3rDtOdh586VsJmGANHxncNAuIzwzi+9A4sWB9i
CIwsy4ie4hYN94rWFo4mYt3mtaR8KFQy73RBAsI8fu+EHIhxOzfAhzvqNlkDSgaOfWu/0VhHvDaz
x3N8E8X/BJLa6YZvLnDGdWzMhNlzxois0nCqE/52JNQWgn3PvuerFDSH2K2T6TQcSQQMYuwO2YNn
7NVLbI78pNP+rHDsoNzFZacaGCYfQ2rJU9ZCYpCyLD0rZ/igW0XhIiXnDY8f+SRXYZYRrSLssEA7
2Gidk56KfAhNjjM8nm9v4ncfv+VMlUgqDfx4sRmSX6KnopMxQMaxKsl9PSmfccBjGCb41o2OULNV
LFyXMEXu9z3mhGs5O2U9WHM9zsMbysBS9yjN9Eu5kQVw34wbgxkSgpt6dHGAyLu6DlFUx1z/EIhb
a3sqowFl/epFcdwiv6ZrZ0wA8e+2ZIWnyNzSC+gY28/gAFmUoGQuezjOSe6dW90e8cVu+yvDir3O
WfbjrAShkQTo8Z9Yp4EUZMRFa8rS6lwExrTdomDVSKyZTeb2oIxEaxck6N7EX4nCQ5ijYq3AXZIX
bueVrPGautKuo9hS8dTtevVTU+At6XSgdIvekxXDwPVWT9PmfFYpyo0CVm+ilLAMYHdGsF59Q0+z
zrH6V8pChi+ORk9Z4+Vk9MniNEWGsvCtdd7kcq+RF4PGerkPRvGCeVchMZgfqWQhypoM7Y35LTuI
GBAk+oXfeUK5BlzEJOGQ0FUJ4P1/b9bLJlQxgdSX6uoX93GQpSV/LePTYcwQANHrGNlVeGX2z/cg
ArKi8zdQNUKMQzsixKfibjdLe5S170xKKOW1y9T2FOw3NyAyWX+RbCU2pWgtJfMR2CmHJFUgj1pQ
wYF72dJJLLEz3Y/OUEdNi0prTZq30J/xaDTCa10eenwrLAKass3zDbPP7UpdauY4CuKeK5vWJvqz
BXRAhDm/HUWwgTaQvlyX2CLXy4nEH87RBUlHKIpuG3yY9my7NJfZ/LjcpiAVomqcjk0XDGfCIYB5
TvKTdk9HN8QihCZwjo41Pp5z18sQSB2e9Wr+CRku1hFfD93uTvo0ovfSu5X7Psn3JrFqo29bsC5a
BcwvqFHAWQw2k4ZTfQSLP10rdCjVQ3AgErd5xZ3GKIEqXjCIdkOIjzJo6JXJMC2Y0lUKC40K0jqc
b4UjFuGATH2w8C8kxyEa8U5sj690IumXsuOH3kBnePWpiWoL74L1u1qpiF5+PwVVNS6GhE6bOMjA
SIxYiKFKF/syi6bYAi3gEDEpmTgGhDkRPl3ldNchPzo8USoyFALwFB5NzvoYvUydGKB9EXkYI46j
KeYeWAFIOqk2Yx2TAsy//Iz6L61nXr+JKfabclIRm3KMYLlLvvsXCm6nRK2L44azeP8Z8hWIjh/w
n/7trJOw6G8mmFOHrMfQrQM58BygnR6AXQq1VAupcfZ59IaNHkrYenPEthb6++ReHWQcsAAkRMBU
Z7cERwtZxfyX0SovBKAALyeV6VPBtWzGD1ZMpt6eB6h7U75hbH54H0KFdtnzy910a8wUf61qrGab
hBOhWde2c1PP+86l1ocsOkUX/rmR8CtxzbOb2dIBfYvFZU4qA68rT/EkZVw5pA1zCPBkjWgHBSQE
IJvk/2XsWGwnkLGVJ4QOsGlCLnc8EMtjAh5hRHvMlzrOgHHrJIGRm8pfwJsBNolar8up76Ql9//k
gI+ckATLYonBYqdAS0UV3fFglqj5EmdAGUEXGdifE0WzLV1FOAiEJMdKabEXs+HspKvqGne+81bI
qSvUvr5E7YZM6lwsfm5bewnEdn40KjuGjqrgphak68YowoLBzaIn17zUnTNmU7GlGoh0VxduleYk
ZpbC5Lg7mhdSNVK4yMFYIiRT8GXTZlVXrAvJQW3TToKjNYjqBC5lJ8dkv3+k9RP0qC4t0yqYq2tc
I95jQwHyRiMMVBFA4nsSKbIyyA03XDsDBfWMn+wS9yjIp+1/f6r1/ikl1m+IaYi9ELP+irdjbiVf
d/68txzkngDaKeFCTBnEc/7cUwft0OT1YThReeYUJgbzDAvf/8NrGhvyHzQaI/xCBkiFSQgiAhoX
Ank4XiqR70HIx2t/+6+Ndi3Y7xxFVI6cnAQu8aBCZphn1deb/nCZwzHOThYShio6Ff2x6qJoOpfY
ZYkvww24MK2LVb7tzUjzyGr7ROHQlxGW7bQshzvmYQJCo11Ty0mMYs7acA4s9hdtVKuk9sVjd8ce
mEt364IlsLD7+AN788yUEN5o4sKHZ6fALWvYEeOv7YkTGymVQR6+9ed3sGOFHq9AZodrlLP4F6oq
gw5WSpzU6j5ZrzVwtP1QZtdaYTqRAmwcakvHmNuDSjzY2cVYXQRwZ0s9JvD7oA52Kux+klcBnAwj
FYMvgVvelVxa/qM6IrKHT8hM+C9GXbtt4rafZG9tqU7Xlj8fCATfepoI1YNfT5YNJscavji3Qzu3
ccFc1+zmUsWo+v9rgrbbfoXngN2g2rd8xUfxFCeidWhYLOZOZFyCGY9yEQfOt/APtUzF2Lx62JM3
FUqoJBPPQiOHyIo/fh0wA4aWxrgCK3SsAfA5/tcYh/sb2vySGUhPUZegXpPYZfq2zTFsTc5Z5B6A
BxFkcW7yuhZVgmjdnP5r4jT3yQxhnuGmTB55IHrRB3wk5oyHyskBAfU2CoACuaRfaw9KgYJbZJH6
oxYmJu75L7i1LqRiyMJIcOyDWehLr+CvERNs0CGblhHc+jz5jwGSPFkc182ObsvYwcl1JKnFng1/
mRnrSTyXobSfB64WbsNtb9Il6LiUtRASLY1vb3duygwy6YH5P5aRljguybgf4IMB5/8R1jahnjsy
RXW9VEfXeENHs4AKFWuek7tOdo1hGsu12Ij8IB/eSTsQgg9PB+/meHJO8s1f6xcWal6sBWmFQUqG
gPDppVMb0629r6CDdrjXX+gyLo06AT0kpFvlHPz0fQZdCXgsIsvwjcKkn6EcbiTh0CSRv4mQuzlT
pIkMgj5LfgMr6mNflmAuoZAW9Q5kaL3lmMP6MzAezOsk3E8VrHlafZdSrl9FV0GExk2+HoXwvZVn
1zUw3fI3siZm6ZKwp1g9UrOI4mStGMpt6umurakpIfC2SqSUqJLxTdvWC7Trn3e//eyFs4dQJDu9
lWBPLpLzkheVGgZN8WfHg1W+NKH0plC2YjPmVTIqQvzqAVGBv3cKjADHFDEIxAszOAuZWeWgxim+
3yjBsjJ8P/jE1V29FFNc3Tw7nhyoy0B8y/gnh0+x8sxwi28sPGS6eCL0Y6hp1m5gCuj5paW81hWJ
TvAqzaxxX8H9rp/1PvaudA8t7wMivOjpkjzVEMtXSezoJ8p1ozbY+umr5NsvXr7UNiVKscdAk2DT
rJQ2i3QA2HXI70uEWnqN6qWBkU3C+UKDym13VK2xttsglx1Sf0wva8UtVWSA4Fmy32X4aLYqmYP6
4il7J9vF3rZhJ0183hubtRPix2AATdphT/KRLaDBQ6kWFt1ayEQRKEEWBV3y+WAsCMyG8ippISCr
aM6ONMatyICpUVYlmz3hDglTNK+5LHqAixzhmawaUpCc7Hi3C8duOPjlEJ/5kXWxDbzmnp4UcHyV
mVS6cMvf+F7h2ZVvoqSwEbFPU6e1Nwevw03PmLKXTw6Ru5qYPJMC97ZvLbbpn1D/5XxJmoV5pH0S
H6FtCIEGxF1fMmZBNAWBRHWptWLtsOUchENeHV43XDwVzJFg9UdcRoQbSnyfB784ehEjnBiaZvIJ
QFZkKQI8GMkzlM67YuiSb0zhyFAlmq9Wph9wTGinbcj/xaj4GaRkfOsvwrjVua4pUJ3tZ5Ruo3U2
VpSAPfOlYF2KlTF1AES8PWljD6UsfoQ9/IJ/WAdBBD6vxh8MJvevrjS3c8UV/FNHGtzUGG8WnKve
cDDcCP3LW1tNJ7WULNNMSgs0gn4C2Y0mfLtmoOnAKAP6jaodn37nlTSpA27I1MRzZhPs/g5N6ogC
y5po5bafz2dUbxYfkOr+XdNj7eJJkVEbpTWEzHgXfkHNIw2tprcB9zusIfuKSztqS3ahOcF12zSq
ZPUCaSBj6aD/z8KwmDNGSnMq6A55bSY+E91K+TwQd2W7cyHAZD6yM6O6OwgcuVPV/bPumTTSGZI1
H9ormXDRe8irY6IKh6eTBHssV97kuc65I2rzoTrsOaYkyUhUPL3hfEZRgyszqgq6y1iaCLQLb8N8
BDUjGEUZa2tn99fdD19tVulwFNEUjQeejSIJQMLsGL/FjT68xBzAFgT5/0Fc57qE3NmhcAH2sCqb
2L8ujh5T+0vgCxW/nCxS6O1XPdMG/vqx7TnAnmwvh8XvtWGlLQZdEEFAd8hj7IGt1Liv0DIodepA
MmgKyJGD031usHi/qmD11skGYCsiP9f9DSMdGcu35F3YQSPHcjI9r0FJNbvGrvBCg0icuq/MhEnV
ujjRIpXedCXg3xIgzxbhApSVAo6K/dc/Yx9ai7mRPyEP6omPYEGb7QHEFkFs17RNBwb9lUG5BY8M
3h6+a3Vc56wOu+92COtY+6gK5NlSupjScxd47CCYTkeL2e/7di8xFAcBV8u9ThBdavXIKC7oDyge
MceC+fv2X0qELtreU6r8bh6HAQePtAZkiutM3DI52/24JfD1o5BM/lG7UkGZutn7gB62Vvb28a3u
rG7ksERgPQAvMEgeoyk3O9ry5VClpqgKSdPT6O4y3ewS6NH5z5PU0ImjGHEXcnWlVf1++gLilPw/
wf5PmJu9MDouLSPzJR/jpEWlGOn/vnft2mYuOk/qjFWBhWmziKbE583lbGlItreS2x/HEKV5pvqs
XdIqdKnRs8Ra1TjosCLnP010dfqJNEq0WQgo0Xg1vf41NzihiOFCwL3SNSqnEFS6oS8CdoD5/6Xr
9Bgt3JQBU1tFCt4chqC7I1vh0DvF65Jpk+hBS6cSkMc8dN29HVl5/Hu9Vv6M1/uG0SMz5UR6/RM6
iuA8zUSx44UuF45/pOkToB4SngErXEHqO0qVvKN5g+/+PLlqiAMIC724FBHcZ4Q69wTRHq9pFwAE
qkcxkD5kOg4QoWfuYg6SjO2eZucCvndjRtLMF7bJofk3vPvVeNSnoYfjZfoEqYttJcDMzkbiNkVQ
KSr9Xdgzm6Av0nNDIvCdKERzw42LCMRFMBu006Ez9F4iJKh6h/xth8jfyUW07F2Sig+vpohxTX73
wLIOK1yRtkydIboGXxxuP0T9GbbbZdCSdPkQ7IUFe5a4nrw+5I2xWywqdC7PbBRDo9UWYZD6jFp/
GJCK5pw6o8ylLNcWdF2+Oy5as4RTrDsKTgU7vj4yIoIuYCo7qSYpFZkaws/bPKaHEORK+yRX7pPh
Kv01ap7gj2CVVFubsehzwp1gAztMIpQtlf7vAsdVPVjAVHsvhJl97DNpLxJitvWgFf6i4NIZnafX
Pf5TsC7DbDFPScNp1Xv2ESaF6nng2Aqy/rmLkjWvUmt+4/77+eimhAGiEAqQpkhTwndds0nDt6Rl
lI4tkYVU2aJodpkzWcwoXVBYa1SUFCPGl77hTHZQzllyvp2RhV6cIRHMTCblI8K5hNl0wqxTO04Q
xp+8ZMsZYQ7ZiZXDNCLlGu4s/i/tpzmp0tEr9+KpLjzNelDcTy1BIEG7bW0hiONMVSweMiHLCyeQ
z5omp+M4j8BNbRm99b4sBm1yX5b/TYJigB0Uwo7Igq/dV9e64qHiU1E+Nid9TpVpRv1FZR4hNL9y
2FZZrxAOHBdceMCaS5IrB5iusqjk1BrT2NfYcTEfpdfBxhkAXu+eSxAdelSZUl8NUD1mVR89LoUQ
jQOiEedsXXyBH//i1zP+JwP8mOezW0JtzXaa4+HThaRa6aVk4V0qLrJwdouLQz0FyjhzuN/KE/4L
kpSCsNpgiZEktYFPIMXK3Rnvnvs0shuGZJtDyaSytZZwo+anFqz5Ck4CJ2HvXG5xorHn1ADPyrlJ
9EnrJf8Qvf22OPd7/2iwQKIlbChRic+X3EtaiMgp41rTqazUg489efvEQeKjFsf0Gx+3Ll2mw36A
hQhLADzm2+KLtRNigMTZvm90/IJ8gVjrEbEEbqSs6415sjRNsZj1K7A2XaoW46EVkJySPiWAPsI7
wFUE5ai3o3RwSzLdW0eS+FNFUSSidJPbpv1oUII3fO3qC/KYXuKFqS7we+uco/0juvMv6/z+A9em
P/TsydJngPRPaRNhHHg9p5ekgsGGA7I70xVQbtvuKJkkMat8yj9a5CsAIpWCfwaH/ioJQLg4BBUp
/Ba0eGFECkbqPXa0v+2f4ZnIiFA+oG3gEZs5dXRfCvDKzZhgGuOol92OmrlD3+nTjzRDOY1jQOAz
QS6hNwIPLsq1CRGNVqTgB5gG8z4N9VJj82eLyL6Eewlff0wwH81UjeaEZ0QAWjoYuVOUZ5WonNGI
l/7eSFI5jlsYAEWFolnCYiOTyASSe56d5h3r8jubQiG031QyelqXn3BHXVp6+yrl078AdKaGmsUw
cpEifkzsGBvlFNV7Wyeeua5pVr5I563owX5jC9eFSVw4Yv+F+CgdnZpADRulCZoPm8ETkP0KTJ7i
dv3v+aOpjP9O1RfxZ2Tpq6g4Q3geCwPTv6Z1ITm7yK0EKvflt3wL0c7CDdhIhQjuIFiFoMqGTVc5
y/TGwec/GetUEewS/E8M7a9rQT5oGH2SAr6I18yif7VyUrlUl/pNem11R40Yus1Si8w9FkpNZJUB
HMOtS/6nNByPGeA4HpxDuHHe9+FN4CMCOOD4m/klbIP+r6/bCSpRmaNE4hFTXLSiOdUBTTAzSLIi
Oz8y7l96bSZWj7y/M6GQYA+R9trDbjl4ufMbMLdJcAYUqWzHjblVuumtZ58R2IhrppV/hWNVFHe2
nfcWV0PuVYnJBuCj1xkOuYcDeup2N9d7j8CXaA90luye/fro6B8q2nc+75O49bf+qZ+w4l/PAipR
65w7ZtnfpowGUdmhvcaeJCOeK4bdyBcae6A3TVo8BuZMvlaW4msh5YIbGZjWVd7uuSKqoqKcSGhN
qdpB5/6kzwCFMeCcsPYuBtErRAQ76idwdxlApTauTZ2PCM8PsWxRzLJfCvjsPDXqzBvcXW2rf4Ar
FfGFA+MEwi6cLJQqXqVCrxYNqbEE96lTiAogmBXiCsXGDvfwjWeSPMfpVJlkLyFgclY6dwvTFtgl
kXVRoh1FdrK8IwtzsFjmM3sDSoOlRr/Lr+eMPF4irv3s0eE1nJlyGsrBG0o0ON2XCWUozayCdToJ
+e8jOLKTHto2M/b9vax1RYmWaZNTkzthJMhozs9E4s/AT8VMCj2FTLlk+4yWTzY3Cp7Ms06UgLfI
ahDXaXVDDyWJl8Rtz4vGqO4l5eotezz2hCW08SwFoMzETlDnKL6u/xmTCCkhDNoXZT3irCn6u1oy
upZQqND/rV82OAkGUJzdesZVPHZ24KxPvy1dtsF5w47EpuI4E/p/VHIxM8DsP51esLtFQM+eDSGC
cqGr3WdBrNVYvEkTBOevZKBhMaJjBJSO3ayKn3zj8/pwdYBVOQOB13CmxbvX7DJ/Ijs749WFLUKx
m4hbMW0kBxm9mk+SjlhSUeSKZIaffZcYiV7QZYJqKB3NLYcULIQrN9tMKO7L7ZwqChoTFnW5ni+g
NL+h6gzHwt9OM5Y8gxgUDEpMQNfS74R9RGMOZfTs6eJd2fjFxu0abgqQ4HNCV0efQTx4jnaNSibj
fn+Sb2UCdiMCEfCpd6PEB5uhb7pPeoLAI/9TdI/2ipeqXE+9vofbIByF6Y4UXj6Vwu2R7IW4ewVn
/zzOXvbedaJVl+9lq/OzDg4EcOL4n/NglmB/pxLt6v2XBJfLIwEjZJSehvlq7BrtgDL5dcA9h1gh
ojmrp0PXtkZak2l3MGFNL5x3mfU+zlMp+rYhgSG+OYbVGKeJeHswdbS50PDvesEgvWIwIcD/7Z9B
EbJw485mssb7L55VuWYH1HUWNJAVDD71ytXO6by7bM4QVTMNGFdtOY9rCV3mVwUjnY2XqEYAiJHi
dco92iPf7/ZPKUh9ufwKdhCAl1Mf5Pi+kop1sqqtVI8hw+C2OxQthE6nm6Sl/lqmisHVYxNxJx7+
NbL9aTk2Pz+ebO7OMFCdxYjo5BU5NxfAoqPPJCCKHusGyN3fvQkCv1G02R551y1BaQr5hGmajzLL
fvQZuGFTigC9IkRHfZFHl7goJgNS2nNE5LEWK+4DQ4Ievsca4ylPVdOW229znapBpgND8bZUIh1L
6qrmXwzIXKUezBiYSA8yUYWJpp1nyhWad9szav7yVk4trCKtIvcfU9rXVNt9zO/FuAkUGItakrNT
QFLEdwDxxYPs/VFjhHYwe0zBHeml7JvBobBvHJtF6060vqmW9SMP9xZnVcz/AV4HMQV7aBDEmpYs
6PxPab4cepl2QeO6AsQiw9hDHl/qmihHGYxpwhdNbO0yAeUlcJlFSc3sZxswO9YgT3u8ORA9nWFE
hxk2CsF3sB4MNogof2dX+/0vGi8nNuhhU7SJfMbuZGqOUMTCgQZWg3K5e9MXd7FIjVDeOunmoqPZ
Ze6GOvSsBF4JKb6LVvipAyIpC2XCjLp7c6SgP8zTRYN9yqS9pAyqWz0FNU7+vUUIvP4z6tm2RqQe
vtaavgplxETPkuauy6eVD5z+AaTBnhMxcRFDZPinkT9iUCZWrwm0FzQgxTbXNNaL1CcI5XblNAuY
axrJTnPNQtWg4nk4Uq+OII+3EQBqRCesdbK82TrALXIX0hWbpCOCZXPh3eAn6E07hVn8mxwiONmC
rP+gvIqfhNK7Sa+g1IoHzUkTrystw+GOo5OMLA3yQbIhTqX4ufJLpLdm9h3bYHK6aSFvEk8xpneb
YZyllyK9TdQX2KHPB1XuGJbXA14RuPwgpvvjuIGyp1B80OiItzRgbA2w6GAMjZN5bUBjPTMRXFIs
l9kJeyfWX6DDoWoPWu8OmUPRWBqgaoGdgi9Rqg6PupgbPIFuBTWsgJH1c37Kh2SiGZ73xGcqRS8j
CtELvW1EU0XpQdH1v/9ERrav5B5IxfHTKUGm9DKP3df4RkNnVWitzOvkLFvaV7wQi2JqwhVadTIe
qFhMGG37jTaqRBWsSCtt51XLPazAASH/TfxZRrD4rpfH7NqWt5mr7bTXMaBfLpOB+zAF/WCfBgfq
9OMIkV31HhT8yl1VEGQMgSpP2i6ncVB6wpP0UlLddixMepOifAMkTssC3aCMO0lMuzwUWiIGMTs6
2hecoCfwq5T/fZIGHvm7tJ6nuPOrN0DvIgaaY3SbhqX+PFXex5qbNyk55qf++rCWckzmqSWOOLKs
VkykXcDX0ZVDlWOqb6AsZMPsSMcXR1NIlUNlWU3dzv7AgWR2/TnjJtP4k4fL56C+wv2n3qaYehBu
sJo8rpNKKQ19m4EolfdlznA4N7Hx++Nbb8ZCVCalGG/XBo+XqMGG35n1bf2ZINe1D9dWAoXQQILW
ZFMal7V6OEeMJTRT6pJ1dqG7SNADSLL7jwFdC0XzzLa45G6aDZbFtOVeXgEE9culsz58zDIcelVT
G5U5gU1apGbZjutDhEomPFxKYSnigIwJ60gTx1y8ki6Y7ILnFG1uMJM2Db7+pOKK+yTA+G5UjsSx
r5uE7nnst/d03izAwmBfvrL4YaiH2rEIbB52U5mgha3So/PvMKqIWzXdmMig6Jks/w2W0t1k/5v+
gCembnlmxS9wU4cwIo64HFFCtJr5AwCkHVxNi4HQ+tvQAvLIiJt86XrveVOaGaxN2e/AQ3e18JBE
05aE4NxpQWx1MqDP74FJrUBBk3JU1tEo8emrfuAvaNz74oYe5h7UqrIuuc8nyCFGmh60k6CJ1ZZ8
jvpckXa8zymquRWWnfAhafPDKj0u1GhlW/HRWcq0tNuAJW+CucJOcueeT5LjXaVyhZpMBkKAqfj+
RS4hlck/Rec0VlJxVwVhvWgDCmVNnHRAaMUsrzF4Q8XAQK4woTYR9rEEhkSfMDsH5cyEiZzv6yAl
2XqyVCONRig1zZ29BbwHf+/EyklGO9gcbcYk4R0Tb7dz+Mxy7D0jUHRmop/2m7rwKZMDrjiH8tvE
Ueznye6mwqITpM7UjY8l9X863mYFzBU5+nb4K1CUco1oquXz7XbqtulQBKCJq/eLn4/IaSvmtU6x
fW+p/oyairf82mqNlxNMNWdDZplrvCy6LvP1fWHebvshla7CW0NJ6E524esWbJhpjIEaROJtgQP7
ENN7SdbalQsBg2xKBpMINzr60HbTzX2jZ2Sq761ZpibJ4VefZpU2SETlkCHEPSvD3M3CHZNUhjBl
huRwY34ZleZ2VIqo6cqH95DQjUwHZD9AflpX+DKpH8eb1bj1mG/LcFSjVkeWOlFVzA5nuk/ujrd1
+tq2Ud/3NwKFPurB+Y5QmH9MSOH3SOmtzfpTY0EAMu5YVzO7yfI0oWAOTi4Y3BjOm/69ugkqzPe7
jif9fymG9jrk3dMp23OCI7vHN2IGyllcEOWT5nF8VAbpy1DIw5IxywMODFKp9q7QxlZpL53G303U
oxFQWDLNMDWnhnEXEohTNed7Bh5xmE4vU3gdfaViLmlyUXrpzofqbi0iE4CHZFhUr8RlqQbgfhh3
PoArdcpxHneJh2L0TO51IJOg2Goa/R3Ans/vsZsl88zaLYm5ilAnXLLCGT8SA03NUG2TTEoA82p4
D/p/3y7GXRy96BXg4wE3X7XD/zi7uDDU9SUJJ16ep8KfW7+MlY6vwKaLiMTzIXdnXfhsHKvKcKM7
o26bKnCWil0aRzm5ef8xDhC3M9PR2fBD4XggWndmEiNJoQoxo7rMbLIfdW9W/Cn1Gc0MEgKiWgn6
WucnOFxPuCaXl5vSfKRG7jtkJplEjr18Po1Wv0hfL8Jd/Un8nzcqX7FpHTNDeUIH+GGZUv4AT4tS
QcfUubZ/zXRnTYrwphTNQFXnreYha5wtvaVyG3fWqvECC/u8Qly2NvCIpXA5Fj8gF0CSsK88q6Ei
AiG95jTfqC1vIRFMb59xnl2zCyS/TpUC1T1ipUtF0gstYJqtbBsrc3PiqiQ/832YmoSzC96+lBaj
v/lIU6b7cFtXv2KrL9z8bHo4fOpIyGTOQJEGIIGJ7j3ohEQnIp9O7bDEd8ChjnJE4IWGRhopIAM6
at2X58lNXyq7vwkv8+PIGU3WzJ9oxpA8cFgSEUT8Bd+sahRr8kWMPMjvl+3DvIZPNBCTGX/e6U91
vPEodid2kQiFPEoWycNxh+ThsChzUZLLt8vTz1N50jtARfSog694OIZ6Cd+nmzzpVs0L0pZDaLIU
U4wnd8srM/DvOyXmvfkCJwowNQUGX/v4zRpz1/L4EcdWUODsVjYqoN6wdjw7TsuVBogrBKrzl3oK
6KzvpjaeUgrxpSS4rdO3eO+LMhEwO91JdsbO/ruvOjE7MWqk+eVyaMzuTWOuS64mOypIpbwogKfw
TWnuwQ/yQboP3wQYg/6jG1AVY0GRgUil5j+DiDmFrJtGQvwVlNUf3Vav9aJzToLbKxk9bbfDznM7
gbkhoCAnSpwPn+/NHluPt7mSdP6SeWa95x3bqG0U3sX8CSYXKynbXUWSZITMKvtBXC8CDvV+g1OK
dFQKba/Qwwd2uuV/XqSgMx7AdU/aNROY4cP9D4bUaqaz7J8oo7++z+1wftz87T8NLjYgMKvdeeKD
JIAGFVoafKlGfWLDgLTAZ7Odv49Sc/e2qJcOmoRBwx5pdB+cLYIWPBkL8zCe3/Kyd3IwUMb9tQRT
mnVE/CGUQBn9SeJzlZMmraNsPQpccG2WGV4iFQei2n+VwJ/n0bjDDNarNPZwdIqD7m5GQCZuhfoM
pkinktbBERQNeEjuzNc2RYZepTy1aYfDvRoLB3wYqYHBZgbxxQx3zO7RObBH1TjOj/xro9TWms6m
rqI3+bRsio3BxbesVI8gpRQFwdzobeRxc5JF//OhazCrBcW8rnBrl3QYXnHlRTgyQqveAAREh5+B
0EFe5e4I1r9zhES99XD+3mpj2JBPT6CB1URKkYuqKXZpq7NKCVc80wY3K0aEcIaNuTyFeW3JaLCN
GMA4Y+JDhbst+XXfU/VYJ2n8nMCASp/eJH3Tnfl5umWX3aeIlHbo25+Sp89x15jxVKb8hybIY3mU
PhTtYfRgvQu9Fd69e3s7xy5q/aqKIc/0wTpdnVD07WO7sZ70PcEBwJwv19K0yfH77nI4vHtosNvw
1otjEH0pFd2sdkgl1hpupTleReSnZaeIiYgf3ANGvBCPBqM/x/uxm4NgcBVkP/L+umENVnTe4UjJ
bFnqXoYGe39jmOuWTmIvyqi5aStQd0bdaBRzNWiE/Z3w3OC3l3HEqdCH4tcH4LR/w0cs9ZRmpCki
4mIfp7Q0qhrpogc7YrV4F93Jdw/Byft1dguVIOo/XQx5GYbrkoAqBRDytO9Jy2QKCLMCe0JmIviR
pTXTl8weiMWjaEgviQ29YtwbSrisyyz7J840BI00BGAU95ezB3whr3RG7cq0JIw1ax5CAUDHbZwh
h1HI16GOHZLOJ58xFZIUDrk70Wbs+WdDXGzGkvVjulBtjZf4iV2r53SM+OhRaO6UxkFrDqI3h55i
MGMf/Z6n13Nch8AWRFFHjRQADc2OXOiclyEULB2hv1TbeJZO6rudqcQ/jBpLv+cBJzkBgHLV+qCD
H2hDdy5cFphpYWWZ6iN6AS3enWgLf9jiJvkoHc19pXvTjvPcIxd99e5Jo7n8bk2tKd6P2hIvBwBA
Tp8+YS5mk92fO5/hXMBAKDWIBdjl4/uTRlwzFFdZoTI03hbGP9+RvMkejC7oJQFWpMHUrNLfqnAO
OUsGh7eyWNZbX8ijIQzwnAZiRx87oikKBiBze3o69mJMUX/+hHTgoog3eKGZQLbFwy9cH+JqqQny
IB//X2wilCwZiXIxOr+8c155UgNm6Mdgzys8U8+c4gY2zuElTVpZscCTGwKp3xFjsp2p7zrrXATH
6uJvlY4tVUWjCHN4siIpHAOJj262dzlwCc5bJQVh4yn60TcrkJ8vVrVX5LYWevl3UgnMOOWXVMSw
hsRo0sUczY/3trRLFuXGrfWDzgg9IsghuWgU+5fRr0uTcHxnDso5bq+Dd69TTVsY/2e1DPShEXog
E7L9qc79g8dzcRtjraSLP+RoW4jRynI8n9KHIaSMV+6eyZ0J4xJKqH6yeessODDyxZXfhuW3V0Ej
V9wcoOYVF9Hi71o5Y8ZpzgPDNi2WrSSndfMQJx1dgrpmyHtp40ec9jS4mkQjkBH6v4Io8jNT5kG2
+VogRNm5rmEC8axcXrLwaPeGkM1+JOC+08GQ4J+m0+EPYXszdCiLI/UlG6v6M0lKf47/3AiMVnqt
8XQuSPffWz5lEtsO1iGkk9rrcbHUzZyk44K/t/LyI7xtKbuVSWsbCvn4/ZCJ77Cwr8Rl+cjhFqTT
56n9eJfaBCz7qbv6CK1FY31SORU257X8VS0fleBMG1wYV1uhpOB6I3QTQTCyM8+9jHEPZEYhg5SR
sgujYfTx19Y6JGOSJKoz8WKOLag9nBCkxcufC2Ff7HcSzlSYCvmBtLvD1xN+masbwvGll0jot7KR
p5XHkVf7kezKK0oFaioLy1NzOXIw5wNjrR0eG/8cBFQHU+ZGpSsO7wi53Xg4rUxJhtRcNRUwUMoJ
2JKzWbIfN631/Xqq0O+7yfBwzgqRW6/ff2uVcmg0KE39Rm41+7XvsQPX1uWo/+yC3vygw4uSvOTA
x/kjT76zz8CMdr5EVubK6mdD1nCvXwxAeoQ9aHSk20YAOY4dt/E3tSI34NJhD5Xgr9beSovX69ku
UbXmDd97YhOcOqYt8USO1GcB1cYa4Sv9aERn6cq2vX3KBKzGhMCmG/fZnKJVD4BDePAh1UqHQBcu
NXPcxjCVN8pIyA4D87T/e0WNHVyVzxNCM3xuvXKaYhuqyUgPMkh7ULPGoD2NPwNJIAEtqt5BtOI/
V4kHDud7+XF21T12e930143TNx813tj6IcDyjBi5SOmosadyDEvxhXllRy2nPDus52WYKlnYMFYU
EF3P/gD2+iHLncru1yOHNemM4WL6MeBzttwwSJYR++TtD3G624jY/oBOQEpo+zXP2+AiEo2vCPev
erx4U1uXOSu81lbdlrddzJNTbYF2Q0NTxyBzscAZC2pAieiHcAd9tXyq+VL+JA434ODCtYHbFJFD
m7YwtDQCgGPUFNU3OwmowDu56UzKOkbJu/pipfsuqMAkBPFZXe4IWsR6QUHjIaykfUwRlA1GlepG
BeDW+4QcTjYwdld/znJFq1Prhg30Qi+6P1Zv+Kxr60titT2eexZZw79iIKsDFOJ46nxaM35/NP19
9DU1TFw5EeAuykfNpDpJKlW9kS1Jr0WwIh4yNN6VPYGoSRtrDG7GaNpAwsJ8KtjPfGanghhjzqdJ
HVYKdMhntm+HLsP8nO+dusfVwblLN3FuBZ9LUjzKFpwc1/TKsgNEBD7kYEk1pVeX144hLaccEIj/
v7d0e2FqU/brkkRDky/L25hbMV82Rlnj8KCp4OJBeFs17mS91kuk2D5Cn5fpTkj7vb94pPB0axJC
g2AsMyHplPVAOBgqyGhkZngShGI7RL0PqFns6nHd/+P95Scib7nljnPYI3YQGRswcP4hXzPVu9Ij
M2R4rRQirJsGCAsQyDUXWLaTig6+j6tH7uaWY3ixBeOhrY/fg0UpgxQWiJFKLj29bOyUVzpSjVYs
0qUHeaIKW0bkbE3V1bZrpYgwjoxyPf4KkW4BLBBXOCOPXPxc4u5NJVRG9VIBoSnv+ksj+PPubQgC
RhXYbMYipfQLnhd1u+rYo8wAUGqhg0qQD385Xy1oGbnoMMVeySxDLe5T4c8lRswcQaslmNtvKFP6
m9UeyrB5OxzrkqY3ul9Kfxd3ok1pLmNXHK2nrcrxvLGCkvPV4WqRKvbmEpUgJwbKJg2DWkGXApu3
zSu622PkqXD6wSBK3Mxt8N+VWCkpadGjX/HbVJdJoe6JgNXQVSy/TJGjNP41UsgBAglLLyvUw98J
tqrjhjPvM355q/hDx8MGgFR7DTUIhRcvTSh6P5FkoqvtqjhYPQN2Kpistt6Rn/dGZonbaZDf2Jd1
3RvI+v2/yG+5N+Qh59f+91rVbeKhqR1mk1w4H14nU0cBxm1JMorzwJa++HutCRLy70ihVY1ll4YU
r11kPyqNiITrgkl5YNnDe0zsCxIgKT9VKE9p3JeFxQrYwaxTBm6tTD21AuBVNOoPFdrqq11q2DeW
luYy6SMRbzEoUsMuc74PmHh/c905rbfp34d2erqZ4AuLOiG0upttiVrIapZ5ZeIGF94Hlq/V3Hnb
3+Zekf1G505ceU/bJwLYB3zgc4EYebWovcRLZHqCW4Hd4JLcur9oov3z+gzPwpeCqlqAJZbMvopw
TCNNBi/LAkyzRPlHhTBKz9X0+Nbdvn1n/M0p7ZJddmtSlIBug9ECIw0kDGkFWID2AIJClmA2Jp68
ib4lP1c9fI21KpAhtTpBlzWiK77kZjMAuxUoIpSpt8gbpzu4aDn5a0U5t9TuTs+uZX3sQgy/eps0
mFhtUCfcxzVBb5u6uxMHAVLFc9XBR7yjpJb9MLEmuoodduv50btCaomCcwRgleKATJNv5PI93VZc
Rl+iI4oHKsk5DbJRBj48HNYA/tZbFG6KrMqnB4/chgTj+wEBJLAW/hFaix7NK8lcKD6v6mrMKaGh
o8nruM1eRODAbuhMLJhkeBanfK5XZJs7iZSV3GwBLMIely8SK5aSVIVVg5T9EAxEE9AyXj+WF5HS
xC+6OkOZz6rs9KgY6DjU5VMTcQxeqJMnac3AwUEEwg5QLDNrxnAZRgEktmQ837s+sHpPp2MtBAYn
pomcBRsj8rqfH+4/+Lq8jMB/MV8DVyVx9vWvTtOcqYXDOxPfLklb5rMCP6E2lw8tMxLezXRFlj7E
Yb7fraxgUqc5vQ8NXTneXPCw9muPYIMlqJ5RMxTfvF+uVK39JpbQuAjfochnr6YxYOcXkbcVdkl1
tY5cSnC4ZABRM+MNY2fB1Zn1E2cqk0aH2ThHLPKVFcTSCLicCzR1NnUq3PH8hqittqX283uxXPP/
kI0kgsvaxAVAew08p72P6gRuWf9E44TC/8PrR39pf5fXb7MHo0AEjyQVKyP7L857NIWK4osQBv+m
+57+hozOctG6w/a8KIM2MoIRisnoC9SQQqmTjUAMoXWd+PtOwIvcVSG8KCBNWavvjh0aeFQlBPsX
ejsiFE6bgCakJzWKyFP87jtw5/Tz0GiRIWmb7kMNuk9CQPQRr1hExxmSNmSRUZGeTqn2QZ81Q0y5
1+VB2NobdHj6yN7ZxffqB6w8fJmOeOn36WyMQgqNvTLOyXDReiDk9ypS0o/xYHi62teX7wD8CKDZ
KbjHBk7RIZKQtvVo9yhrVx4iqB0eieOwsrWeY10bmwSGNOIRWIbgIs8rHAcf/HQj2r4umF7e2xol
w6fB94JrGKqfMeHCrVfw4A2bPZf+RJ4f0to04nHgb+tcahsl9j9zoDAHfzT9Tl0o1ujkENulNxDz
zJqdkp2OFr4jykntgUUlKuYYxRs+to44SL+6/jndTFEVjX4kUVertjE86U7lDiZ1L54PtczV8R1s
ZRA4Np84vBGDPb+4Y28cPVjfpoXSssnSxWjuf4WeTMHLnr9CU11j2c/iq79BVMMYC8DEPuPuL9wp
GY8IpPzZ6f3/id2XYr7sNnsYjEdELjF/nTt13nVdy9QIHCyS1Vn1b86G8JWQGhGZqX4OGlGie5GF
+dLH5+YJhCwta/O7ae5lb213dYm45KTJxVMazal1UUQDN5Oms5XsqWgtQkdd3/Rz9pQ18bYKmHYG
aPLAR9UisG/hSGJaUxpKmdIpI2Na18j5AlLu1L9umIyFvaVhjU5dB9vTbf5F9izGQvp/rriCLT7o
h4hv4Nxl/2Kv4xn9TdHFd5UgryRYaQuC4V0485rk0fKpPGmItLh8bD1RuqyS7BITmku86gRQARoQ
ChFTou6rKEDX7oapndMb7XrTgVynAJ1rkvpaDIXYFUp6dPNkicLF75DnTjoqwbxXKM/PN+eC75bH
fGqEpIlf00lbOAYFeZsFtIPnibGQ+mJR8nP79hkf3V9bHMGWUWB1OJAhfYZH3TmtHHlCSXDL8sk/
0BwccvNyYWnhlOjt1o03zuibhzfIxLPzOGFHnBXol7dTlr+5Wo1RS0KHWTp8Sca+OhhRg82sUwmr
6+gC0P1X71tKGp4JsOTHjJrKTxv+hkTAISRNgWxzBtEpKxRO5MQKBjn9L32Wb10CtQAqNKJZ35+0
V7/aRrSoa2JIAjn3UGDFVthCcgYPJqOhVQ66huCdA38dn4YJEZb4ZF8vod5dIMtFanVhrGeKy6mf
Y0WOwVMQsOcJl/Qm/ygrHfae3s8unkxoX+xYo4gejCfapKUM9GplpjEpLK9cVdIHeLykJ6oe3osh
OvMGohyo5dD0Qfj0ywKJoHNf4IaXu/ud+5Jv/8MrZNxgvUVx2B/v593W4aRxL2usoJ7DmbWWacet
2dqM2JbDnjcfu7NA3zeXcrQ4zJ8CedigACly9+2u8jpd5PpS0srnS7OQ+9ingpRywAygRgTW6TCV
251nxDfpKimYHO6zxga/mmOCy3yIsuJx/StFErKIXLsLc4qIVMXKuqaTsJPryTsWgcycYI6rwTRH
IXV1O+OAxvZsjaay/aU0b9ZBQN7/CF2Uf/0k+8+Qm7zg+wucQqWx0ExRqD1RYe/Za+OyR+0GXDTW
symTHsQycdphhGQymhxXztDkaykALtf8Z+hhpMIxlbkA1LG67htedduAT8ALqFoW5q9WY+iP7pF7
lafkQZ/OmrlZ3al68lM27IrBLkkT59LaEGCxibDT4FSLC86CEsP9l4iU/tSt9+sZIV6FlgAf9a61
ILbEoI2WhcJYJ4ntnZ5DtLrGHZqx0ly/eicWJo6D9On/pGda5tsGhEE5B9wlpSZdpchpX3a+f0zB
7RFWQMvZSDj1UAfL3LxAv8eapTGWoAwYXBaCCPKJLhiIfL0wYDBvnzAUXCtXZDO39x1Fx02bONlM
m72oNb9c31jKCLgEdLaogqTpH5qOr77Yvzv+A57Xahohfva5a6p6lSls4AQ4vRdTwX7+UtLvPcx7
MJaUK1a6meTNAhFbdb+O6PdDx5kZvnDtV3MXqYBGP7EAsyjHTffixkxG3/A/dIGmKCt/6s0ps+fO
02mJjea6umyFhmBflCqt5K9bDZ5F1fktvZ9IdG3mSF8+i7PXvrbJQokiln40LZB0fUIw/PwvqC4j
WHODRbhaLD9XIXP60xIqwiKeGM81N76kC6fxkUfQJoW1oTRHi1lmAkwnhZCD6llCq9C26jvTo2Z3
q3k1aVoQ2N5ycOaHKNccOi8KoU1nOJZd24ywxl6Hp78vT9+F+L+5VTcBTNHotMBTyFMRH11VOu+v
dX9j/gdH8TGIBeK69u81BMPPAbpP2fW/wEiXDs6Jy5tCokutaw18/rjqurBG+nTp8/4d0cdNCZdt
eKAxl/iUR/YbEMsz2IYCadTSgRPk8tcyAUhA8seJzFa17kmlvFnv0Wf3QH1YOeL9MkhHwfmzztRr
7z5oGAjI/F8YuMwvQhrAXCS/u9G9aGui0xgliecEcipeYMJFF42m1Qo63h2tVQnNut5wl8jrN7qL
3R/tc/6btKC71icxEJTeptSo806k5A2a2/2EsfulqZEWFdFGfCt+Gsn+Bf1fuApK/gS0iREM9QL1
5o6CxmXorzk1yQgSn6+Lv44edtD/IeDh+CjNHXo4gjDx5bLs3haa3MmJ7ZuoHvEmDbersdE3cda7
HM225FiadNVvwnZ/4DdXjPTTYH9Ib6ayFExAm2QIJd3fWSGKa6PzFWifIktwHH/5gmCyxTWQ7C+y
rs1/0idoecWBps3IxTbSla/A7OOGWljecbcSAJbY5ismtBWIlzYFDsl7AHNOhoS3a2Sg9WbDAvH4
I0Pdvq8cNq5TLOU1Q4G1V5wxeFsDJ80SwgHYTgpxAVy/dzMk+LIQIp0OMzAravJZPesYNFZhSuby
ytgVgFQGgtFLLVqIWzQle+vWmjK3VxMvrivUu9KhhR6+QKeA17ilWh1RhBmhnn2NU8fE2PAqrosd
9Ozs7lhyLwr9FUL4ZZ8PDe/DB+7mfScFEVtJkMXURffIWB/0Sv1d+iGEgp0g8wtit7eVZlXTuhp2
kWIBwZWRVCRbHYP5Rz8Kk6BpE/3brBGVtWr7dk8S6Y65aEj39ujTGiJXOnKgrW/pdozCr6XNMrzC
Q0A6tVGLAcDDJLuqGsYp3ipd0U+hf+9EYMbAfNYhrWKjNDwKDJWtXflIC+811VpLjynppKGJJ9HV
VSNCJAd75FKnKGxrizosMGRiVCYu56FmiqVbbL40OXEP6vC2WDhO5btye+hIm2yvbHDBVUhjivx6
JYCirLzBGw0LOahIOtxtM86ppEVlfTQeb505OippnJpYQapQ+9+lZaGXDPzDaMOgf/Ywy1yFajUt
qVmANuIJF/4Ud/6x4vHoyzGevs4pbahfkudaiMrDOwnxuwLNTlo+J6/VduBuLz49cZ/M3ZmSnugy
dZcxKVxjq5fYrP3ukhxNaBkJpFMEnKesR2WQ2FQJVEqrgJeQozdHpcoi1wHc5uvYkf2M8Wi0SYt2
cWwv/Ni0USY+hen8+udVOzOpTyiOWCNCspgZB1gfNXu/lkX9axZR2EzhS7yVqhFPKfLtIJFiSb1w
DQzT6s8j8tGZnLaNEqtytspSxyebzBwaMi3hBDZRb85ScbmCZ9VJV9ENxqIvcVal3Rdf9Mu02cp4
lHBnJ81SDelTWqe70Gm4xCFw8oVONuml8PMlR2YbAa9FoW16JdfQ+8TQa5aL7PNiYHofV5zBMLGO
eCTLer910kE1Jgc8FKz7Up58zb37DDMQvOs12EDluiiTzSQJ/JWIrACQUbleg96txdd8YvMefTlW
jufOgKKVJIhuoPb5PQylRO09Vqdts6I+fDPsckVu+sR5ycxmR/uVf1r8/VeXkif9el2kNlhzq1Ee
m60iLRI2of8bScfzaYMFO3s/un8IWSiOhKZcnesQIsFhWgSbLdxNESMhGwP1iQDyMLni9KhxseQ3
wxpdeB4jONOwUSVn7I6aqT4BOujKRqDmCQRHcs2MO96pirxXnScotdy2RR8ZItX3GSxjDjslW4IU
+8kf+d5qRQWBSKldURxQ2+Dtv/gc7EJ2b43kL05ac1zzWxqhEhvM/tYBAEg4JtaHuq/PnNyJyELY
dGCV1BHDjUfrAZXJmQKB9n6LD/EDzLvYCxGd6XFw8iQ567RtqfaeM71OGApIygpm0t68qZYfU8wG
2pINdNTpf9LBVtNq9We31M2zyqZ/IoiDqu1omTFSEZZHcgV2PYN2Kxz/2feeNmolZTLslvVQN76Q
7zavTnCZVn8Nn4MDPaZ4uB6bZFSi1kop8i1f/JU7O0Qm7qW/5vZ2vg4dyyNgvMADG7r/gjTqjWvy
u3hNKuNa1vvObyMI9CmZ/6wNkOlkfjzwROZQMR0LxVriWxPozIKWmkyd44Fw/FJWHLL//8CcEa1f
VhosNwKCZZAz2GhiGStEtG2EDiDZivJp9Pya2VYCD9dG6UYfExOpku+CNgyEoh0EbDThFT9zKOzh
kOhtDIQskp401a336AVydd5YKfLQJ7qVVM5QrOAFad4KeEOyXyosWZkFaXlD29cTVZAfIkVGLWaA
cfjNMqm40OvS7JUbkVVnoXOAwF8mXDIDu21ECk0iGX5SXrwibqdkLoqLxSmi0jPBL0eVp4PmiIHV
7IoqvwUnWWZsLO2sYBsTx+LH55kiatwEbyIr5MP0dfm2vdxPA5pJHSv7V2EWIXbTYCWmAGEssd5+
QnuPBSZDGv2wTJlIN8aWJeovqI/jr8JI5LjKuTGCF47k+FiZeAaL6JMN+/8l0fY4RA6QNkfDq82J
CZJb8t/b6pbIEouIJNBeoQR0nSOEZSBvuVH/MxqvKUSzry2TWY0/3P5wYVvtnXn0605BG/dthpDV
7RsHDE1RT45gwJ040GYV8ig1VtuxToTxxEWfCZG0C+dm/apefweNzQ2mFzyLY7YzcBrq+M+fpVxT
k2YokwpbZqfRHRcAUm8v8+PCoYz6/sVNifti0BeEbwzYGoJAKeq/780XDV1emGeFH9vgR33V1Lw5
9KLDw0d8MYMwBMxGdXwUgAnFJj3e53StfwZZhmOBG9Cqq3Ha/gf1YmU4iGaqpTeNOFVonlDwIWZq
Tr5BZcPruC8uoUWQyh7fXNZn4benEE3wEO8PF9KR8x4WR+seWJswFHi81IqhUcLMATa3kTZIMv54
9/DdziZxB5HGv4FSiUrYGrMP46lJC81GhD5mxOLcFW/eJCf2Quqc5kWMvHUq4am7KsfhawiBWVqo
7eMStmY+4/jUGSVJF9ETSV96M8QGzMYudAz5StyVEzl5+ZIXQBDsz5cVSZNASy44LxRSuAc+0mlz
YaNu4WrT+zzDCXI9ZnmxDd3WD7jdoj3oaFinMxmQP4EiDYtU989ei1tni73p+FGWNn5PQwf6FAPO
+J8X+6MsRgAhvWm3U+deRENH3agj/Kic5fm0BvF1FiPaNpBYQBmiuTNUfokTHwvCo8qdOi1eXGIg
IzaSBB84WIOqgk2r+CuotQDstU5Z7IPd//O8Pdc6p/gRGMjyrcf76M6RDEpqrJmWny7WX5JI2qZ4
uVcgbkxMbwqMLp2Rh955GikhJ/L77fKL+ss1PExDhKbR7wa3/4+tjbqSIZGXCvcnPFJGg0ZCLGfl
jCHJoUCSwkn/+wxipaPOkEemqnvLj8YLojif6+vNNqfBkUiEzBz1Rgwekd4o5PmhTgx/lzX8nNmk
bocI2Fm6A1YOdoOfazSXK7C5kHSJqLrm5NYqaCGdY4kJC+gI4VznhxemA5LJEEfFLXOsty4JVV6A
z+zhHvr9P3+cRukhNwo9ekW5SINGEl8i6NyhPcqppAKOpF0N5hNtcVyY+tCxg/Bb4ujVf/q+g6Jl
MWipe8QfwDnXubm4R5m+zaRtXTmEyEnqBuJh9ugsYAMMkY+PwlkXycw71KDQYXujOmGce4NIBVSz
1Lzu1w0j0KEc6qzxxPIaobA25U6xPcFWKlVfu/fZ1W3SLb1OlODR4y53Aa7IGiGSasN9kOmpqHwS
IOCeE2E2AQ0BtPM7payAGZNv4eTBr8qSBWwiSA+FUbG+BG8U+GPUvFz0TLuLiIghuwebjHcDWY4J
H6//rW4fw0xbIVnaDhxlr5872XBImuWbAWCR4ftPf/9pdfZTJsf5APLSF/t7saszMmxQs+KRE1tu
cpbRmMHGxiaMkZFmawQOa8hvqjbomaxcSBaneIbCNEZeFk1SXbZTNEi36i3Hg3hgaP6i87u1nbrE
bCI+kTgQRC8Y0PY3jeF7Uw9L+TQnb+/aP1FODmjc3dQjbcz5NAdv+Wp6y+hFDwZmZJ3U2CzpUKky
Hs+bnRqYLeyVRm79q1w4nwyklg4PsTR4/+KWiTPB+ktgvw+gDrew64yrIEcH/UkUcXsK7T4pxfHO
c1YjaUB1y5NR7i3upkqcUbgYdAugD2SIuYB6deLS52U5nFUWbsYJRW84+4fmjlPi/RqQEd9Gh1zl
6bdKr5heplaUCcA3iR+59JRhd3GBdPxdMRT0rGhMDcosifto/UMtLpxJ2Usq2JV3B7gfEpx4q86/
GCKziHeGNHrpnTG8fe1bQUgcxzWTVCVFi7ATgqUh5dq1PpW0s7rlAyKA0fY9PxOABfdx0RXaoCvs
GtslYhcyaqDdCjbHMLg2kEG6s/G42T/KNGfDbnDtDALQztH59kjmn2PDIxNUwtQ7Wylp9RnFiCj2
+jhDKGr3VvOVlITjZNbXLym/ZSg7dLfTtzL/bjd11N+UcSc2bWn3wPFhstmOp1Jj9lVMqlbDnNcO
+zRtHXWFivxT7k5kQ9ZZPvo//7opWbi2ARIs9xN8rQ076yGNv6Odhd0V+lGdpGL6DlJPPigYbwm0
6gTxKKfA8M85zDuy0GvkJuk2EHXdwzy2fz10KzF8ufdOwA0cfcFSrgDZYMcjQSQWRq6EpMujQt6n
gygSF64WbrGcy/ztTQ47j0Z+Yv7Zxp+0AmsJ3DplzR4v2H8pxeVj10258v10pZ8ZjS0PR7VQhVzk
OLk2PF/n6mjFgwyngiNBaXj+oGrYW0EmsIBL71CeDMqvSNeYI9BLDJ249xICKbcg6VuJRuUserpK
05WkjX6rPlsuqbwLfKSMt5ZwEg6FKm3tTbvhWZA0zaSHKfg+1F32i0CexT0IL7LPcc5qlAfitnNu
DFlI6jw4wWhEVXTR1xBWgNcKUv6HzlHHN5wgrfHOtFmtJrmu9UNbotgHkU3FvMR5tQDwo7JUXlZ+
NRWFjLkb6WJAuRJ/6ubwPh37nBWTb3hxYgbzJ6XFNRhmGKD3oCXjznpupMan3rl9Vbs28zjDKwDC
UOqYm7H6WyCeGbMhxW8jz+Bmn5gl1iJiuzOaKzGpi+arckEMauufB958RD4DHZecFTyTY5tAFUlv
CUGVl73EJEfefdj825jd4cFoBFiG21RT9ZK0qwrkDKptW53/cZ44JjM5mvBuh8Zxzi+QfFazfOWt
bzmR9q+INV2ay63u+J5lU6pOKxZQ5AVGd6tnKtVYxU9wgqR4VNjg4lpsr0lJbmQhaoVnFl/9AwzR
lPX7pzz7MyhaQu4BCwx7a69CxkUCrEIQp9PuDs36Tz7PXjpsH8Jbx8cqyK8k3VqBym8PXD6xlnGG
Er8NHnqT4cVs3BA924X2hrOHIXusmeM//WUbJxQyklujMIWWsheUN9Mqj1BGhzs+FT+9zshLzHRI
TldVWzLf4gUby5+3hdHEwOc9AADTJJZBk1diBwnVPeZ7ZpT85oUVtNDe/6OwzjqnHDDKAtdBwdXp
c8rN837XKXK5azUhYw/6XLnNzIB2mHiNWAglGdYCkaf5Wt64O8/kuchVvFO0jFeO1UeL7FqAc3Xh
af9sz085izdXUl3Dkw+IaoBzcNbYuVKUooUb1814p+toGM14T7nDfslXewHPX8azfFswoaBp4+d7
KSS9V6itS1NIFKX1SGP0pIYhWbzf5R/U/Rd0Qo5CHz0IBUYIHjnFAVO09gqHE+5w5qgKEGKab48K
ZEOU5PIVfpMKqLHsOCdgfGPkexz7OTZ665BeCkTIHmWwrZpTY7aKUUYm1jPm2JCY0IOIBht9LCwb
+CRBZDQMs0sKx0WKp53b+gQEN4r2DvVqWTPx87HGZLHclYkm8wvDf1kMr8N3whQTmPgTc4TpIqer
Gc8K1n4cNowKkyRNu6qW0lUxKWJfML+lFmDiht6jUVhMNCrD2lkt0WjgSiNzrlY1SufCFg4VI0qm
6DnTYXy++Cd25zCBN/b8xRm00bRF1dB/6NM0L/RReMl6p0IuAtseAZ0PmH1/jwqrWRdGEHvSF1cH
Z5p7d+g0JDt9j1Wf/KNtqKT4Yg6lpoXVC3Ubn0yCN3iel2XpnXr7IuhkvW8vK4jBw7C6wcab9QLG
FGUqWzW8rtbyDZjagUilf7bsJQf/gZpRMwU+VVd2v21GhrnLbQbFc81da7AUirBguKBh2sg8Rr6p
/CQJMHZw7kGC5uGqYVxXHnaZetUWvNDmLdwdcZgFXjxm2oITHP5XEdMeU5vENLzqmZ7nfyRaNJXP
1TWRFotUWu40d2eipRZ4ICrUUPpfEw+9a8T8PRDd8VYUqD1N96UGCxcebU6Woir6JqJyGthqGwfs
wA/L/iixteOMxOUhwRgmyIDILtH9g1UAxfPOUKlWnVCUVYbisgvUzRX3ZtYvn6sBBX0f1DZLa8S9
f15TgaG8Ndzn63A1kcT3FoWw3D9r3aVWM8BJM4UkuMVxuYGY7LZh+iYoXe1B7gji8FC75K8eV3yl
yLu8KIYGejefg4Gk5kRuwTEK79Qys/tYhBtUIpYonmk1DZdZo9SVCzSOTkSNzdi8kJsijZHOZmo1
t0PyFzZ7mFz9P9R/3ZEydDQ94Ugc2Bstc3HPqgJzs22kuYaZooGl3cQs5/oqd9C7K9clyE+Q4cbG
7+IO2odTgfX3tvDi6mCUX4nfjlN0jhLHx+DKFFBu3l3gwokwskalVHuwbv3u8VREXlAVlZpbDs1L
TNG6vFpcuAOoif3+UIrs6WWjjRgIbQ5tSiODOSl55fVWGSANGPnQ/uy+e/x2Yuzv9FBQ6PL43xAN
fLnSXwbhSpd8Zuq7eGhsoriZv4+RJIt1Cn9SJ9tkYj2LqbWwxrJdObfwY2L4jt71mD2RKi+zeCg5
W6CD801gMCUd1p1zXH2shLM2iUj1yqhWLxAG6aIb+LqAdmIW08+llLQSQuB1vUifkdo9smrhnMzq
UXmXRjTGuEschLCXubs5lydggxlkpRN+5kO6F1GTOZFtt1DrQ7wNLiGKzRaXfi5wXl9gv5bUcD3H
vUQYvUiXZWJFuQX8F6MohgiD2luLS7t1s5ajC5wEZ8a97TLKg3BG/MhDZdFKrzqZiZ2pdTC85Rcc
qzy0Oo5a6AV9vL2rgw9VTKWQMXNTFuS3icwdVtpymtV10oiUDzNm52lcJJUTXN1Rh4zqAhpWQbdJ
0S8Ls2+tuKDiddRAK57csCLl7JX3UNcJbqBH5OAaSGAcofG864b9uGLBu/35eVTCy+jPN9RaGmI0
iCQD17nvDeWlb1tc/cNAkuPl/5uMgG9YruQL7qkTBc0C0WVuZMDpELEZi7zBRlT5Pjki4mC7sff0
hJa59J8SpkwjFM8vBQ6V7SCH7oTIGBme+Wm23WxsRxmyx3lmp3rUmoC+qWWIrVYGvONrghsVL/bo
XBYEbHaki/zUdfDSTkHuhbCdXIF4g+DTXcTsSIx02XujOPoEbzL5jHBygosr5h6sqk6tYUcHE27G
iqARO0cQAHbjX0g5AkMTkpQNVnYT/fT6Q+3RPmwOfcy1wHTuusYF/gDULCEAKne5vYFUCT/2XfAX
M22D+9mEZ0g8KLUWQoCz88dE3CvjhZ7hQb37l6bSKUmmZs9wvsyerFQyz7Q8372tnCbgkJV1jm+C
OTbmyBO1qKyQTXKtWVLMj5RI0znSRCjEbuE+stap6ityILCxG4yPooHmmR3qAR9Go0HjcQJFiAnT
rV9ur08QiDHHj2Q/Q9VUH5fosPp2K/qP9jbcqQuNX6rP0gpsOJV3tQHT6ZkSkY609tALZW2LS+LJ
os5HO7ZKUksdh1rHNGq6zfViU455C9bkT4dSg0e6RXQxs77ESNjraEOwWbWBiPc5sFf6mAPbo7Q4
wFx8arCZWLd7W4at+dOeMUMHpFxbAZ66O0vXPYqgMlDS/b5ERmqgAncc8cuZuipfEr7XOCqcogjX
BYCVZxYcyXctYoV2vZ8wdUajW5aGJBEVHX8IPAJyrCD4BNl9pJ7tFYo5LF7z0vat6C8p3h/3EmMc
b697Bv9er1TOrtucy79UnmEvog3VRgFD8jBxlgO2VRIHs+H1Yr4renH3szTUBRMIVGEzLsYk3Sld
dp61KeiC3Vv4daehefRhqGglcB4zn0Gl/d6ebJJWQ+Wb+NyRC/4S+xJM2mjoJwnU/muAWIloJt5S
HJu7ZMPq3Tk1HKR2hi4cfViV3DGg8VumMa588kXvtzlqNrsOBcKVWEr5bPIVFbaigX4rtYFu0l4j
ITnyi7kL98RhxBPSsgSJ0bacf/HfYBCPTASR8fwPisB85YkviMjJ6jraWTgeozQh+Fpyiqoxlx7Y
FrNiPaTKHWDa8Sr0p4+z1phhMWmXpTyKR9dsQAkHg3RT8Hb4P1sEwHdbXB16SpwpdromvpRI41Ue
zB9jAwNGavuCSUARhNMf/L8KFKKyxRrv/B4w3Ht34N7yZMGSAOdhbJxHi1B76W/v6lthQAgfRxCI
bwzzLEuhG+BUJeQankxfMoDVHhQue3QJS4ft8djzx/8oahaih8lpX1QLSjwr7G8VHG8OteBzxTHe
rsx4b1sLIr1VZjiZ5JfUoTuc75cIoLNe7zQr+2jOLkXXx4j3h9wcwg1csXOrqozZ3kc89oBJdL3h
uKJj1ph9scF2zNYK30VeThLPyofLrUJSY34Rpfcc/BwXPwDNO+2oe3nK6dvUjI7JWDTjh8vAZtfB
y9pSYal2ob40PFpf/+Jj5000SV2xohii375VaAwMhKbiKhAw3ykuRP1Ra7GvtXHNHGRvS0ZrvzGs
G/9dFZOJE8EZf9qGqqNbmoRm0pg6Ug2Gkwjbkc7yZ4aKUG1LsAc7zagD1P6Qr8eu7C8AKn4Hkbhf
z/ZoA6VWYecQ4LqBofj8hFfjvzpSR0di+5kEm7JU7zwZW3hJYUhEeRMK6ZYDiDBTvkDTWB1EqGpR
lMXzFxHqno5CIYXHFA/87mwIi+pdYfi6hbQcMR8uxiBDEP9JoZdDnvWWvd1U0/5RXXH2Xlytqjr0
RtvuikPHdPxcZ0CPe2anDUWd1SBGi6HyD9kd5Aot5gyj+Fou/CeQm5tcLgwxiXHBop1LeIqwzrCl
87+4XfUmw9Odp4it6WND1M+msC42FjhMS6jpUsEChUp/+OMOA2ZFjzgRbmBUYSUJ4iRtilD7e797
UgmIWPHZ2zDTObFW+RxzgNjp/LQIdnvxlKvgqAaleeWVGK1an9PNNflMTE3kBqNCLhSlYvuQ745F
rlxx5snqjEn5BH4/x06Yd4oA2oQr99HWpLA5psHaA6ALu7rfoIdQIdc764nry9YqgLJ9tYT1CBeN
4XxnqoAzBPTa3y5zxazI6I9H0NfpWBFdtbmnXx8czrqvPr+v/i633cHIt77IObwJb2GluYEv5Dht
je8H2ipNU0kyhalOavRLkNGDc0HDOlZqB9PYFWwr4+NiE1PX5Fji37NDeZ3YBeVt+S96h8II4faq
KBCfEeZZChEoLCPwC1BgxFX8sMPvCqJI5rNAI/Nbjbabqp6CHT7jntai+qNoifOXWm2iutclWAlv
+2hOIRB867sFzwrEr0kDbC+IX2sTq6AgVUN6n24hX+8XJWEIya7DtwyvlCtGdzfmp7t7PG/bYccw
fgs6LIF/qe0F3VmBh7jNTK1peRvFBP5ARs7bX4coUpr1KX0kDixPXUPeRuzsYVTe/x98QHnlNFq3
O+GVxcHq0e8ZXOWzjZhvJaQwzimiLUQIEN+FoP2gIvBGFHgNxTj25H2fDrpJNxQoO0Vf9nydX3Sy
TLGpiLUEmc+fMhVL3m6nmpE8cAwW/Bf9VXOdaqIxogUcbq6wATlSx4conyH+uiWvYiQn8vS2HMNv
XMGaa8UO8O2CA7dbmbhcHyoEsviLVwgqpizIlqYhynzotTV22F0Nup57zHl0IfFMEWn5I3UqdrsF
CsrWmUKwe9pPK5H7C4XOVpwMSCbVhz6gPIywzMUJsqjeq/RrvzJB/6xIGLdQ3oXGys2a/VIm2u9n
Z0i1CVC03KJ8NzVirkhCoyDv766XdY1su4FJYtnE8KyMwO2DokdH9fSkbJkf3biJhk1HQqc16m48
E+UjkmpBp0nrQ4v7zD/UmdjuttI5/MMQhMijPR8E0w/tlUO8mpUTWbn6i0QIs+YL03oXA85wT2wc
akSRnvQxUTDts0p2ocfbaiWNE77knWVzqCW9qgZbtzCe+ZSmdOITJ39P2qw4LkyCMnJgYZ2sKexI
r/+Pg/RLBjIppyECVhJ5eQKFezJ0v5k9t10PZMQE0AtFyFANQhNzX/nuvIjdqhjMu3s+p/a2d1Zd
OrBq4K1CQSnmxfzNbfHC6sg1nF5TpmCrbh9BCIfF9NO/5hn88wdoQrNsHPG+PY6afpWGn1fF5T2j
ANONrsAptBp7/3QEbszdur/pN4PRP5P8EaWca8kC7j6hHnRKhBWIbwQtjj55r6pIp9ZFiLrBE4uD
A/1MlRdnE9w/i7my5vFZTfd7la6SWv82/ubGkWdNfJiPnUUWWyyX4BwczGwG7hxdGUlLpDW2lG1A
z0g8TWYXvc1qJekVh4c9W5Wz6+yZ1rDR6gt3bMK5ajC5QHJywYYA83LGU7jmR311d2XW3DaW5Vg0
9XZNbQV8+t6q5SIbwtvGG+02izEnSK/0hsnr5UJDKQo2ME0mPMICs6dV3nt/4wltw2CfLr5n+kQE
Hv2bZoaXn2Glev2G4yyhOR+HYSC1CO51Gnb/OqteTgZaCyPZJf5clkZm2mLkGdzCzGNYtDjbrgQs
8wtmlOwKhgK5w/0UmgIAfLFgTH/G+Cec07agopjVOD4I2TzsO27udhfzP9vG+E9eLv62HwTWL6Ou
6CVpjn2XKL/A82lsEyWwYklI/tdD84R4Oxr8UXidUby44KA29VeBaCyYStHANu3dDbwFGZ8P21bI
PJM2tLRg5q++gE7u2U7saatYpZCEpa4m3mCGGfoWt9paD+L6xH8Dgw+UYE95kD8S1LxY2JMxXTzw
SqTMHt6UPNcRlGwpykkUc1W2GtH9UDfwqrDAeOKrI0okn4UaQt9fIAz/s1Bw40YZHoiXyygs+IU7
F+JHWrEaIDGSHVkzRjS08rkysboO8FUhaicZSU1dCeIHeVX3uVi9hPHkM5QfNDxKHya4N1Jz/Dby
WbEnW/iDVzTr/GOoSs5gEHyTaeQSDaRwEh+PvVXJhmrtBroJOruP2k43SpomulKpkYmWYyhhpC8L
kDb8k0JtBJ6nDGq5lwvnPM708TxIRndmSABgbc98FM1Gi115hjmwEfGZT4Z7QbKJ+rmeCXdKkCPg
5g1CPy0EZUhmFq8PTtwU0FyzLvscP4ZTT+y0Ttwa+i4pmNZMH2dcwQBRusksDrO5sUnryL2Hl3It
G9Fy4Gz7D/eydCxv36K+UhCQzWIint/38/CdxCfJYrss1DzYCkWhLD9lkzej7BzatUKNLPqwuMz5
K/1K+s3bVUNTiLC5+4fw665fEpo98r5++fy51GKlHTpasRDnW5gIZNWkgoKIdwwbIFNuYvKS3X/Z
iF1dm7gzomJdsTLA4wtAegUpOtxaA3BZXQtdE2G51YOgDmhgPqvpgxpfTw8fHUzrcugVepQi5g4z
Ej4t49/Y0VKwxUtjvYi3jMH8m8KGUHkB1N6tVEJhJtK95GUTgQshTRYkiXUNP8VflqTdk9dR5KXG
3UvISeA8BhnLoLVdUYqV1AkkhEnu0rBrQ0ruXIgHEmyhY8VNnS/XEFy/KOODg45tbtCshnI5roD2
yIagaHW7dXHtcBzlMjraiEYOGEffQajNJlIHIDvv/DoVYqW+MR2epsqDJJuD6fKmTBqHQvcoP7Ib
CoNfkcs04Dx3UifQkZIe+G1NGj8nEvforRWpRCdhBtxiAY52xoRyNzNby2fvH23YsdEoTUqiHm7/
/5NkYt1v7PQ3SUx70eAJt4/VGZ61NKWr8oLbQcEF5yr4WkZE4cjrLyYjfyeR52F0ebDx8Gf4mpO2
M0txzFBHf5Nsery2BEiaMjiqULzvcR6TWDJ0yDHpKQM2QQzEwO5OrJZBdJ14+cA2JVmDVdom4/vd
hPPcbrJJbsji+BgyzDW9I2fmL0jTylK8fjK92Jv0rHjqOxkD5K8KvelIEmNP0YY0jgiCm8W7Pg17
8dPmtKWckIv42H2zd7a7xwR93D+uH1c0srj7kpUXRHGQrW88oW4t2g/FPbDzjPFQ/ve4koYL87R/
CB1AS64/9+TQYvB6iIxJdeuVrSuA0tc2VEfJVHYBfSBNU+lBVYOn+MkQmJU+pCvzBWFqhfCNTgG4
2S8Hjh86KGcAe6I/H15Am9Z+N+343WEzMlO75SdTi1mVoFptASPe513NyK5HkUlF9nHkIBcFkjFy
XTqovtMu/zfjhDnrgGLR7z1Alfw1J1BbRVJA5LEdQhzMKh7Cxx/B+3qRHpPcJZaaRIsyexZ+JQWu
hTexq7jfoPjHr/PtY6NRXthHXHldIWi8OwAUJgcsZO/w6UxNSI6irVvFPgoF9ACSQ7dNlgJQCrtf
hHINHiqUgkCq5CSExXxC7GlaC8taQFKbMEqns3RYPipAMHctlIaOv/xfDdskWvyOQYw8bptwfSFA
foTPUctPE45y/9qAQw+M67LyTKWh0SDywNT1/2uwmVcjwJmtihNIPkOhdpXQ1lbU9+VPTL84qdHL
czS2ngVW4jnzOT37Ngq4w6yi70Vt3J2lvwWoWk0Uv5Sew5ccXvAbE8Vn8ZgihEUU2AbWo7fa+bUl
l2VFlnUwS+e0MccmOS+y0JLFRM+jSJY6Psl5J6yq1ZmXBVAII+Wi8aEzdSyYbk6ayVEgQILUpqtA
sex0A+6uIA0zBGJmkIIVF9HWeSHIKCuNzmwaHHaAY3EhxO54JBy2OQyZf4FTPghWdSBUb+pfa3rs
hTRHjCaYaxvu+9a0Pc6r63gBarktPawoHWsCRYElG9oFBzix31haLBPKpxpkZPKAUvsfzCsP63Ya
W+gHH9AOPUrBnjYzQZjcKdd+7Ra7wJhb3T5IKnwS/9eETS+YHcq5O6P5g75oqWQBKdJEcYPotmss
eGQO7S7vpVQ+EhPI5EDEgO3fnyns3V/6Cm08k/YmGNchbd/idwSvbSulGEH58sWukdTEqmBHaPrV
N8docAq1LNqOr6B9wtWgA+iPCokU7odI3gp/zzTwYpKiabV8Y/AyaQb/KGoO3nkQatsWWb/mhc2Q
+fRjqIBMEDvJvxNjiv2a8j3xwWCeOUOeB3ILLx2VibCqaJk++T5XfPLbCXOyUisjgQoBCs56zzNw
ZzkO5j0MFQUaBJrkPSPwNe8Q1+fRs6Wu96Vurz09FiAb/wM2qWb58IqXK+mHeA3jDSWZoZ5tWqb/
iEUgwd01YWaeQStiwXtytXuOcyfe3Q6NT9yfBlX3wwJpQLkZ5FtWb8kgHQSy8oBTkG++6YTQB/sG
jhF0ys+GcaiHGgQLOtNLNXfDjKnPID//bBfs1NmJLFgMfF4vaNxnapQ1uB8YJZx5QgmBwKgnZ6/Y
hvi/5FSYlN+SDk05KTYe5MDTEZBcd6Q1ZewXL351J+fx3R4EtBNU+E1pa9y00bdEOEFcGmO66+Pk
tmAT2AZobf/K+QfS5oHrwYR6X0Id+6sn8HM3L09YP5q3iGpVPrdB1wu7JDwTiy6S1E/GCKli5Owo
pTLPWbUb8pT7BceoT+ukQLXFxmbxItHar34paNXXJU1dFbVXMAd5RIz1bmMFvShmr7DFnxUEswr8
/BA92zYxSZvEMbeApYzbxegVDzD2Hqp/i5DN+Yf0igMWMukZjW8JzJALmujSfdzcHPM5vF6IyHUQ
NgLOAfjqEEVOk7e1oZ4kQKJ/7vyvkqHTuWf8PT+HoGYG51EA6KUyUkwIjyXI4hToqN1aGdJIf+M8
EqCm2tM5ty7WoD1bOQdszd1MQZgZ6M5iEYbIiREAaHBG2q4Pu/0Uyhbwls2N+Sjnl109xX3dDK28
Kzpe0rhQIOKdxuj90JK6nK8t9KqunG0FkkIQs7s+iArbUlr6BzIhRZyTw0wzCDS5f8xt1MWXmxtp
fbhLPaEeaXta0nxuJeIf+IagntDHwKJO00Sb/5CUJzAml3hPLfMis+D3CwduSgj7htsjuHV2kxrh
aZ7FjzKFtkXfqu7R9joX45jk72N0HY/H4c2Rh/44qjWKWh4ny2s8geeFybq9TwdfC7p5cCWEANsa
e/UUO58DKHH2voUHbXv91VHZkMxL+PrVp4M7A5m9WAEfh4/m28C9nInW9EjVTCNXPBCulRpKS5hy
cXWk5j9Gj29L0Wo1k3UWOUlZkZQwVo7jADBd3kjfRnUp2nht4WpVrCZyVlU6gJWrfPD2/aHx6N+U
Az11N+MLpdRoUTOP1Ac1cK161eDmH0mxxs13DEZRfgIyI/eZ9wzuv6PqtULj1XIUH9dU+SVPJ7Fs
2KpTiKPmlOo7yunyVuRX6YhELs9tORYSN6gYvF1Us/KuQGjuHRvJ5dg/Mf/8H0i60OvlviLh77Dz
74NnSwSBXL5IUtfkqblwrYWyj2q09Pla7XHd2Ks4IeHEqSlzUBlPSmH67p5GbykwXALDWuZGcXGm
O7zFveCF8mpoxhm0tW91r36dComkztZxuIvlb1eKWav4OFuYYyY9PNbrvUrIP/WBcKhRzFRYlDm4
fuQc4Yn7rPwQKmD2dXg51hgQS3As7wxnPqGDyqEV1+5ufKs5cySaCpsMbUtKeqTOIjhtMaZwEcVh
kZ95lRlssGtja67WTCjaX6o5pNKosjMqL+bUSyQh7WFnnxZi14GLwDAbgh6e6uHoMMfg56JGiwyK
flAg1Q58aikRl1KDSuCBg5BhS0c5bCQ+yUzYDABt95Wkq8KKDusZnrSVGW9l2OAR39uADzc4kIy1
DBvTvdy9KevHF97rhHG98lEc9bSM3dQHTS2q4oD7YrUWAJtFcW5TlRcU7xdsnQckWqLvKZ0q+pAZ
p6EDGNFfOB3OZwJnrtPdRsIoHfysBaeVcYmxRl/eaU5Siz6psFsLr8ptWl7DiPyGvEAzUARW+/6U
lxeP1ntetTJG7pdKWuOa4Qpn0DvttSnIkGD3LU1CrgOLuEYlmKr+XiAHRVEg6yLkFSL420uzbNG1
EdYuSRZRLBSE68TnawFFAPlQFa/n1t/rrCLE3SnpzfsPb/MgbGfLcmucLrHye8HIYXP8EV+VnQ5b
PGdhwwKqszNzsJa1E8UpvZ0Oxw0xwJ3zhakvf738AUahL62DvgJbO8dMIbghfwqcd/Xhg3ebjzfb
oWywgb6JP0P9fo/Wnb/gImVvlD/bFEXl8m89HvN+XcPmgz4GwBAPGg3NEGyqoKCav5j/UVuYgXG0
JT8ENQ30VOQna6k1WYLC5BiHIll6NmknYxoXNCRB0byFGzIPIQd0WlVooWJnRbSXbWmnpQi5gUTb
yuZQFT62VdV0JAJODM0zprfzxAoB5vL3BrK9eaTP1K23Ti6LGWKw5ksD/rowucPf+ShfqBDqlbtB
+fzpGNafZHvH34UqupH0zIiz7m8Avn8eTSUcVdTXXyFas9KjS4vxZqWRmy34+fkMYZJEe9xHC067
ZMT1irevrH4n/j0VKAsKkkPyLh8t6pICXT08NE1XeI/BrphgqsGaCYDvUc2sB67A6e4ZlBJts5rI
0YE+DFLRAU1ed5Wi0Ue0qllDoxF1SbbbwXV9P75yriLeKT75Flq0IvC7YcmW/1xJNdQCzgNvxZSZ
HMDC4jZ8eAWLpkkGP97j4PhgxGWAtejtSsKDXUej/plMhXchjeYYn13hv14Wpx6ORZOVqLbT1oDv
McyEP4ZNra07cz0QP+YeLQGpGcNvJ290Rf2WBIt8ci37bIOiz+RBK8pDk7R7H0IT9K4WyPcIgbW7
wnDhpblxwrZXF2evm+ho/MZnEemA0glIx1cD9Inzcw0rj6FEtC81Os+E3FoxHGkvKdlOU6fL4nsK
sAcyso3wPNwK6rJBVf/IoOtp5v9KB/O8SqtGSpFzU4KXAU5jSTNV9ocR0jYqGwuk4a0PTBIyrXbu
qzW6x+HwTuJVhXDSqDewWYlh1WivbxFiV79u0udysq2Ty05R6mJwwvFgIaGXnXNvL54V6TX8ENBb
AKtiUBSuelUQDZgZ7pzv/Gp/BEBH6GvlWM6J9/uwxL4hTtwJ5yuKkWB5o3uASxKd5Bogv2DRB8G8
kkVb4ge5KujJU5eI/lQdasG+N9kR9/d0jRHq3P5YPJ63xkBxjNpyOJzktIh8GhiLbdOB2Cs92EPE
JET7Ha9WNt6icTuSAUfB66r3GA0s466nYoptQ6KOXjCK8JUsN4qj+fFuAlLvghRhnpqF6zi5SoH4
SLVp9/i5PW6RNYj8X4zidQNwZcD4RMtf2kMq8MJNgz93MOCbhZaDB9uIsFq8B3bnJNjshY/nVato
rNSW6HvVsRcT1Z1owSICcJycKXvNlFblw4A4v+QHRl1E6KnaCoefWLkTJum7vPDV/WwyHfk2pWOo
B5PSNe7GawlqNAjxrNowK+pnmcLoNwwfgeIcfE++XXMXyeAzwXpkdYe8Ob6kI/8oS7EcyHqp4oxn
AbFUkk79FZSVkpS5pywG/HcXanUHN/Az0MOtwChlzvKJLX8u715+oQyQWdyw42V545qz5GIY3/aY
sketTvfWHRpBAINHCb12Dd2i1nfqPpiFFCc2SQ2amH/vKNhfoxY/8IG+EvvQRWZydNz1s1bfGV+7
ht93VB5yg+VauBY9iCP/v04wXkMvhKl0VJMCTTbTDtlyti576Ah5jI0UPuoS6qTBlQ9UX4b0gjX1
N/MWOV44kBQfEAw12K5KFfOZv3xYB4yfgmoUcoVR3VBuKQ14nMe2CDstmjATR5I0wdDPIod3BYx1
yWLSUX7ggxfdh7mECUm+kNKC4Mx8IXeb981QrYGcgTSPcX71zUiC5iNHdf/kljzC0SadLePxJBTW
qLEIbx49SNrQAwMqf7Zi03+BkiUbuw0uj2zBwfd3sbv6r8bNrsKwDH8A4pi5ocn6CpFKGOYvwb1U
qzFYbi47yamYbFBtkhLEs7S4eY0cySSOBRUuG1xzwcyhuqqomULDZCN+XdtOZ4UDJhJg8DWeHK4L
+wQjSgRGPVGvpIDtNkFz/apGGOdTUER/Iy6rWBzxpyFpEGVQibFaBH52h0Hn2kzcz8loc+o4lbWm
rKPB77CnP44NvyUqomHvcsEDRrL+Hf3Sj0F3EZPsRvaMLG9wO4qXMxHKRfl6248SEW4GjUezQwmC
udMT5gRxO0myTCwwIKOhDnxwTkNLvQZ/l+IASSclset7NA7eXGuCqf/CY1Z/ifsQJlO5wzrBPzNm
vIkn2F60chR9lBSnzeZlTFrAqexqMxix7QNd2Te/y5xYRgVthT+9ITbJiluUXqZK2wprMG/Flr4H
tXxdyqj9aAT26AGoz4DDd8f3xj10ISl0QHUy6aIlOtUmtUffxYetUpvrF2mHYArYXIbcrt8gIFxL
wXT210qbTc9GlHiFWbSpf9xcT/mLjtlhUL02i3qzoKLv+ypGn1MwG8y74nVY3YuBdujpL3EqcgXo
OMEEi2mNNULSRWp8LgNSuDm/ku+vEVKcD+ewiC6UHGcz/oc7W7sC9wmIEy+mGXEbheskmusMPg+l
KDclZabsy6RIg5KpplHMGsUYbXgpYw9EqFWQP9aKSbMcVIO8E7AGQtlBNMrFKnqEBTqUNZhS+kKD
TBc17a+RTyQPnFM52NQQt5Ay+17y6KaxNsyQ4+68siNev8AESsimKOeCvE/uxFPBvOVntykGS8DU
mSJlINJzwkhVAmOGvg4Rlvcq41XA/gfzoBn8uvHXM/ZI/XDqmJuSvwzelDRJxGy+mJXF6Nb0uvYN
sMl6E3Uox2IFyKPQ95NQJ4KQtQmc6P6LBBmOHn7F9V7LjQvTATreNZgqGZ71HxmOpYavFLIkCiWe
ZO3+S/i3iUJTNbE87fsnk1hgGxiJ4obwcOGFOphhwu6P4C2rvanJuJ1qmvUvGwrHbi9pno8heCDS
Ai3IpS9PMB6yH3rl3LiOezlAPOVwjoe7s98yhW/EXvaMT1qJD1JMsdo1gY6wmiN57ab8+zH2bsKp
s65DlOFCcQ9ungjncdGxXPCyj3V2KCaipr6Vw0DC/1K2QOUHKvgi7a3wmn9Omg0pf39c/snY5zt5
19Rlxb7CJ8qOp0qszbk1BgqE0XNfia/pIe8X4U80JJO1OCPngk6iXIirP2+6ZFQ2BENBKAPiqVbq
ZEa9pUd2VR7BzKtB5nKz1zOtlqQ6sQGsJx+fCV7U1Tn+kfzK+21CBFoy1xVLoer5/TVzZ30d88Dn
oDQTbUbrGA5TfgSHWeC8Ww6AQPGlXUSwH3pYxUAO2az1lmdxp9d+eQa4F+GURU8o2nEqT6sMjfgN
CCSWrcH1aa8kxJw6oDKzYjWsaNnSxCn5uvmjXxkXW0i7JSZukvmp/HRrJLMq2yBRNg1Lf4Nj9Fda
t3YmxjBXrHBsoqkvaF+XgtBo1/Pn0DuGKTFqnGbraW+v/2bFb129sU7KLp7x9DeKDuYwl63zncLn
7nQ7tTnc55Jz/5Tj23dQO8CnS6JQbrx1zBKIvI5+2HB8E23m1N9echro9pIJE7CSuobzVDvfpAfv
vXFVCsDCO4X6RIulo9cjaGbBJrsk6vSXAcPFmB8S3dUPi+pCBdXCVbB2abf0LS+MK+8Xc9lEMVnO
uprtC/BTpDL1VsI83Z/6xFIjozt/CdyavhbB0fkbbBWAtcQ4BnPseyvc/nmNggfICtJQxI9XjhMJ
T5XV1U/OAo9HaO8cf72LllAJdCZMxU0IcfFarRedIt3TVE/c3nUI6K0TTkrXfwEaYHcYrDKPf+Cl
XweJUB2ubEuL4aJtpdXp63ZGqGQSYAiPNJPJeI+FobYIaiRUmJY/tnTYgMzWYHu6l/+I2rU+QHFl
pQJxpHBKl61Y56lErcgUhJZfkmyO4J8IdbXOfbzHs8rfYeHOy0Xa7dDEe4IClTbm1f6PEitf4VIb
WeYU4gdZ8TzrTL8puIigAu9I2+1QKQs6dDNUI6yXNUG05RAv33MIlBZNK4q7/zfAjvH+0bWR5wYO
x7W6GT08ofNlsaSp35wzKnh4knYtD93wQJQxItP4PlLxjwyMsCZsP7K/IIGYuiwyOvI/NTWaDAqE
3YtyZu768RHbx2J0OGaZ6SZ303Nb6BEiBfJe0X9kdIKBU1OUTIyrK26/DLGyCGgPDdeSpvothdLy
2ImmA9ZmBd+Pz7hWsAgy4bd+0lBf0JgzO0JTZrd3XxwVpqYO3wng21JOjsACQBRdsnmM5AGe6ave
N9Pq6fQrDxujNCRZq7b8XNjpzLi6B+qm9+cJ3r8/GCdlJl1xVY0c0eEv8f4D6MAwCZBRVPCWg4Q2
DcTbkGD7EhYcpF+lFgD2scMIndbpOlSvc1rANJk0uh158Apomo1iZM4WkFHcUajLhB6WvLJ4GT9L
u5obtKtBrI9mI3fAFViT2vOX81Nhwo8Uu4JE+oFA9RxVPW1J8gGv8PTssJVzLHdCO0vQz67yvJ4G
eDo4p59bLXijDMkoa99arr626luQ1sjt4iOBmRArkyG2nYlIeHFffLaqiyCixspjc/ABLHIRCKj+
UUBB33STls4W6Fg9j4H0DZBVc9hx7HEg6CQvkXXOQg/S6JFJJHp3HcEiQrOWxOfR/XTWTaWjn5EB
ftkxzRk/Nos0H1gH221k4Zj0zlngaqw1lbgRsJVdNEbfyzkeKJ1zwV6bK4H2coDxhAxhWlxBYL0L
U/fXEXBqKLtFwBgiiuH2Liz0GZErSSleL+7H+yOLQKo2Jo5v/goDvOZkYQMQPAUMWZqxdDdQuplN
LIk4Zks0pXI9GCwtJJ6tKRxWbvGI5yWSFC724B5eVn3T0RTZ7zq8iyDkf0S4JLh4SU5KUrcfmYKe
omJZeNzsJX1udGFvQnEn+I2PwnlMfRsJ3oNlfBIkEHeE3VTM9YJrPivjMr7s0AB6f0f9SKZ/IKb3
HPYs7ZXtHPgPl0sR7i1EXiULD8003MK+fdfoLr5OIGOXYDmPMKMZ3X6zUHQFIAqqJceWOzDYcJEm
14QiFHm7g8OmzLreoooucCHG0guEaP1CMtVO7Uu3S1BpD1jEpDxw4XhXEpDGQNXSX54cqZg0Y3UM
Lb00qJ8pXLlxsk80eQCCslYQC+ZbMkAKAh4dvxuCDFapmUVaEN76UEh4E8fRiJiU71ZrV0Ol7iIM
m0N1nlcm7pQjcXYm9MIvF2SR5ilDygP+aoY9X5srbGriugw3I0vdSwsGlfq4RjNvf0KgXtk2XhHr
vSPY+SxZlnMcqYZ7+MolElpdXo3+y6wFY4sbsjWS/pksNnIBxF+Nzh9RPPYR6GFk1Bf/1sgn8RA6
aefIiPJjPnVLPSotC/O7VEXEcXqDuQBz0PSEjAVjA2gUT30Ds5Xr6jzJ/rBuTTQ7vBWB25kQnwg5
v1HEbKXZgSpX+HSTpyqeOuWf0opDtQKzcP43jW+/iIB5H+ReF3KJC7V6dvzGuap2y4VMnikWu+72
mxk5QjZmtwk4Rkxle091Eo6Qg2bY6MUPj0kSGQj+GhfgZcL01gJXBBInBORLBmPf56RzfKbG4vso
KU9tXHQDgYSWBKK2tsGHcD4jm4SX5nwH6mBdNMlG1gZ65o8aKFh1xTCXsinTutnarYpgGYH0Djxt
e+Oksv+Yh5ZPpbf055GF74j1hKz30oYg/2LBAHQdzrAewVaDRnA70bwApZQ9OPtwWfG7eFzTNPEV
+SBcvUgCVhB6jo/zX8s5ktcYRPv4pEuGG6+z2UaaCzF81Ug6loq2Y++txTVaX8hhDWI+TKjJrrUZ
4dko1RqmVQ6W1jIgG7qfL9gnh01jthYqzInlE1ace2X0+WGrScoup2HSN4VlJslWJwO6qboBxIF7
/3PGpp4VTQNBN4UTQTJMDqGNoXrZKPhIRP7bZgEA/lmvOcDvneu0EeFeNKQU+12kDAxRHqKC8/nT
XnQv5YAHxKLBg3jvYSNpcc6A1tLfYx1QtV7/YAisJzRujnVbNeFU3crYMe/w9x5o7rYAsh7oXOI1
qRA1GpDiheizHcDwPEPjcniz9/Cw8WhlP3JUVcb0C/aI9my+6yj8vbCxkOyUd7Ovu5rrdBHG0e3D
DHhNh3mo1s7re/+FNVA2TksrMTFmJCsG0tQhijpoRLeO3rZWM+RCGgV0jBRFnMKuWHC2vlMh/zrc
rjwCjKFzHq5e8DsTO66CROQX96d85eBM2/qUk2q5YLsF+bizwadHYSHUsHHdYh3yOinG5jXJtWoo
M4iyVGEiE/A/vlNJLB7SXaGWEuDgxpDyHh5rlEqRmUcOBbV/AEBPBEVYeEYb6DBj3U92VZQBhp/p
CkxhRdSK8oXW3dHpSyIIXLWYGOgYpm69NDySrmSVKGbrv78ryRNlPwPxX0zBRvgKrGQe234hepoH
IWioQeJVT31zka6YIYIHD8pjOeCKPlPicOFqayIYAc1P+KbktlLa7M1t32oxoBj06AyJhAG4/jQy
yzeHdal9LZ390Xtbgxi70+3mwB/fUfSoDn7TIRlTolGxDh0sWqmB9+Nh9AMm+5T7er6gHm3cUpsU
ZfC3C83j8uHHqTSz0DPggMn1JjCAWw+Pr5boHnj/eYZBnLKAwTtvL45w+8vd8428V51Ok8ThbBNg
fq/WNSH8qigcLE0EcCHZYCoT1raqGu1dlUbTjatB4lhcN3xvX7vvGF77+QqCPMfG21PO6I0vxjLu
e+XYfUV59nce38153q/dWrHyRkPVu8orhTpjNcSWVa7WLenbWEV7KqJvQZT6aH8U4ZA8fY/UeFEQ
cqYEr4AMbFC2LZTMoUeBVP3liCeH0i93IS7DqsPRT+DBJd+yq0AicxBuhiXbeYWJ9YS91mhP73o5
eNIW+Ia3P7BPHESed5+515GWMoP1EHLz0ncfvToGsZlDz3XkmEEK2IV+guQgoQhdqDnKLZvNnk14
wr99UIP0M+yxXplAY4BJoIv9SJwSaISoswzZawMrWdv1TE44dTvaX1HkEkIGJCLgsAUplqun/m/k
0t2rYaFfMUdHsn8l2nFGePaXDbFrjuB2ZXRHwSOSNOYAqDk5ZVJlvDSvEWOi9O4SyIX0Q6ECl9s5
O8Q72zxNcaD86Ut9IXw8/8MZMeia90jdQDZRpLXc9nhL/b8YN9daRF2o0+ufxEmEAxWzN7Xcv/7m
ENdYcSqRfLQSmWJwVLOfc12HPuEuiAieq6XOucHuPgl2DvPW9h29eLZllb4qQ6dmcVaH5OUdQiUO
lonkS3ejvlpe1g0AtIKf60qU+Rvbbv3V+Yaf0uaW2WJ65wshLdmFR5iSNiBZ+tpWX+bfEkwNXWWy
eq5YNCXH2JCAFTVLTzzMolhblbC4M8goNl7SFGZ67/gOT9Rsu3UqIo1+lTVPRThnjKBqgdLgonc0
rQulA0gXZLqf6p9YW8UxDijmQNuq6wDCOLV+39uSOxIpLOCXsY2U5+G95TWOCs13NUCXABe7J7LW
1BtXGHbRszfhn7YILwCeW0RJWv12tTjhGNYTsZqdJ7lsTI/CkWYPrWKM2XahxOTJOQzTSzkF8b5n
um2jnPoM+aOcPkQepnQLyZIKSg9JK/BkgB+846fkiabVI8JLy+Ty/kr4bF6j1uPUnp1lxVekfbg5
XaWq6vpgsmQ0o2qahaho00L5IohUD6+55DBZ2TcYeJ8kTEoawbTbgAOewUFG8ZvBcPCJBzrQpT/q
zakiEQvla7tDDjo03d52P6l2CkTgr3ZxG9sFbcByeO+3wMKRcyMx51xZlJ4MwJncjzk0EEO35qvn
18REAhqsZesztb1gWISeIOuY/oW0nnnw3k4Y8tqSyQvA9+Iis6maCPpbjTdJi6kUa83dels7sboq
oT65ufyJtYyzHh4puAq5NRo1IAbXzU3HgsbmLaPylh2jq9Hzfgfbj5BdoR1hflei5uEaNQMELBC3
CWMYlabSjlKR+As7P8wmg7E5ksF5fL9AM0/GlO5upO6DDYfdWS6hIjdWKnn+wDcb81NPxwnS/s6A
QlnUn4lYemcoTU8v7Oh0SyTUWv2yafRKFgEXTaR95bY+H/3GNt09fmzFtg/exuinegZfMbO2ip+F
q4dlwFnNF9KwYZiScHemF6mWhFQOjjm1qKHAMij3Yil5jwnG/Aw5aiYh1d50hTtB4C3zYG+6dKPU
cCyRGT3YNvEVbxVW5BJwjGftfFJflfIb9aBbo6pRAbAprBgHtPA2F/wVaL1FiNwfvAgN4+k1bbnZ
Tii94Li+f/OJN1uC28YMwJWjtqXsbUgEX2YudtvcE7h/5XwuVZ8ai98CQAufbAxr9/IlFpbLLm4d
uiH51Etw5XxLvTNOIF61TMHtYCN9s5J07M2lpvFSFhKEvWzhT4eNuT5t9OSH8y28HBM3R1q61bCx
zH6cZa4KMUYdX0aNWVB7mlyYYQvhXUXI2lvaS3gktfu4b890D0mxfrKCe1QfYkgkARgfc/Oy7lwB
JCgQIFnDbPh5evcBh6tPztjHHx5Qxd4nbVkhF9DbalA4BEjGW9rv+dR9B36CI0vUvAO/U9FNT+yh
cIQ+ij2tO4NJTbSAY3V+92nOZ2iUPmgWXC0YibDmWvqqWj7c9Yuxs4mFaoW0nZF1CT1JjT8qAF3h
cRsfsdptVfZkx6RmVhpwAucJcKXwblPN3Sd0RJv0OlaccdrMZ6B8EUiLfiW1Ca6ccaOwKhcA/7MR
LH14XI5jsZl/dLTw63nJzT98pA9e781Ktk35LLeaJK3D4WxT5N0WPPRfc8ooNXpyrlZ7s8eAbdFd
lzz5TqYzzq0PBYNbr5jJAfTquNoxpKwNBqPePl2SnbxZX246gzm59LVVdPTcbbHsh29z51C06YG4
79k/j2RXeBOTmFQF2IZ7aowZqGIRY0yXyenazKBuEil+UokT9v26G2g98/gOlUvd5tqBGoD4p79p
KLWSJ5ebp3nWzeF51qAlPW1Yz4tUZkYk1OoOZ4CxZPIle/JjpS5313Z7nuR77viRUmIxHETvMkaa
03snLJze/N9mREfzIYXl4RWXX4NYbPr+PDhKf6csim+l22YeSJcWk/v/wy30zoHiBH5YgDlh6b0s
HvG2KCq7kAeXFSUCrVKexiFz2Vil6xvqUEnwOuNYR8vSuZ7E/QtHLiz9Qw8xs3r+41PoNGQpqThF
a5WetEdn5FBEVIXNyiSkAEO3cU6SxTuYEvOPuvHvUcgW3snMvKlr5J700zYifI+umQxBUYL1Zdzw
f1k3I7r7x3Yv0u5Lg6U5DudE65znLBTWWfUJ0vyLnf8SFIO1Mot896Q4hKbKw1JZF6me63Kahb9g
HN2Zdt7rCZFnXTO77ew6QFNn0aP2C3chKJsQN3BEpkRBLCWycqxwJrbdgwRfauSIztihP+Boj+Tk
qtPEgv+Q8YnTuGKnNxE2Hm2S2OTal3BqUZgL8t/E00Y8oPhb6rRWwpN1EOoZ/1e7JYK1zaVQMwvz
ODPFStEnCmko+HBwZBy1m7DU+FvT9LThKSa+MXNtgDJtsGZl6SMbMjzTHwCpY42ZNwOl125dz10x
zFv+yu7P4vl0xEzRQA/rSr3F5IGbY5BaYSt5RJN+h9XpSpUMhDwHaMZiLjg7mjSQHcYmrBcfS0w9
mmQfZNp2iGYxJJ8JnAvF4aePRGQh7Z2pEspPGjv9Qf90GKuIYJDz/gQelnap6xXuuhJlCVFY0gZM
6j2OTRyRLnAe5QCFTM/jFd4v3yc/IWu7ZMtCpF6ga3lzAMSqQdijw2dWc5KpnFbVFTheBKKuVAzR
O/y18OyRqQwcVI0uk2jvJQuBSY5n5J8FSmQOmzqOL1tMTet00ZX+3ctTtwGb+QcxAmYEWjRtE3yg
JjE/mJgDAhu7NJPgqPUTfP+y3WRwBOiZqbwjvUNEtczj/AfR+nEvPgEeJ5dE6qN+5fdHcIIZE0io
Tpe9O8zMmiMq4nDHI7Hfevbmnj2S9fIpv+jici++y0RHHDB/8q2dOXJigMFW2cQ0yP70pUil+bmg
DHdfLzvnjgPD77yTBPmxTqtLedCMAJPjqrjspR23HVliv0F87WTsoDYEPqr2Vqrl5rYombuZ7698
VUMsX5Iz0d1RdR0lJUnxn1INLVCdUlTeu1cayuu6hWFIqNLA9Id9l6YDhl2mx40vPjDjYmYrym4E
QGxyoSjyUj9+mt9kTRU3CoEZS1EY9egWR3NgSssX6M+J+Mq/L5BDCUkGz+25BxCgOz0lPnXBZClI
00VBnq9Xe7aVum5YYYkTQMK31dT5tfca3OGZYEE+87/LIVkqRdfVRZfT6vf7dIXA+dYi9NP6hXTS
wBMjSLdhESAN+Pzrakyfik6uGDlXJ4NkrqhgZMz+dWoVOj54koup0FYIPVbJe1LY440+nHO/Zga6
wCCsLa3xog3NOFRCbu6m8zeJCbcK/Rf4DiUvVuch4M1OzXA9KScpskbggPFGuPSGn/iB8s820MBE
bY7FbZ73BJuU89UnQr1O5NwRqhZJQoQRaEdqu0CTwblHKEE+9Ps77wDFL7rhRhAWYjjuWmCuArYZ
QnZazSalH5kJ98iO1b9ZgCsszg0mNoM5hLttlgEI5DW+5JnaU4q2snY0yOeJFZhhtlJle5rG5mDf
amkVsfPx93QRw870RaMc43lE+btZ6hWnBSEjeKjK3W5sOSOrecxhYConAL5OxSFLeZ+pvAuTTpjF
+satbVamY3Ij0tsdowFhDJpwJIuhKLL20pmmhJgZyoUXcrY8mxYrWHOrpcIGBZIxxbqyO80wjFw9
DFMR7kma6g45z0/5oFLusrfTz1LZlgt9FcFS4HsC8fY8jS+O6rbylyiQaWOE7rBHo7bqVQ59WrzL
+OfFx2kzpOMwGiew6BsK5wbiPItoHmqx1ucLowA9O5TfkpnhbbGtmB33pdXVvroEESybi5LxUCiD
Btcx7WhpgMYpHOhGx90W8ogfit0ejiRFBr3wK0k/6Exo0ITnuEEzjnSJsKM/J/Xq05+A7tsFfSK3
SuVvl5IFFhGngLLd2lbOLw0dZElwPvmTI26zw9XM8OEYs6uTM0dtieTT/xLo+CZ/vLYQ6xuxmwSE
B+XhklQK/B7v4Foef3EASZhAPOg3AwveROhYSA8TVaBWlJV/l2/mKHFQN935V8HCadrfSlWiHZ8E
sFDAW1tU8X1B261CyG008JG37+5+fKY90LjVx/Uvq7anPHEH03JYZmUiS2WN2rV3mvNgSDgxV4mj
DJ+N5u8ENbZMdncO3VkxNcqmZwX9POd+2qYPM/4JoofxmboThEG66vUGX1YlBdMaHoTorRr2H/Ad
vWJQr6JyckMnWrFUV5A1jSYbjUg8LsAxVegcFhq/G3iDLy3ubmueJHdHZ/8ZCpOCf50PrnJ30P7S
84jLPduTM4gvBDiRBq5OPSAGIQwkPIVTfNSkL4T4S+9cBRQK0x3iou/e48825+kBv6Ve42O7Bp5Z
KUXRaRWIcwbl4qWq0BumYHYidary0STbAFkXJdb80iZzcllS67r5KxptR9QtT43ViRQGIB/StMbW
FrpY1iQ2/dwL+LPzsBS2ziaeQ0JwSHDT54GGbYHyyRQrLHwbhhj/i1bjPPxp+N+rn3hGmIEcuhZB
sOW0tG7yfyMER9sbmrkZ3XNwrNfOkvoKgMZb0C7VjYmy7Ol0xgLzS5BE4uTO3QGhKNydoYcXLhYN
eXCUgbGCGYrkt5JSvWjOfhQ+b26LloMcZSkOf3ZQAI+oCkw2Ep8zH8ma8GZYRWdmmV39F1efe/N7
RGUYo0fhF3O84mL0yY/Cz3AmTR4gobCRs+7qNhnoNNgwaMoXrXBMKF9rlpLeA1S+FywDP3IkcIlb
fqICmH6AGz5HvxOfCnxbmJR1jnbKRRzNiJ+6XA6Q1uxbDuMlQzdSnG/FLqOEt0CfT5hOZWn3y0Ig
xYfgdz0tAjyLsV7u3+Jg1Uc4wCAOOpu2lfHf6wuVVUxJ15TqLNyX40dIwlUXnPdJ9kLn08pkmM1G
nyfqBKxz1xe8CqXSmOEisjQqTNxVqU/x3tEZQqolyT8em/xfF1NV/YW+NslZQj2aX382Mcn90cRZ
225j1bisjYqfoyF2bS93+orQMdR9HY2EFkPDCiP4SU4dixkqSAtq45Bc066DyN17EkKpNIeP4NvA
ww0AkxN3c3J3/ThehyhB21bOUh7LJqIepzTejMzZlfpJCs0DZb4a65BMtuPrijuDbANmA3rlq84c
uedVhw8B1D/RsYpA0ZOFYWC//WHf4EDdGXUK4zO98FWPyErbqR3WXp7ukmPSpbw1NkMxfUDuAyv+
0aAkZBfCAOSDcCook4SVlULpCW14/ejtrCRXfqkH1abMveHVhPEW9vheY9dh4h/aWaqctMkX/vCO
pWQYjpuZPRGoVZeRHsid48ZizDlF11qTU26fGWTe7g+8Ltx5lhCXbfCQVBAJrTwFxvuM6owLY1En
7F602YoczwcX92c6acHjoFK1S8MgwfRNK3xYalOIPxCtx7k6JwJ5IokZJs2qX8QZoEXVRvvMi6/9
unuUKD0WxOF+wnPyzeOXpdx+HB1+V11+FKv+0jqtsPO6pwKjuG3b13lfb/nsyIaUTZ4KwFGf5Cs1
T2d+z9ehvRxnLU2/QpfYqGtWfc1LFR8aEJRn73KgSAGOPCG1UK3qfIo27ccXy6bR1SxGYNa2HIab
L0VmRG8dv4wrcejHk2nmb3Ean+xdB+ihxyiDBM0gEqiaYC+9zKbSi4W0DPlPJ/jDvV2f/l8C1eSZ
CsTdOc9xTFqKNKamky/R99wpQq5BywAHEYPxrSEoIcphbDArHDmGVL3ApM5g3aDr31DkJB0KkWsp
dkBjBerd/H06dctkHxLAeCVPboHJnpax86u27dXS+FVX5At1N9d2B76h3AC4bEQQuy2YeZIxIzjn
7/04S+SWWih0AGTryueXD/1gGkKLCgVMNyzex4UP1q9R4jRlSx7u23SaGeT6AUPky1waIxCKBBHg
olWI/tc+rifHKwzIXxMFEIzTrAKb0YsOQnV9sL0vMkicRdqooV2hFNt4dzLn29lWAxHqqhsG8nWx
oPC7Ek6jknUZuzUMWATEpIQ1QSkBOOoFLBm+5LQ/yBW2agtyr6UhEb+ekzePeQRXMBFfp+eXA6Lw
ZycI9aKT0hpuVydyG/2wj/TNSRQINJMi1ezRoZ8XXW8giTq/dQg4EiyLkatEomn+RcJwvkt+vjT1
k3ULXdCFVhUtWDiSQGFFwgjU0gi+jA3GOtW5GkbGkH5wGgihdmFCChzzoIX837xbItQP0ddB2r/t
EezSRgPNPdV5eZKK3wTwKOi2GLRIW+HLxRYW2f3GKhWktxCHbFYkHOOccrBQCihac+EoQhmp7YQY
IFO3eCvohSzArz97v8k+ulvtG7VVhsbPRh0+ogI1BYP+iE7JZGeBqqcav/YwNu9WErYy5YbrVa09
eIRdXEWj3Bg+Tj6cjzIV4h8n3AvlEVrol+l4EeOuW50mtuKfkJGac6kvj9Ijk/u7EBTyWC4CzdXV
ePRUn/f08/0paNH0OyYE4nI7Vlcot6ZqJeMvA6F02o1Xnr5j7gB90wZ538WA4of9l/lPkY3XzFgz
bJg6vow4yJ74UaVxSCxgrH3Km4pDRbPEYTc53Q8gguZ4jTdBXl4JGbAo1TH/FNMwaQpFsXrW8aqU
Bsl5Af0qeHcLvp/dSDxPhFuoVcgs7YtifIOQSL7A2OLUgPeC8j9zYZDSbmI8DxEI0xman8Jp5RS6
w34pfa6IzvCtDXClON0LZ/lZ+fxaaGH/E1YXV/PwUqxcAc0PybMWMcStw345xdxpRJddaSDbFU13
u51MJ3egOCsbXp97qs2EIc1Ts3jg1hO0V16QsqR2QA9OluRIFn19Gv9ZajJZBXI5kGgyn9sHxMuk
X/Z0vKLIrOyiOoN512JDWPHxFDlyhWWkNvXM+q0v7KZjNX46ExOu2GPvMgYVw68VlHtd+OzdrdBt
0JIoICTD5p0Z5plKyDemFljpuEDKN8Y6TJ4i/SiE+JdZEDLaCEuZYJr15m0YtPaklQcQsPdd+RtK
hu+S2aawEPOcUpCKjuBIOUptUhzzQfRIylRLaPmJ1sZZX7epi0rabEqk22Gzg8MgOA2mWnR1OLVF
CjD2ESHOI+3yWjJJZiuAJqPmAi5H+AXV8X78vQrAbrUdcELvAyywFA4UqY3CEK614A1E0vbAnpeC
pOuMBD16l3q5l/RFIvlu3uYGDJ5RgPcx0BHW+aR9zhw5cFQvNvI/RGy0wVsydMm6d4XgFLTsM7Fb
qmcjkaZ1rsx0psvqsHgxiklj88SwE2Jv3IJ9AsslBmrcTC11Yz/7hpdhKgnLIrR3oujR9rLV5+mW
E9SJ49oF0PVi1bUvL291cYSaPPS+nJoIzjj5jkrboITv0OyNB29kQBu29KTz4VGKV5OaYq8lJWT6
RURgVjKgka917VFZXX3uVriuBFoQJqiJfgw9RSVNioVfSSTPXfb5KKPavD4uxAg18J39KA/wvuCF
cy+SdDs4keEOzn3Lx4LpPXQnOYZOGJiKGexxz7kE1b8cTE7djnbUVGtXatbwOZRNFo5YAPWMIFbR
rzGK4P61Urz5yJVPCCVvpxKFGxlZsh3ARHLfAWnUzh9C4+6idrAfozCNy7LHMrZ6Gi6GDhxS1L49
jxw9aC/ccAYC9M3cG05aEZh1jCciVWLroQsWj7fJiyciJP2xue5++njOrLIr5Crf71tvhK5l6I1F
ox+1exQXEBdf0EcpfUUkJ5mDHG3+9HEl0FaTgwwT6QNOjdhHfMtUFNX5Qt3acDXDuDJ7oHZ4VdJO
A78auGtAiOvLewqt55hkR6Aw9QJpDf1ipOgiPIJkuVfxM+J8tBuR02W12KrN1Xc3Xj88ZLoUDvt1
JdJOHIRIu6JfoOz9Mbh+NIxzoKWJv5rN2fsW/fDeUPlTCcuTofek2SbOEYpaM82+mjNxkef1HeX2
C3ON4w96od0m6BdMx7Agoil+sn9wRiLvpi8kSpx8yN/Gp3hwbPvpdnHwVgStH07+ntHiCl53qsNv
dfZCeqQTAWW3T6fgv2eOGOhYc0f7coXBHenUcwv/+1gnCYOVEB8csLk3qOaO/dqCykSb0idanRIn
EM8ZPecLfTkYcOez+0e2YLlu63wJXmatAwNbl3ieNcl0lX8/JM17W2AEnIG7BtIKeU8gtwa4Yq6Y
Q9y7KPfV3FvWWu8WlyOfUjpgejvz6v5Leeu5lZQy/d2SRdB18TJ1e+1Gl9bHxUX9W6AuFQ1q8tyu
mhR5/QDKQ/JcgjNMT/ZW2vManl9FL2K+2cALYk5B7N+qRvDMELbRpqrt/y0Qez7f0B/mOvhu7AJo
w/5Jy9ObLYiIXgZNQE9goSd2bTVth3u4/AGlSSvMXOt/dqyp7OJStwtXhofYfu40Jtgfkp6+QEfO
gYC+6WVVfW37D2qdYMxAINc4hkWbJhahhWWf4LTLZmsxR9MK7wI4FIWoU28xKtCO1NKTx1Zhi2zB
OKZ2AInkwEyujad7g59Wxb3LZ+m0h9D4+H/0zUb8NYia1WBvV0q7A2V916DAfUPPvlxYFQP7T98u
ng32DOulGkSjrhc/M5rRTEJss2c9OMVOb6tGMkKKUjabj+LlWBAVIDYgwskUinOOVfUOs8j+Z71u
iBEvFq48mEZltfO/igmeY6UHt1VA5WMm1o9f8E+mqy3oBbgRXifUYwI670EjdnOpGUBVJQv4OOMf
I9Y1YyX+VNMA/OdsQ9fP37OPnMcko9Ti5QDSJOmfcgcRHZfKWk2JKs7WK/btw6B7I8VZi+s+lGUp
pFzYI4Sj0Ec8sV7ycwlVYQT6egEVPfGlqhAwkj6N3lY1mCFxrNrc6KkRJhO+nNeCAwA0sFTiz3wS
tMSnXthICJJc2r56R2qVmO9kAFqTbjZlixFtKAHd2FW8LHZLR0Am1dnqbSGqI72v9c2buLoaG3gu
NqS1RMkb7qb91oEIDX2EqRNx5clNB2iNytYulScx+aD5pQdn3KiNoQo4JyCTYOrznsxStZgaPda6
20KbfkhF4+mV19DsTAhRxqn+mvCkWRAha6oSzbyXfXJ9Qc5gHQX1i6uiyCl4UgMBrR/K2bg0qR4r
3gvS8U0YDikHOR+eWRHhv7VTBE9gZ2cWPQDgBwPP6MampHu5z1kUdsYYZRwvuvavJmRytU8Q/Bf1
65rwdBMIDU+w0aXajlYVK+58Q2w409Stg6RC3BbnisWGhf2I4d2C1ZQ/aPT69YL5jlR5p89c8mK/
oIGisWIPuHyxNzQ8HBSI8aHGVCn/OIuR5vJ7fGibi0eNzvkNpw4PsttjmCpeS0ytK4v5HbnstURs
/w+y/Pp8YX17JQUfEzMmIGmAoZx/UvvUb2oZYc5Mv+Ti6mXjDazchIbYiodYvhP5cQjkTpkng45/
NU3CqshJkShSQfOtejHkueCfMx5QsAZgFI3QQ1TNMWKhg81Z53GIILJmVNUG5+C/Qs7emu9BgBg5
EtFcfgClHodIyG/10wIhSMLDuVZyRhVqyYmbG+XTt3wsJK1rGL0ySma2aeo7UW14Wph3WBmcyXQ9
Y3CybPEYwm3d8OS01YblCU4ur+8sZVh1jbiS5FdA524G1YZB0QkKV69Yn9eir76tUroNQVf8FnSJ
WyaNY3s47GJnByCv6/ea94uWSYqaZf0uXuUi40xki4g91xCtLHgN8h5cNG3gW6+oMAZhxg9QtBtO
Gc44InFDbPZ/5uU+B/x/lAHueuemuqevFQD7QA0ixWaUEbD3xvBdL0F/cSuR1pr03n280D+FmJty
9yHwAINLEoDpeke/Cyp6r3AcG/9sknvcwZgMsMgi7/1NyscH1r4X7OCo+gPreEmQnqmmwB+ZwTns
GKdkf/vz41lc4bZMGGtLsshqetGf8szAVHLOXSWPACFcB35WbJJEvOV8Z4VIv3XIC2FbE92E2X7r
W5Gf1/TLYwCVyoeG9ajm8/tqeiWCFhH6RXpjgArxuv7SA9pCaRUywpSAyxkKhI5TQv8Q60jqhtZp
g/HoKIxbwkkzPlGjSHLzThHqkhcqCnbTu4pIX00Ae/aCb3q5RN1sy1myyLZ3y7uzB9VN6/XDkWVb
koa9cUR9jYv8VUvU8NR3jJXbAEDfGGVwt9ReiEMcAzGXpgOq39vzctu8A3vF/ZS+HXZ8cafBSS9G
maysdsx8rMDrnZWGs43dFVW9dbj/h85Ktg3ynZ50BJahWtAhQdIl+UvMfVxQfILfaGSIdZ/oK/LU
AVzX0OXzed9lzo1WJ7vMxRsMz3SXUEhXezWk8uCohvjk6w94lhwhGcko5Skb4i7VbekPuKEjTYoS
6/IGWuUXQ9m4mO5uzflz4hBCrZ8dxNPHDXx/KodYEDb1ZCAmTK13Nn+qIxEYYUEa9sLXc7MXoO0c
pOTjSb//Ep1iyrMV/qnEGL9QYlklpI8X1oa3YIBaJV2T4fVsVGob/QkmsFrKAQc8seGB8FJRtW1f
/GqVzDMV7O/d2he0qDGvqiy5UJRl8R+JSEPphKt2WsBYtl19d3kHpJ7Ql5wnS0TYHdYjysn7AdSJ
UKpBRREIRdTX1EXRB5qHtKq3LYVyI7fxTM/0COJc5r7qszh6ecxRwqK5Wt1CBZ8gE+M10BLn3fHA
O49AYPq1J1z0HgchPCSYpzeRVYe9/+/CWHUEsgyeltJEbXrtdxnhEVzFo9CLt49CcQS44AQOrB9o
nNT3aevO0u599dSjkDO1z6/KXrmUNhCpS8ewtuZTgn3ZkoAkXsAjS6e93Li//oq0nwnSY8Uz0jwt
6qFOyQwORJWK/ZQ+7q+EiyRabuMi8U7XM/ICaQXMUwKqrv7Hkk1+6UMwGRtJkpjrsXhG0ffbpWrU
fnLAiFi7AB6i5g1j0LCJ/QHjuNKOiQPNNKVLKe3+kRgR3pqzIGFzkhrZ8DgGCnk6rjfrThmoVCi7
RdLj+k7IoSxFyk7GL9X+GofSrPt1e9GjGjarej7s90l5iDGoPxD/BwMJkLlmQJDOXdH3GyZZOljt
cpPiMXQjrRszWG2rnx5E8RgyfaMI/W6cR9O+Q5Esozd8+eCBFaAUxNgjD12ei4RSH9FD1GRfl38t
dtN0uNtW0M067ou0HKOnTlIK8pSCyIXxECZ0MReEft3NOU8vdRUXKmQ912u01/FkLtn40gmKmP5q
0oZE2BR+gpjxWu/+p8TDnD267mapDbUT7rHeBerH5iqZEifTOv36VDeCv9gu+7bRAimA2t7eSl1Z
UKMpgiL1xpWHx3ZBkqVGryozceSZzKo+B3COc/xWPTOkDYUtjnIJ0QZ8JljIrPjuG+o3sN3vJQFJ
dQ6lMgO7zfRhXVz/YFwuEOCip0wVLUyosbdNAPotD6Fd7pTsEsToRnP4d80Ikj9oCNTYjbjo0zrR
nxTrykvcUDjL/i/iDBa8Xrh8NHaK16eVgoFNqZ/52p7gJSDhWT9sJ+jPXiKaPIUKddVfLf9CBkLW
ON2QU2SxAJWfNzV+NT4+jydnVwlHzJgYrWr5XhtOnDkWA8ZC45yOD40gNrGI6qflvQAdOPqs60m7
yYW534pE/H2eekkRvqxQ2HPxtwSLLg4JPaZgT6MsU4pqVvn/0EoKGTcbhKW8iYuF/u250nQnNzr5
KKMXrILU8hwhGhAc8+l/qwMsjDD4nh1S0IfnrsWTlY3/5tayeSIKT32203NS/Bbp3qYlbUkGna1d
2AYHH56iVpMD+oRwGDSigJgA3uwnnSnu4gyHH8rwCdq3Ffqtlra7hRU25/Ja4bmtKSLokb+V9Rlo
4p2EhceWFppaZy1kEoclmDtzdImiAQa6/BlUSuvwt6WtpupVtOC5kLweG6CBU1teazUrS2sP7uks
8gcFuoicHph1RNO+TPp57dcnm5/C87mH3H4VTj6XS9FaL+aMsAukuu4w263kzMzzbivJy4Dx0lwE
FW1OjIFfZkBHlkvM3riI5RiGRt5igQCz7QmEQ0EeY4bnXNv5UiMXrnTm2b/TYACqZ/t4hSf+RDC5
oQFjtcsUKjM39d2QfHdJDwaRAwRu6teXC9HSiFXkVibMWsBa4p+37PsUPtVxDq+9Mst6vSWfQBCQ
qcT1v0+ayVQrUS9r85FTr6FsL1l8++czCDQE28Nq5SWUaj2UPoGjAL2sqGNdzM1fXquBV1INnJ3M
I24iGY6oHxlUA+2z6cLoERwqbMFC2qGm0EMCF78u57x4yuey1pDC5LQxYuRIIo59vIQ+wMGALpJf
PyxhA2qCNHTIhY86OrIWqjLMTvCiUnmcL54XaS4dMqgo9ucvxhC2Ynooxyw18gCt8ppCS5U+qbOA
j4kOf99S/XG30dwXlkWUijqEu1b6GCgRw5VDy3lpPDNM88v1YyMxP8Lv8bID38TZJAoOvhIYS88/
0Q0iJWBTD30b6T96GiTzbIjRAWSOQFEL8br52fZ8OjgZAXbpUJNyjBI0Es7GiWFh93GIqy1rGVPC
0D0mbBcecRInL+41I4BhvBeD1lIf01bzu6mEMQSA8RxGvcdQujxzY9HRwKh7hlLCPkIVjAe0E0FJ
cgNjOGHGKMcCqOMWXvyCuqeULRdvVEnP7m9u0G9OZNxjWc/6E/o1yVwrNGoieKn7mycZguP/DN38
R55tToaGBVIKlTvWOr5ytJYaat/RtWAmtkCx1sl4sq2uEML8D/Y2NcR6SQ7dXX5iXUYAQgzyNvG+
TnOaWjYYeV0v0IBcV0HI7GMQV7bESpS8NY3R9Xpnw2S2+2fNRdieWIwptms95/WTBLmoqZXtcRPt
33eABDqAA5frEhiPCn5r0wyExBj+kK/Qwq3SB1EKB344AdMwhKlmQRTL8aKmB9cWe/kLPcppAcus
Sok0h8vQAHohREqnJ7hajaLmat/wy994RJ8HLkvmlByoDgdiTFOFSLJSyvQ7Sq4WKBi6Schz1l3y
H0zfm6zT2POsTmdAko+QdzfAx6in6xtPEToLnKqYzTQnKLT3nneRJilcpzLQpuuHo8hWfHecxoVf
T8rFk2mvTRR/dtrWg7xLLOGFJo0ZU4inQnhWbh3JVDNdirAWlsK8oDgwIgnFmPrt1Caw/mRUwFjB
xkEzJXXVn/jPyzHaqX9siZJwAKMHJu7/LNB2dtLxe0Cv1enj71njuDF0j3+JOsf0IMICqH9ys1ux
J0qejxK63r54ni/BRms+YoKl3hCRkB9GJ3DlZ7qfth/HXTyrwANy5DHHr46ULCE4wCBvXfXd7Rph
QvLLnWpraWiAmLxCk+8ihmjinsbp3ZY1epxUWpGxCxnKSW7Y5MO5eIuAwdSOozh1luudSOA8O+/y
DFpQtUS/Qp7DCdcnlkej/mblNEz39iBZyZZgKXt90SRHcbgstHsyCWMSNVSehs7tRdpAA3qD/1X5
TN9WluB9iY5yPp26AlxNCF7ZmpDo73pkpPwoCh9RboX/3e7gS/myjK612GeSFDv+ohpZkljIgvfT
2C0MXJ0PjRK0IbIHlDupeAfJt1AdBCeGbX4e8/Q46ZjYuRBPDarL7crFipfAeX19Fs1z8e5kN4gR
NNzoLoS00Sg6w7peTKCCVyfH1NvIxhJuieMXI/cCv9bJOnRQ3LsbU6OvfSRNRG1o2F9p6SXS6T/S
iMUeNmghGhvvLHHCj08/gn1Ih8dmP/e8igL4kEdDqQnOSGKl/UOCALKwZ7pxJY3M8PUr9nVNpMUV
ZoYo20uBI5a7p8sDugnaO/eTpEu6szOYw1lHtrsn/Bs+cR8TwjJpMD36iJdvawc3kECngoDvq/lk
y2H6AwxGtQAaClw7/fXfRxUpoNwZ+hQxXgMU/Gbd1ZPrtdEPeihj6RFXznpyzu8rRAdHbNhHEv9Z
vgTt9xN5s2Pl26OTp8ieXgoqnS/q2tSMfjDJ36t7AJSu5YFhENTB0YlR8QEKYQixeMuMi4y8HH51
BgeaolcLDWQko+Jf/uOT+e8dpWot/GFFFXjHf4bSAPufdDrCmPC2zHbAHeWIpZ4twmyNGJojtOG7
EivmmgqVgXIvQYnXWkNPNeaNmDsTJA6NxFDEQwbwJSxkg6yNUUJcYOs4WGuHHLmP6DR3ns8aEZ1S
TCPSXiyYLToKX1aoPbFZSj7Wkuyosg39Css4tiwGOplU4FnGdDzZQ2jD14hPJdsCSnfI5Ufx+NgO
hnY3SbZ1b3z5IvmJYEcYN+tlFhrNtbYEDOfyDDX4lUV+RBqF1vKxnA+z9C78vpUdOIQPIFyQyKr5
R8Ed2VmtzyrGEWKHYK0hQThtD9FA2EA23QHoulCrCow34O3iCbpw6QUIbf0NrkbLI8cJdVzsAxhl
j7yKWsugtGCTWKBCWkOYNjTk5aQpjExS16I+xr2gjVPx0NjdfbJA38d9eiSDyp2hyGQ78JVtrv5N
G4pVOYSp96+P5R325XLRwtUcpzRjJ6GZBgwtVwy7A+LAWQIoj2J+52y2JwPbUKKQXpR2yy2tG3BL
BGHLlJW9RhcNt7CHqDMCzrgLHeCqlisU6O27+E/BhT3KuslwsusecYWe66uNB+FZLzJhajFRgZtj
BCEUJ3ZK897ET34oO5jbzxUBt1V3DFvfPJ57zd/C9cwxb9fNmrz0LrTlwcWsXn4cZjp+NvSm+yVm
6GzqCoqnOniA8yFV/pTaD9I2SsPzqVf2sv7kshg057ZtqZDg9L+NCNS8ehVS8RqvP581s8ymrhVv
Als3lm4ubE5uxpeleVHmbsJhUReORZJq8gd/m4v50kWMQZWoNTdlihUf57/mCiPCD8Ke5LoQ4oZg
dMS3FsgBL88/9EuK8NCfCeNAg0asWMaxcHBQX7QZaXKg3rZE/1TO88+hZ7CU25/fXkdQXK93Rbyu
AqCES+B9KlukOSsPtSA6aI1ePSwgwSpJFW/TIptgxHW5gKozlVBOdDLQ4bhzxXMpB28EYbvu5laC
F0pljcjMbOr7/YTQgjbUn+Qbs+GExvpBUFqmNWBATE7chYkR5vh3vUQp7jTZUuAZrF/3Lc0fays5
a9oLKZIdwkqeKnTpnjbeqSrKq6TeD4uZbpHHiRZTXg1U9Oq4d75ynlUJqP+gkwCFBVG/atBIBGJT
ctdTPfOWtgXrYtFzNVoJk/mTTMJOQEohlbmvMeilPiG2yToGe89Olg7OnWO4KuAX5eUoQK0ntzPh
pBR+pmVNqvF5Kky2EzK2sp9Yn0TVgOzVh3P+ckg8ledV6LPX2a+TtMPQWDUNZluyBFHVG1lmF5Nn
vojJs6RBPibh/vDxxSL0peRM5VMEJh2Zg0k5b4mwrRcIaP/xOqpdzLIS3paNA7AEXVRBdcEjCBBV
fgt4zDZRcF2oCOcHT+4sWltatec7g2/lp8L889I+lYGH5IqdTnuatDyeKCDPR/9Z0dn0Sy72QyCA
xoU9+tAv5KmyFfrLcMI1vEFdd8P/gRvTAwmfprAB3fYLSAXLsFuV/lc/2vwpQi0EiSCWsYqvtmlX
C8l/Q/WhS8i/31cNMn7rIeR6FU9BjGYJ/pyTi9aOOtfgI7kCIRzl5m8pKKx4yTvoHd6rxzFeTJoB
rafkSaXMQuXkuBleevdKB/RDd96mzWwXGaWhD+1pAAQzASxXzn39h5n0DU1coRPeSlz+7WBJow+e
k3Sfq8QGMK2yEcC7vkFjl2fbqOGBzIrf7qGciUjF8X+Lh3BRve5kjUvqwp5BZGUR5V4YYtKtbDMd
Ku8zoIxPd4cI4VE6ZDQ4D7o0xjgyp4cIfaNIIVeDKyhPMFr6tNIGimXxe60BjNrvXtHmJYRKhrmj
sbY0fXfPcl9D+deJg1f82NUQQNneTzDeIm1drR/9XE5kGj9r7TQ/uuRMJ7kvbaHYzBZhCZL/LCsZ
YITat7VsS7Piv2XCsvMek/IBVThULnFLRDQQ+WMUf01ryFYk59P2crSDpbP0ZcOfSur2abnbtjgH
Ff9UWH2p7hTPPPRwfHD48wa23ZjVnOu1pQ7S2zssSnm55fcai5CT0inr+saRouHsFb+EEs+sb5PI
3UseyBaYc7cKENNarVKiR39kRMD6fV8qKTEcx9mwu4cd+6UyUY+HaZkxfDOQHLAxS59B8KuO1Jzo
UqehP/bHPj5i4/Id83zU5cVTrMJ/hMweJXNEVvqY/KLdYu/OuPNufcVBd6Ntkg5EM4bHCpHn3V9p
hI4zLcNW/iD3taz8lBqc7WiweqQpt2JMkYmZ95NezTMqD3skFX8/hXSRKkLX57JtKFh5lAPg4tQj
W2ea6ME+Kj5p5Df5mFqbq0oaj4kOrDl9wkPUU39Gip1AMQmkoq3/7FDjoxeuKNYdIahQ8MZe+j7N
Uxf+Ri7c97384EfCxibVnNCRZM8Pxz03lnhafvykv5YXh4Iykk5fpcDcc+0YfN8wRJ+dFU1gHmd9
9DL26iy0llUKLXznavG+POQJ6TMqKIAtFVNmCTA4QYg8kGj4tf6M6L1jYVYBJ5qkuoe6UaS5u9nV
urW2E7zENN59Hf/h0F64I91Ay+YPcSVRMne2fAPxc/WFcN0kS7XYGic+PBw0//R0rLK+KWpbFC06
BhzVn3nxzW7nY7av+4GRezJTzZ3TPy0IvHmM/G9KWgJoPxZWUrNjDGzVm11uUb/urs6dpoDfzwPE
Fd+xR1Vk33b2H7jLBWK8CccBgXd9xLm4SLkOi0lcjZh2aoaFhq2ecd1uf2lp44mLG6gOGQd92wwr
jqUfGxrTREw1jsbxC2zOtprUT8rHOEBZ+dkrY282FJXZhEZFOoBd3DHNEHhW/icVGeJPuv4QGikx
FRq+Fb8qKwpGVGCcHsGafxbn5h4hFx79OhmMOz8rMJEHln39zSDJsqbRdwa02T++KAYuxxv6DVTY
n17UCoqSenjhUix9hqqIy2nyJcp79g/YeoqIKcfuEvjrESEJksHXg4M/Q29jVVjik/l9nvruVqej
IpZ8Kwg33kGjF/xOhfFn+LrdwQydKAQsJmZY6mH4nb68/y9X2Q7vMDQN0gufDn05ql4jYzpNFmpK
YAr9B1OVa0eesTzd9XNpPq3E9G7fNfHTJPUJSkgMwMN50cx+12USMLHhj2jaFfiXFNKnSv7Epcwr
lmf0wfj7nBE8JSQ7O4LjqSNgkzAejpyiQYjx8fc3shvPpjlUYnwpyqko2Co5XZkP7aA8yrehoKAp
HV2Sv+cUkCIAL2m2QVh+ZVv5u5NE9Ee+wxBZfsy3PoNbBi6KF4C7Lxcpvspn35J1Ve+M+AZ59+Ki
QBaFdKD6u7YYtdLhWPXDNGEPNKInSxb5pGYhkEDMKQkvCLPQuycedZhEOdltnjaQL4Pp5FuzhPoU
aapfbw9wsECzYIhgDl8FFcXB1bQKfKoorncW4mgdfwXTa1DgZ4hU9f274KBMFBwmojEubZ4m0m1E
eO3z1AQocQ/wynU3gv8+u7XUkx/PXyWA4rRXStCIF+t9Cq+8WhCcwyEpXAp12V73smfGqyJje3Ru
n5ODhtRZdOMsccV4lCp5kJAQwwvA5thF9cB4vcd4CHllJFHyTqY9aVaFgajF0Z4CHBd1cbVyPqVj
QndzLrf9+9ATrN0Q0olFTCnLxM58OyKyLWD4Whd+XrtVvfZ507/IJu2IeAxWYT84hTyu9KjxpLtK
B1xszhUfgdNmiBUfFENWPWI0BDjgPxun8yoeW4svKQbR5C8XUd6o+DAWM8LzB1bxaOR1T2hXePq1
KXrKiocSzbABL+Anlv7vyx3r5gRWjetoJEQwhiNEAuuI1L0SVy4Y+dSTCfJOiBS6LKScROpFgStQ
bFT0hSEL/xqPNp1iKK/1SkDOdlBnXbwc7TYzeSoVNdx3Ok4wRFhaOZmUiUg2WtpwUoUHrorKmmRJ
dK1lZ/xNY6OKZvHjovqmRaTG/aEzf8WDW57qqaalRL3CUEus7tMpB7lOrkq6+aSP9+4yxieifNh9
x7TqNStPnofl2uERfT9xO8UvqSXH7elNCwx9B5BiR6Ixb9aC5Mfm8Bwe1Jdrb6YWg2Ec8zXJ1yjm
d19Y5MLUkS3tFWN/pe9LVBBATx7mgNQKZkiFrFrMZJkkKgnAziE6Lvqd61JxGsiGRD/AGYScR/LN
x8bNqeCbxCei4L11H1y1dj4xC4qFk1lMHua+iNnHmrIjfxvWM3zNrP7PVA3XJewWSu1zR16DOXSU
biAxYKJsWcPy+ScP3AQiy52gG3UMgPcmONUYmR8OjvkRU3D6mmkU2Z6ovooqZQeniiUE/ebMSQn0
cFqF0OKK2NflSlCbxzLcQdAVr7qCHqRK/OcAx62Cnu0B7hoUL+AVQqu9aCVLlZyqigJ/d5En6XNJ
Wi6wGaEiSmv8vYrwFhFZ23bdr3kOt9WbGhU7ISUbG0op5kUkLObI5uv395M2La5drcj4SfD+fbNl
aVdiS43ABSluX++5V9hFohbov75/Sdqeu1Zwd4pvdfqx9L3XN9YAWbSfC/oYSijrX/VrtfFcdRUV
1nzEHCleA602wqLCd4NitP+tbCWyamaJ8uCRX0UHlcIPDfDJpARY4lUimo7Ji4eZIQFDFe//EFgN
Zq1FNmghEiHgw/8uq7x/htaOjCVRt/kRGPub0A+snMf99UasHWU5Xlytr0NBzr5+tZdiOitdDJ3K
QvNBtit5AosHQA/RDvsVltJO4bcmOh/DL+41GKeXYCAYm8KMVPkmIcYUVQvgBGc42LKrARy/Cv2w
tKbNp46e8moYi2EL3PkddZ6lYE8WPd+gNtUJvF5l7GOraZ8Jf4eRJt9YSqcL6c/iBwFCKwOYbKja
O6tL3+xvusnoC15mDOfjivigfbJQVu/19dyg1nRPf7JZxUQJjM1YyaPza9XzAKFrAixUVoRafTbg
fRVRODSoTlJWr4WpOesq3+kiMdJ/ooaNN/Ly+RVoQNy0ttZdsvYFHOfiRad1hGOo3dJgc4mYuZtE
xZ0ZB4kFi1NsvuRemoSlK+aPcD/zkPYM7DVLV7CYDQxNTzQmUPFqdoFVTZZ2O8MT9fluZu8bfg5v
sD73icEni5ppOnLsj690ip+0F1dw5KadVRrxi/2VByBe45lBJbxnSy196WIFbxsxSx8mpA9ThFXk
xCnQpVtpHwVZnQGbjQftHoEIcF0KgPhzpDuwROYqIMCDg1jTvxGMbjJaohYKcj/K/mARELY5/qH+
T5XMIUQaXQt+jQyDPGBTa/NVwoUkOcKvRykngFtYWXTrTvTbzVjje7RkLd6wJXY8Jh8RGNCYxSwg
QhwAETD4cfy77wa9iQMsGwrd7p2FqbHwsnQA6hxU6R7sIbMjhYY/PKEppD0+fhJQM8e7FWxni3mx
4BNuNMVlimP3pBEr8UYdRBvOTVL5w1BJMCz/2LXzaM+tOGFp1Mu/6SSTB2dxmSLtfjRXB2/eLRek
lH2gK2JSge66RryIi5jbZC/MpQVOroRcqzKIvC78dWBg5yiekw5qwYsgM9l2jrpCOt6ar1TFKshc
JRXjSOXtr/F8MXd9dUMCnoqTYwf1BBRlEv9Ce4V9iy3uBL5Z7/Szo4O44yysPxVQqRwngcs6JksX
meepxIb4vW4/2U/8HAcznNdtIRASEQoB0o4rLn5/Sh+8XEJSNiR+kQq647OxtypwdTMk6txi2K9D
CqSDaCQSDjG2XdLQ9UIl6n4IaypJRxouUREs9+PBDdbUCE2NWO5d+2L/4wOS+mSvE6eV2hFSR4A/
oYRH9Rw2FPfBKyiY+yCIvRsT1BhDWjmWYWh7/iQBB/VZG+Ng/xVkwNneh1FDjuDx5qQstx70bP7i
jQXchnxSXmT+OlBiUQfGtltg4kfxGuvmGlrBSE0joq2pz58mEdLQdMVvn9H0xit5cTSYeN8eBItO
OQcdWw74A/Z7VtR5NaN82rQOrsgyZKdYr+EChylFXMlWhB2lyVFkc2V/DHIq4zThtwqLyNs50IsI
GzvNgVbZa1a+ibSmtCYV1bTcyCU4hAKelcl1m6eaCHyOGoM85DTNrnRX5QGSqGhG072YrGXABdcq
ct7HqM2oA7Mrzo5aIi7hOaqHavlw4geRg9HVgQ+Wmc/Un/qwep5QOjUwSAdh+WMalV8S/cxg4i0I
rsa402sGkf73U18kR3WrN0dhps11RqyTiWwa5VmjGiUmO26CNHYw45tS2fCJIgtV2dqiWtO40rPo
l55GhH1r6N0heaK6PSC3LRsrPbpJjhMhlbvivONr6fApzroFKolAtXgM1mp9S047H5d/Iik72kRa
bf6Q7RIpU6+zTRNdK8uxUVQtyV6z8qkSQTzyDfKUJoIhtsRmagt4345zyzhCChAmUi8IiUp/M/Q7
bYCvp7qozzm4JWnBbVsyqqhxHPtwRoiNTABPURHfM6lRUG8X7LfUsKZC3eLjJu7gWubX2DXgcgsw
ovP8vQ6nr1ODo6sn6NrYOkpkF7HoSycojXE4eAT5XPpD4TpY/TkXGpbYQu+04gtwt7pNy5TqRc0W
E+/E2GjCCftkoX0OibXztugcOzkAuza8w4Co2r8S758q2Kw25X3otp3Z6WI8HIhe/5vjSPxr33Au
XvLHuw0lWoxR1rb9aqjFUlUmMmhdqtRcVc/70UqF7BW7Ur03KpsA06g7e0SLGPzW+rv2N70i9A4U
XykIpVkVE+0EilN09ZcollADMmWaR6scvSBekEwItiTdzPOgAoMb9JoGeyKPpg8TWCJch1L96bLZ
BuFyVSk0VKo9Y7GVmHXQApPvNv/pf7aOJoxu8r4PGAX7wegvSU2BzQfKAbf9eYJjPRyPloYaNUUA
bFStwkaT9mnrq3Aj3B8Kr1QMIz7MJhrnxU7CqjsuCdWA197hrDy19RDdPkRhURNvccqXiUTXt6Zm
ODYLavqAhbibh1w16rNZyPBv6DNdtBNkIoeBf9laFqRUXv+RUMzO5pj27Be1YlKEzhG7YlQNQFTP
zUHjxO7Kd0CjsiruXAkAoP19lH/CTny5K0xxhks1JrG10aCv1ndo7xhswg20y96sAcJu6SCVIq4T
CSCsUH1va8IHk/J/00Bzxj0Zje7/Xycm+Ku2hwAlpUIdDpF/numvp52yeht9mzl+/VxGBtSecKWe
med5YvzmKCEnlCgz+pF5ZNPqgygQ4+yfuqsTMFWQdDBsTs2Mh1MwJs/DJjH//3gPb//BUbpNz/C9
Mmd/MRKCedlRRsvOPImj7aBoRPkscNjUL3tGauc/fb0cANhswsUspbPKXy7WLPHGmTm6A+4Dz3b8
ZtVSwoNqIU3LimNRUGl1S7ijtAwFeFqONMy9HoKp9FGl5iXjS1vn/4y5b338ear3geZUHRZ9b1TW
9KHYyQTQFJ7DZzt0lkQhQ9nLSdHv5O+A9+jNrInH/3fM2Nxp7HV92bO4kiB/bLwjMgcpo+NCXn3T
5IQQQi2+vuw+qvh3qYYMvNifgOAi0hxv18uZZZecUhEFOvRsxbX7Nu29x3SdKQ3WgLpb/2/l7ams
s5rXlgwH3DOFWnKMqhNUbZzr/5dZBRYcu1Id1AjSlepdNq0TsiEHNCesyxq0oxpBOfxY9QXKhDkq
gX9HvDP6S33vF6wvV3pjNjeBWUdmTq8F9wMFPL1Uuf9mX5614TkmHtS9TBCPyuAL3exoZtDPL9vL
3YqrnC3UkH2QOEliqkdct85D3X0kCpNm+ieveg5QdIcC1OCfPs9GH8X7okDcMKcA9+HL17Rf8RcX
+xaW1SMrJ83alX9rhgA6kgQ9Vq6QDKnuTxIRvdWLm/LCZDahYiPd7LYHUunehNioY8DMfQz4AFD5
vUYwlZGCUyzpu6yIcEtKaJQxU31xIRNzHlB1k7S4XtSvOFr8XtxS8lZLLeLuBrwndiJ35GrMb1f5
MBGSwZPaIDrDZRIMT0jOrdNebvUEcjqIW/QsovKg+Ky5EEozChASPFyXrwKIi8Xm+1AX49WZV37p
vGnzzTP0TyguPtQnUrIiQSxoYS1+IVwUx787x7YTdPDomNifk6yTOcjyka1sxTVhyduUCm5/pRaX
dLijZCBTNVHoTAC+TmotmBuicnQW59DHIR6eECW3VeYBwJ9UTDovZCkc0XzDIf9Q+q5fUkbHN6q2
QGrFzFedW0QQg91H7TE4h8DIQU4AQOGe1Z2j7znTOmnayamP4CxviYy2yyiKCItvkTFOwxMImN2b
X5PKKQal3ZDTIrKJ4y4I0DEEbm1iteLmi9Ds9oDVXMeRudKbiLPM4oa+sxQL9wJ1j+IsMIP8wDNY
vlapNF1f/KkqGNETNtdZkvJ/QcscrZwyQAdaCyABhhHnlR5WypyRkYLuuTWAm4mfg4hSx22/d9Un
jxiYeIxCUir7+piT7rNFvU9FfiNlSE05TkX857GPPcxH1Fm3iEEvINQVuFnvH+M3yTrr/0TZro2L
autwfMt7OQvp70aOJ70UFG6p61g1cprNXfD8WGr9CryJMrokW7u4upqLaHz//JdmXFtaDMlS0Imy
CfaEN1d3Lz7pAiiRvrvDQLWHKBttV8lWBilGq42gH92vueprIqUKbKU4DpeKrermwhC5ZR2YbdRN
0E2sO0fpaHGGFa7R6yQhnHaqKhzjzFLBHpqGhztG9QyTV5+veSAsTLN/W4q8smrmKNEdDWgMUEcY
yJFOtfmlp60+rXkhtiS3gzyP1vnMVuwxDZbHUjYLlG9JfrCa1nF4KJfPbTtIEKEwBg2M+lwQjGhC
TuAIvA/lwwQZ2Ivh8GPSASYDY/TzrNU2u077D5oJdY0MX6BbH4iU7gfdE8N2jZmiXuEkrRjM06Me
hUgi3ADAD+gGFIjNCEaYB17pa6gOA8YhybXFxLEtaYI0tSnAYPkTG8AEvZdZHfxhVVQ9I129g0F0
Qo7VKmmrf0tdtdw51dgMimIBIF/x8AkoVhC0994Td7zyvEwbrnu/vOwD/8QBZj0CM5B7s0KCuTbM
z1zZ749qb38tU01IAdWbC6xwaqqndaouLLkszDrZqxcATye6JLr+DkWp9Ap9d168Ims/PkAzynwj
H2oiDhjLswAFZqnLc/IQIol6OwkcpZLfhv9adOYM8l9JUUTL6/743UqXDUFe4Rl/EKkVwHE6zISM
tAKocTu75Mg2W260wYjxhTYT1Jtjp6ef+B0c/rL+pdxmU2Pwpi6J0WrKjLHya1lWDHs53DOcP+rK
B/8HkQ0/dRvL5sNZq/45G5F0GY0iTr5qgGgfkd2OxpBTZ4pC0zao3wvelzrQPv2vU5gE403RVCns
xLcMJsuHEcTp0je1Br86WDIx6oP30G/+9jVSMb21SViRrzJ7LlnzBa3ZY2v93ZSxdbCab5fUYW96
6Aj+A/trD42MR2SQaLccIuHiccxOQv63ouYXxyT9WenM9/FHRCvZNpPWpDB6iFDPsWnfoV+aDOhq
hc3jNIWn1vSESuUXYo+bE8cBx3UpXhIG36MtFi9DNdP6i99USLIcyiphkc5eRPch1CyBl62M+Xba
0mysvjN6+9Iw1LVN+t+nEkVTAPsIhmj94hL3em6UgxYijUeUevyHPoX6R9vPS5NGKshJFLwRqoIs
001+bPoHRJlMo6XXztcPZn/6YslNXaTzxOzb6sGNdW+fJq/4zJ1BB7Fo0ri/NP3wjHFDHjkEE9Hr
iVsB8kLHxkptSRdYfQCmPwMYZdi4rctrQDGjxzrmp4Q2shNrf1gmqCkZ+wYCtq36U33vvQ7E1MPl
PV/7OFDuOz7rvv/uDMSkhEkZKFPBktVRJnajRO/DikLeaBEzVzPDc6TjcxvW/uSby5HNVgU7myRW
D1P6GBahk6Yt1jtDPoPlP7Dm6HQXjISKU9aJ1uqcemoK/tFJrKswB2BCoCaDQM79G51iWBnIjOeI
U83C1UOyW4XQEpSCaafUNd1JS/9WFlI0ormYrQnOKHIdcL9FK1nqFF4r8kjh9ToOtZ/pMPL7jCDw
DTtFBjfMA3Tg37Hmsnq9euVGhsQmXrJ6IdAJSFPHQyMt8Ix7HGhE4RnIqe0TzlU7SZsgT2vIQ+ae
VKVJB1aaj+PyY1SvhT8AANTtRAPVOl4l9wPnDdeg+0neQMxjZZ4x4BLdv1bsUOLB830umw5UTO9E
YfMNgM22oLbJ62pO3KjACFps/xFQoigGZ41bjsJ9qTu7+nz9OWJqIXuJTp9H998vyr/VpwexzwxK
KJQDXfGHn8mJrWSM6Tb1ce62dxaRC9tpFTC0lvLoS5zxuwqwsX7s0ullWXPDFI/RqoIWBsVly1q1
LDNGAx56JOm9xeSB0eP9xmnMvFB6IcDjfQRCrkATDRepFYian2W3AadP0tc2Hsa2frnfRFdUCVb+
0jcFLd4jKH0AcbH/C9U0ofhkSwGxkF3QuSpmZE8Wv8GfQV7uznWbKchTCtkX7NICDjhAaglWuCn0
YqLh3CpUO++S3OxuVDuoF5iNVyKVYd1ABrOdJrcr+t3L2vmMENB8LQ7hwZxyJEFGbUSmrXHzcBZ6
iPa5M+aLc32PTYyJb6/Tavc89MuEbzxv/Hp6tAD6NciUlcwAZ/AvJkGxH9TjuStWd0qTVfh15Fbw
wLVEBqBw6NfZS8CPlNm6AsFRUHm82e1SduMcR8E4SfH1KSdYzG3RGmb7UYGA0MixxK2HCzeS3Nk0
y8/syHEW80uZFm4WWXXV21rlKD7UgYUgOte/YL2wKnxGXuAXcXdsOZT25xG7lpyiknS8xPfuecAb
gIGMc4TYxR1e0/Tf7hTmLtYbeyUw2XYqhuBMus9IDq0F1/3kwUikXGArW9EZQKm1f2UH6m7K+/Sr
V2J4ohY6K+oA47P+fZOY1JsbO4omjlMOzkgTdirQ+kY4msUqgJvo3HyNzqA5WMnRKCnTtuOd5Euq
wK5ZXvizoVsIlfd2GdJLsea+OaMo9s9ycpcAcArcT/zb7VnxuRpA/36glWQyK0BTrFz4KZ6jhcJI
AuZ/GxL2ebJSh17iEM7D3AuFaJFSrlUQ/W/rn0Qlv7nLjvPaDa89/cZVwCqwv406OQ6fmyltXEKF
iaht1P65Kz9nL5k83ilmEuTrmEIaJKcOfs2rtTwsPCffZj/OI18nQXX2INT06r/qw2G64FVMPusK
XM2Y+fB5SLD3r2AkcLfvAJ1eJhuseI8xaiaHD6X37OInK99JxOPQL1JUkLTbDAQG6E1grNknELu3
4sOmUWk83oOu/Bbt/eftScWx/deQSJwZ4qsmUOZepUL5h/p+ftPZ67vEHla8iMUSwYRE2LubVEQL
1a2JgqzLDNmj415/tP3gJ/h5jywXE6FgRcHIvzNSQE+CODzqGEeQGxsW5LZXlYK1sGd120i3LuGW
6HPAqYs7TAETNkQeYudnTqvkjLctw6E9jxomWExsamIQVo02r2ybp1mdBN5TuOZYNF+3dWgfnrDY
tyPqOOJDmF578WQTWbiMAO32AOstS/ia+natqnUpIaxFt7O9odnQcJUrMsQnJRJ0N11jRFtpdd2o
VcGYpTmUjAKQP8AI65w6iPNSiXEj5wzc7KznammUlcs7VxEIRNoGZ8sbXTPEvsmNTOUrTiuq6R2e
2mkZkyMqVn9OGvj2w8nMdK6BAGS2PE1Ti28rc+1spHdowSsjM3vvX6arlw5Elm5J9p7A0alvaV2W
b/r93kytyaiKnOuBvTgbKgikoHWPCMSNHAP68Fm11khR1ZjlIoOfuoLAIKQiMLY2Sjv3SWbD9jvS
iOo5IZwOjdOqjMRzrbmy28HWXhVpMEYG7bIawhudCTfQQRk7Yg19Rp54y4yHXSDRUl8WPE/IQeYx
RiJP7hQCHdMHv2TQtg4S147+zSOAWheSa1lrzE9tFtmr8FgJRtvxYtFACmkXwkdlNj+ipwS/X29q
cffS5TdZkSyyWSKjvF2dvyzTCGcOaZLk1rbJuYi0DHun1E0fxCpazMa0QTGvSv7IBoILPZQZrRSW
Toem9/lyRcunu8dvirqfXvFskyq1vO7f5WIVLRYd6I0/puJ8K7iKdPmXKfLgXgd1FjM/hSVPRazR
ACgVLn6HsNO498v4NEb+EfgaC4Z1SfBEjNvcfenrD79w4Z5rBUX7Ni3AKPowwdmCiWFZRMHOMoyb
0YQgwZIldK9VMxonrxY8Fj5t18FyWQkSWiQyTDRvGya5v5r/fPi80mmf++iykzhDijJ1vr38by23
ie+8JzKRxWPcIsTxtZuCYjqVM+JgSjVyOPXR7C9/gwRI45UYWbqmzgIy42GUMT9SQMPZHK0PNo3B
A38mYAQ4DgplKgLXxO+HLT4hTIbJnBw0oM0fnBxJXAB5VMi3rFfyFjw2gSzo5W/wK5ek//yOkjkw
tuP5KOr4x/zHuD1/9Kp24rWsyx6TEixdakJDX7R9EgqE72Yrv2rwS5QArtlQy3/lA+1eZa2OD1Yd
FaDGLUq8aoQZq9zOunX6jNGXK2VkqabTzWGLhnCFlQXY3vX64QeN+lVwbDXzWb+s4bsvvVMjoBv/
iZu5ZwPLR9L+lQqBlUrhPrbQjd3QhBKSJhYzXMNkahTqKG7YoGt0j/AnJfSACjxUKRC63IOOVqBB
kw5lG4omZ1yW5yy+XWMzC6lwNaSsm9vH78Qg36DUbFb+49SD5Yx/IpWnGvSk6CjuXX5UxFVQgJmQ
osiER8N9NLrnF5ime6XdB1/HmXOOBe2+Nwqj3pe37qbHLFOTP60kYzYCWWVWYR+OA5g0fX3j8c9y
RALjDebAmKdVH5dnlYE0q4uEOwtg9FwfEt5hgwgimiPErWqoWIMYEP7LVgQuX03JCtq5aCgKHN/9
sVH8N+0rnENqIlgYaWiBOU2CeJgloCJ5G2YHSulCB0aWBKycxtMnA/5kIDVkjPrEXz4NTtbskKle
9dDVjCL2CQVMeOZXYrG26qs9meAsngfgpFG0Q8lS8c5jsb07EQZ13b2BElyms/k6DdDRgTjaIggQ
Dew7oJB/OXshUtwYVovAGvv2W1UbNIVw8LFSUNWJsZ781y54flbiacqM/9I80Sireq0N5Om8NOqu
NNeU7lRBMFM8NGnfwELyfF0juJE4YaxNebpXfKAHgEKXCyPdUH4JIUHT9Y2DZ6Nyq7YC3sYR4C0v
jDZjYIGhaN2FTfjicAfqdFQcs85P4AKSOOlBU+hEvh/nDPcm1RFM7mPe5ezvT7dNtQNRe1vPM/a2
4I0aaomqeJIo+wZmMgA/Ne1o+jX/R2uu6p86tYEsBPbzgv2+VPsUNtDzgTiQfK8kQijtoDzGlakl
qH3vY2dIC+xv2++mANSgF60FH8vY5rMF5kqmauKUt4Lp3QRtrKHnCjlF+Rkt1DRe9wHR6w4eb+Oa
10ML3q3I38TZmwCa7WrCwBrvqI22TMYgCUGJUNEXVjZUhXJB0jBUMPBwOAp4/DW3HgpfBjx8foD5
LScqzReBxBAra9FBndcWH6m0Y4fed4jIyks2sPAWKcucjBrdKjayM7jY+UA0Vp3GFQIpd/mxqlvF
Etr2SRzV5aPuawf2CO16OIlY4tnEt0dbl1/jFipqbENmihb0JKPz2UskVUTU65K6vC3EcrzZ4T/E
SYbsj20d4he7bw1zLn62lmi1iVOI9Zh9pmeLVK9xYLzUDXr1R5EoSswM7v0qR/RlY4CKytYydwD/
f1bQRI4HBugUBkAlmLbCDribvCmaj/L09LyFX2agTfDhO8bqSWgiAzBuy5m3zdVGHzhnA0M9bT6o
IyCPacy5sbxoSoPlFsK27Z94BY3n0WtztOPU536l3xuxtfv6QCgERcTGxM1VetAj+LHx0wXGbZvn
Y4f1H++kNi/imSnDQdlyldqaIvrx7MGQrFq1Pn9WIVr7WheEEcom24WfDtMYiab9vJGG223JGrwn
SdWGAPD4ZJmrr2o4FTSueX4GMx+MtQKmfDed6TsPFMU4cSt0yIU6gsa6v1/htF00y7WfJdAnj0HS
aohavKxMK5XL0vHN8+2h5CcT8rEceblfYef40EHTI6sZ7x+eSi70+c8BuamBMAysyrKFHdCl9k+i
6O5tI2tPXpYb/dqWSVWlP98nC54DBfkNtjMmz/oM087BssitlllSuVR2ZISjdLbYHfPTFDT8KT9S
0f6q0QRr6TVN8BNdbwLBu2XqjwoAHLw8aS5qODmSAM7escMNC8LIeq7JcDuZmVQbNrT+F4ba7WU0
mHPkdw3eDI8zSrXmjAGJ1qntGCpDDAyW4fXSenVlUWNMAqds0MVC4/BlVnsTvJYwMJ36bTcyG4s/
Bhahz/UfY44SACNEfEf22x1QqHfnswXpKPEuZzpwPBpw4sEPmI+7wh7Hz0mNwqAB9eE0lGaqysFl
tMXQ8Dj4zSrn4UhlTjWSwVN37lg6ffOr0GcMzdysmMoE8PqLV7/D5PGvCDQ9Sw46EYIjde1wwea5
DZrWMxTZIIAy+Wxe8VTKORjl+qQlcZUf9il6Afwn4SlZbqfkq7x2nOZN+EZUWZLa1jOg0zyaKfbc
JzmqbKIABUICkti2TtyNiKxm1SaLj3W5/622WpnHyPT0AH2GtSoqroLUFTk4ZNuZNLXfQdiZfP7g
+aMtl+9doPaMkK98Kq4UmUEvliGvfCp8Xk2KYtMY+PDriRHCKH28SUlpNPuvjVbX9ShOmI7DzJtQ
mXEns3LtRJCD21VrWYE9Z/ZWLuJAu82DwpC5jYhmcM7/LbaD3dJ7Xj4cS/kHQ9MPb1DvNVzrQsgH
9HGPI0xVv5D3DWovYo/rwda/oOMuXlAWY2FKxXkAUussjkbfCj9YWwboC0IoI0fA2rEWqWAX7kep
tp5RIRH6LEljyKZdMqtaUQp5JYNQmMnduS4kuZ+qzbYWXLkDFlG+NFTnf+VZIEl1XY+IpESEkZ/o
tOkWOhOL1UthTOavuPo82YKTLB2M1L3IkZ/mHEqIZ6ipW3iTshoYPpAXGUMabp4bMLH89FJ+iHg9
x1LxBUMB5uoT74v+go8JVTuBqUyCkLpQk5BU+OxHIxDjDxesT7jz+sVFTijP1rI6xEZDTKmwXRlD
jVtcDN8o0u28kyCuDQgEr3+69YHIRjRN6Xd2yTXmBB1+izDtwaKjZF7ARuv5v8TDylABcPbzT7pN
TAkvgGMoO2cb5JgW/ir4u67K0uMo7FdgWmuVg8qcY3hGJYO0+/fnfDBgoZnxp9kAeaWEOUnav6z9
okoReUsbi+tlYbGIFSrLzhc3k3dzLOWCknLeMjNHNjGL0G051X7FC/Ds0ulrFvpeTSwz7jEX2/ZZ
5Yo8r/kiqunFW0ft2zEsoH5URQYFN7dFZAWAjwlNnNRnHe6AVUTx1HcIRTeMwmargrsupU0NGLMJ
S3EEpj//ybWiIZhyIAUE6IqWIDEQ7yGeKeAlfeaJMxc8LZ7Vwb3QeWNQl/s4LpDTtE/ke8kPhvHC
USYK/OoKt18yElz/+DFbmRc0VFPFEb5++QdCkogOglWuGAiwy7lhZ4SahEKlyuj1tIpytef6dmk2
9SX7qOO8rMREhh8mkk4NkQzC5ZjUGHkWwzltTM0bCxStH/YApRonBx0w3xA9MTjuoY3NIfw2+sg/
laGDBmfSiLijqQ441fBsHj1CWnmI3Fgtf1wSoUnpAXcFmzb3TzrmbD+IpBvHzrXgylA5/ER5yVWU
nvGD7wEYQ7Dyte+MCJQfDIyLpeg5CuzcIZFGbySc8KFdQ0iQhDa3ThC5Oljgsprsxbxjw/XDOriB
t3EAtNb1CSIBpBDkdzJoXlu20znekQXrkrVlMShoMDjJcApR1d2FugPhnSuEUFwQdsX9/SvlBt7H
B9sUx78wN6f+iIOdjzSqNzA9nmKtXX1FHYTvnzXFSFIT2/TA0183xkroe1UdaP+2iwKfVgWIef/h
8IF7WOEWKdYfa8wNRhu51YcspUacDpUGj85EJpJfHaORp2RC9Siv7l43+Z7gkHkG/k7SGsDWieNF
odenBOUzqC2s1SRFMKVfPhHTWDR24SzotoEo/mqJNTd/ifHIH5fU20c3Z3L08A/VZhVJxkYeweSk
UdpZc19QW/4GPiAjevfiwpmkzzSVPhA8wAiynCV9OXGdFXKOiFNdQj5/c/Jfz7u4wGVE1ECD0P3w
xIctLPms0xrdFzFoQGg2KF66W0biG1eFqliwNR9NJs8bVXIgabHWX8UaYvdkvqYAWPLsknUQ8Kcz
/d6w3Lqd/0x1g+UB8a9OYhnEC+lodFG3FarNqYvSqEr8/IITbSmWBtDN45jhEGgPdG+jB9AsXBXv
Qlq1zxMWCv6GWF/BBpyzxDd5YVaLmrqfEnSUvPlnuGmQhD3JQsKBycu8GaJUnBi2GGrS3I66vITB
4DQWhrdt7IVEYLDXKHk0oHs9O7NEDJCuOLptBt9cj4IJrDHF3RoCQDspmfGEKBuF/Ii7+FUAQCFz
a91l7XIJ9zhPH+sU4UvC6W27d4ZjnsXY0pAYvIlSA6SDuX9tXlgsrjSZcgzvI4g9uL/xyy/GCSvY
uzh7N7Isy6m0uNvrwAfO1l+uc99czri7m2AO28fJgSGzKMVPKjisW1638hMLEor14SyRxzclRM56
0gHCE4Qn862ukbJ1D7KqSTPBGH4QMRry0dhGgvKtbzgP02TzFwQJDdwptGMijag9GUmlAmHGUDtz
3uPhwosV67A3aN7S7umVmdEP/RjrCn+hjS+3tYQ2W/depm47LF5/QDraqNX9154M7Y2wXV7VIehg
pxr9eLDE8qssgLwxJEQ8TNeian8QqOYHrfpbqhBKozkE8EDU6Zc+bPdVT1URqaTVbuJHeGP0nE6Z
vulaN84Vdkpa86ySlleIM9Q6hUOVHb3j8G4bO2kvWdsZg+/ltRNGRUA17JgZCX1S0FMWLKEQSOhB
l83Sshp52GR371Dbj2QMsui+o6Ow64z0PCyYKv7Kqp3sRnMAXyqdz24y9EvbE9tYOFgJlr6m+tHM
V0O+/vTU7miWSNzz3IVDewbuuzv7+6sXuvdX9oI24jdtW/8oqGojYqglp6GFBJFAJrnGNnjjcOhc
8m3WiF+yCPZkQisK/CPzN2ZBHbhmANeZNYPra0LPz2OZlo0JOQJ2zQc8+BOVx3jLl6Ng1wDDA2xq
PbWl5+HbK7+54J4qbLe0WvDUaSu2ZHU7slIPRko8s6qxF/Pj7py0mSFkUrhfubr9rW3gn8Ow9HaL
BuUrpLtctog1p9PjmDeDpp+t5uDQHgupgM2K9aRS6g9ylelnKKhV03U5TgymUeaKjd8bleDyNhH1
pbrUaui88IPAxrpHL92hpioxazwLYekLUBdbPYp9i8NDur7bmqlEfEpZjBve4ezJpb3aXN64pISg
WACG+zhWMLYbusjMBwiMzJAfuJqG30aRJE8Ik7abUTjDYwhml5yond6MRGUPi28gmedLzm5bakUe
Zp+0a8FsSce9aSDhfvUKmyuUFIbRhvSeTrWM+rMvnGNFKq3SsHULVdtcGs94JU+vaj7l+zRW5mvD
3yqJaAIHvLI6FIjBVT9jBXGCGx6qtqDlWz6VS6e2t0uJXrM5iAmqkEHPlsLmfSd65uSYVCOYpLxe
7EFA0D3cWgIe+WX2ZvUTD1ibTe2NW+wKdWmbIP2CnjREo881JEmT/GzWoIMDMwd3ySbRBbTWa9p6
Rw3nj8LpNAxEtI2z0gl5L9gdBLqtGh22s6H9frTCjkG7sh4VhPe40EmalnaiqoABgHLkKfGJ9dFq
LteoA4MSmiZKDLIeWcu8/+2YUak04meLM/c101zfxaX1GBpt9Wd+8wirTwqMGh73WcnaMkw0Zi/g
Fw9oGuX0yEXtBBFDyBToj2iqGEc+nnCFDHiS+bt1Qf6blPjlmKslcz2b4N1+pD80RLb2Kb+GLcRj
z61k5xLwGZS+4A6dVXqBU6x0seVLbH5itTio90KGSy2/rxWTYzQJ3yE5lWBoXgsOi0HtINopXEN6
azoc7CLOL7jkIWoW9klDbp4TFeDpihP55Mbrz8Jy0QF/xbm62AYGrVIoWZjXjF4fwFCDQuYjeJ6h
5SeelR3elqbIX6tClJCg/vI0smrsNSeXh3jJs6j8JuZQ0pkIzwlgtRWJq8VajMih1d6VpB9o7NwR
3HECA80slBqqGldXrgTJ+6EAZ2QEHAtfvKIrVPcDadxWvZz9u36GB6jK2zq8gQu6ByxW41U54kvx
MHJYl0Pxat4C0d8VHQ8QVszhA+AMVwbVgabEiakkxeEJfng7m1/VpWL4du/8j2q6U2bA3IqJNpnQ
m2XcK+f65L2zwEKRhlL+JXExE0HWzAs6rB8aN6hkS0vrcg6IKcSTUdec3b925ZzfxsfRuctCsvbk
/4sQNRwMEnMT8awR+0C2v3nrZhmx8RNlBtBLpyl8/Da8ORISJC82Ye6lrmb4Zpr3bEFK9LXfzS2D
bxdBISUOcU+9x+GYEDr29+7ReQ2NnBVrZscdUz+axCtWXz3S2tTQt2SFfi7twb4J0Iu1dE3b+Azv
xk9K2v8WsARQ+Nvyh9tEw0sg7uewMdbqYmleoAHiZFA9MPRxN3QHxKMwoPtT7cPEWKrkynxei/Si
2KPZkA4PBWvH7lM0EpJmIKmg9aM9bQiA2VKxzH2DUAG4f9PuPJpEMGMDcrUyuFXsYlKDXQ7qOfvp
8QX5yvDsowQu3i9MlDdldrORmchBQMeXUEHfxqqCbQj1LRu/x/U9DHXmWLqeJ5IFZYmIYRcJRlW/
17EjOPmRncWH5rafV+7IOZarSIM8zyUUNhQkevKY/3T1tozAmIr12UQ+0hk5y3zS5KliMcVGQOtW
itnkSZv0y1eMtxJqmhiDijsbElfWJM0i5VmTV8JwcFT0riXt2ZbWHlOXDAzWSQn/BqrVi2ADRsN6
fyLlr/RDnYL0yaPuG68uIRT5FIOst9iN66J4tgEe2/0tqMHf8Ow8bEH18Fa0OPlo/33flgBrNdE7
+o/LUEtmGPqWxxbbvDBVIWRSZmtbNmHqgC0uwaAVY76Jg3dTR53EbqaLNbFyXuAnZK+KHfX2C3Eg
7ls9CEODGHtQHeL1uWa7hf3drgqa+r9bCjI/flsKUKG1qPdTZaUQLTRdRqWgIdqdeBLwQi03jx5H
ZgGlhago/OP6joz3TkzaFcI7iqk6cZZ2E0RZ/YqPF/mvoYCJq7Le/1pJq/drkWvBD/RAEgKbvXp5
3xpCQ+/AfT1JtP0mPGZKVdEASPtoeIHmT9ybqiG9IP7kZSEmqcGvXK7v2w+BDrlymsX+h81jswZz
+ELsBBCWO7g1eimuMhs1ns2rQZP9TFTZuaTZQ0jUTMDNvYQuCMISjOdvsC9FdQd8ihaYoydN0MG5
VH/854SLFPy6dg7tGU8C8w8OujM2H8FT9VsQE5fVEAxooHTm4XiYJWk/opQ9PiRKbQLSfDgwlAYT
pXLVTQEDNQmQhsxtfpB3/3Pj4GBV5hSe//4lRs3pBy01vBh739IAhWXW1xGuwF5y1CVSVwH/hYYj
60mQIr13nL6vpTZ25Sj1ktzXSdxyrizyC9QfQ7S7jc4EWcGAO8ifiMEWhwnH8kUsrTKGzhB+qim1
l8ow8HGFcIdTdEqZKIc9c+fUJZwXpyfSl6M0mEyuzmA9lhaEEFclMNftzqsYRYWeBKD9YBUyS7Md
Xc6yYV92QPuKMgyZQS5J4xs4R3AKLologrs8JJFNr5p0XVdzThXObG3h7oKJp1PGrDJINwzjyoDP
UnFQtd9eQjOnAI2A6xnbq8Nfx6lIex2NavS85NxUfDTIWtNZVvitign1GbpMPSnuKOCbgCEhXHJZ
tDzY/rLlAKmdSH5fZS+7epR9FQrod2NgH1I4I42eNVvvbt+YpqrEG2R+iz/+GhKaElg3Nn9pmkz4
XhxJbS5GNujGUgtT5WXMbC14FQCtbR86HwYCsxvBkIjhYZ8ZwhU5A7IQLS7rukKoMHXakR3pJ53A
ENnFWAvksBBNGVBEuJP2d9RpYEdMmBEhC9VHRLggy+3XZ+4xHCCeYd7zUFrdPvE276evWDG0lHNl
DqlViTX7wJShv8/OdrxrD5ZcjfxRLadHitev+OrkuLDSP2F/GwaONz9VO999UoDwCYnu+bExx1jf
Eiz+nzB4Ny6Chtx8t1HCewGX+Uq72tNRBjVXkU4SUBzdPJS9fRpjZSabInsDCEV8zP3MlaBkVUOz
saa863lSfDVg6tXMdWWNzvK8KoY5kJ26MOjSMJ1Cs0ScdjqO+X3czkaxY6mjAxnnpgDWs6jHE6VZ
MqhbOdlUr+683LGj8wYOYTSEVYuyLZD2opysdfyRtcDSlwj6Q8vgv9Xlk67QyhU63M41zLfyO5cB
/V8Lnq3fSRK9gH13L79G5k6lWrXU/sTiRhCjnU3wLMqnFyDoMX/rLAjDy7howHQfOVCt+3Z3IDc4
aQFSSmWRr2Xd4xRQlZJRuF+jh5BTk/QVIgDk5Phd3jCnuooxFkbTxS8uQDoAjv6CYHzBHaVYfSHa
NOabuxXx3O/Ey60bQjpAr3KkOta3CyLaq3FIuhC4Uy9BPoPRxp0Sts6j5+LUOaSYJYUAUeOlk7Nt
9ENlNp71nwGuaN39Cv8Vokt0McbpG+q3Uv3nxQcbDWRu0TYzdbTVufbX4KP8UyguW6Rnckz1HXRn
hAoNuBbIGBhLX1z+HiJuX+R5igGJDaDeYCH7xeFQLasva/zmgo8mTgDbAoj2I9X/cPgN0NpFA9oh
KclY5tyOO6PkSX7bV9GAOKeNke4ISQh2YS2ers/QwNYFP1zDQ1g9lIJeMh06VEoCVO8dP7p3KLqk
tPiRgIoXaQMdTQSEvXVVgYYY5ZhjiP3eLWq0CJ2Ph6p2GMmmqmCO/qlhEhcpcwPSgeyUiKW4ztNp
Et73vT+EQrLXZXhFhbRM9dl+ei+9W9oXQagkAKa4bKamJ2CE8TeQzkt6wa3t2HWPnDi2vE/uExSm
2vQY4z5klaTTq6pL4n43P/xYFUcg+ISjUW91H+IsVt7uvXuGkAcGJ596XIPkizE74Y8Azh8frDtx
yxsZyVB5CTS6T2DhQKOJBsQnXi6CghltRmbnoSj3vFQ7jSNs8T3iMjcCMljK2KLfF+MtpptsALKe
fyM8OXHzUIjomByDcSUDOAk2pr5q6YL0WO5K004TA89D0vw9vbOm8mgiXKdVQ51hpk3BL5pFgIGk
oFWmkqsaxtmOnUcOlUtPPW0UTj8UW+sxUng6FnovqqkTd46Dr1mP3aJRhWLUQU/XESj8FgmV0EkL
d9yLGLQGjCZD4mmPbElDQpPpY7UPzeTZ5Jp8AMbCHurur3/uvyWxKk2khLKYkgujzmnJyWbQcIm3
qnMYA8xN9yebGA16TUjQ+Swjx7q1MZ940644Et3YasvHlq6qzm4vm+DLoSd8PxenvfwPtu99Y12a
e5YTu4SuUJQc3lZyYTHrtOP/sXuX/KwIyidX0+0+e349rAi8GlB23XzgN/b8L5b/kwZB11/J7jFc
W54xiq1KugkfpchUvXyKu3j3u41/JIB/pc7Hw4kwMy4vZtcOGFn4RlGaa3hZzBL2/wgALyfx1O/Y
fSB1ZDAGeMXGvbp0TC9MKrdUB0h5HcDGwh+uLm+QBWekoq4mxOdiFuhxj88wWHkalqq/C2SM9qbK
xJXufLsRUMj/xS4+hkU1Ri7OGk0okDIw8+Px3X3uDiC3gAJWTqaR9emrnFKRImI/n86CzzI6Qs6k
Z+5bT1nOt/l+02ALbTbFvaNbFwnKCTcXM+bbjAte5bBya9SsVvf8HdPAwLIX9V8VDhQnc/+6WYKS
BFpDuIzXJ3XiuyQdTg+F37WoYXgZ7m0dAy25Iy+5qbNTrXyvgtPgcqJbHQLxp9jPuopZs4E+tps5
ZItMF+kHewdrrUqCPkGA+QiIx3SLOdl1MS4G0fbJvsIkNhNsELt6Cr7AvDko06mICKV9HS5MUHAi
tLPbo2t80yfH+BaNlrW6yVUpkJYnZHzAN4JU7/2P9qjP1t2aUdzujn2XTn9UGaPht3eJnXHrcr0J
IxHqCAYlk2ux3w4hB+c6y0xIWKiv0EQwoeqxZQ9iz6JHBqw0YVYVL8BvdX1WUxgs5/JDjkEzi47T
0080X5TZNSZbRCQJz3xS7kqjvp+C9wdwrtU9kLIiCUqebc/a/ZneoTaFGO3dL5rrGHW98JwsycPB
fxe+SqlyEUTFkVbsT2vmx5jxuF+awUiLQ6VLiB52GHIXTz7B9nPtQBSwQ1GsE81p1VEQdTC4SiWU
UGnHArg9rWF/fQ5cjbaeRknO0aq0Qzt8n05OfPvyJd8cDzShF1eJz58MGxd9G1qZqVNP2KTKOvlp
dXE3ePMblTrz+h3tdIMKY/UTW8wrSDfY0k8rUbqr06tX41E+WACbIGoOPlk8SJO+VHY2eIlAJOYw
bJQu1+B+bisesaRB0tMGyGsfnxbxl4nybgfTVi5HVRXppNFUAIME7PjsPqWvOq8IbE25WpqPyQXo
Sz/gjHADxFU6svRsGVqGLDtWXZSbX7Cjnt6mgbF5yRS5wNsDkKlmdRpcw/JyS7gk1lZIidT+8lZ2
emIb8jrhqVIlbVBQVulLTaNTq/FzFMyCzyon2vZaKhgBgroYg3500P79qGjHH99e1pt/esCZcrr3
KU4qSx+tU/zfbHShLMdto9OXGCQkOx20gqABoQa12C98y+VIdQ3cuh5lEpkTIep7O9opVeJInK6B
Kv39uvJPB5wIBenh2FkcnvxpJ977evWkneu+fmwE3RSgKptS5yq0Lb7wy2w5XBuJcBazEzU9jt8E
fg21mME5ZZEap/fJe/Kpwz3DaEcMvkqOw/8DbqHtNciYLI002jAJvRdb+37BNqT9G3Aq8K4yKuYh
Z5GYBeZjvVfr4pDHYhicWjptL0Icq9MBwCuEHkfTA3fI5YMyGSvnbpB8vca6PJoM5ioMJ3Dk1OS6
8poeKqbP4ACn7fRyQeN3Lq+QMG4SpQcK0KbTQ40P2dW7YQRQ3EGP0tzJDWxNdiDCzEgSwlLEnoFk
6c1ilORc1ohu+0s4HKQFR7Bvsy+X7mUshjbjGqaaL0DVxe5M9+mc1Z9Nw/+9tSaJ4A42fPFiwIhd
+0xTbcgrDAFvzlA3muAGXlXKBl5kH7FuufxPdDuC4t5blGUkBtJQhfYE+T5ZGHKG0cBp9nfZP7+i
OS4VzmEC1aHj+/tzvZMQlcXvAZCluhMwCYWTn+NvWfS1k5AfHBvTTMLhMKc1UBDF4g/PcQluzU5/
6jBDs17g87MBTKn7hwwhy4CLdCLaskprWy84AhKQzlV/aLVLz0h7oRHbY8py1o+0q9ISz+9vXSE3
/mXzoGfMhOj9hJ9AgHlRLW3glFWsPOirlg63meH+ssD5joVsUkXkZ4I57kvEGcnr5/zNwP/1pZXs
ZlEVqRkNH8yGT1jrQcDnlOLSzpjEZKz6yrwQYwKB2bSnMH31e8/58ACMvFtNF1+8wQjvZf8XBexJ
y5NMu+sm2qQM3a4KX48DVaXtsSNcU+q0MFu//nMBZXRxKGCAcKvRjIO0OJdbJbA7a8rT+uBxc9AO
WPpxrqGvVeAhaRRPnLXCMxPRrzEb90EZVBVd3s5voLXwNKrUnCPyUMMN8KO7a+n24gSlvu/LjC3n
/+kXw/UfnDcDdWOP1WX5f9rwMJVS6zpAW+5im9dtfx3McPl9dgXAw5Zd5PwEziMjel+UDOUWHQGN
5ksrvpIW7LvHyPpauaK7AMeu3l2hrigoRzJniItcPkv73xkJMTmBIpaQfGZaJwyRSdU3pH20n3xW
GPjEYGGdqTYKG6nSxDTDFYN6ptC02uo85r1gB4Ns/F7gwXPbqeFhw0Cj3oR/TlvgT4mE7RaDoqdY
upFhsikTQKg87fUF27ss8Xpxzv2tQpMOD+fvpguAVtaiYt8du/kr9vnmc1wjDE+TBr2a6ezv4zDN
jcOZ1Tn0iidG0KMhuO8CrmUNt4h5u+zgt9HD5ORANUWDBELzU1qiFxt7BlBwBy4n+P3Jv+Xoa2i7
G702Eobk58rnijuKwpa9C86gh/HWAqrwqiCrZtM8vcGPEDs+Ayn2NAa+mnCLp70d0SmQoFK0QDq6
CVvkf8KPmnTH+C91HMjtjCisNzwlGI+S9Yd0f20L9eFD7FVnWrc59mZnnBuy3suy3ZVs1kgGlFPS
K6hw2lK5swzuF+WRiknAO3G7CmUhGGYQqngQk+gIQk+FmhMulN9Awb1so5pVz8lmuOno4s0XooN/
4/TnY5s1x1BgVOeo/ZZ7yK1tKJiUUdUvjxzcExGte803CyUGlszpVv5bzYV42Q+CEgHGyUYRF5tJ
Swl27MPOlxbiROT5ewjgDQdujUw4mR10b1cJsqjCONEieg7vF0NOQ863C/K3PUE5ygBfSsR73VRo
QETF5hxYf1z3m0WN4sMMulUfOp39YSF8i1LA+YiMcH/MDWwfRD5yYPkiEe3KnJfZ0owCaNpDePYf
w0WNkd+/8GXk2u3RnIe96Ltlp0daLLUOxctxO/DZBWEJWbUezKsUM1eyrMB23P9bL5pvi3Y9a8y5
Ig7dMuTW1ph+pG3DkZFx1irLgzzKN/Db/DBEc/RL3vvuVBuExA/z6nba/zr+D4lL5QZPmjC8/+k1
Lp3zgmSNS6yFP0T/PIsVndCoiAee8vYlzErZWQhq92r3Wwr94RMIXE47Ebuh7ESncZ3zMng1eh3L
ZX8WRu4Hb3XMch84yaKBEElPoMtg/1LgepCLcCRMVgAhi7zWwexLRusKvjdCGVHQaAhk/wLRHAms
BCy+VbWsa5SyPZPGm7GNKTZ+XcoWRBCaZZUSOtTd15Y2ZjOiKFFpWfjMuKhEcVEp9TzxgRb3lTLS
oIQeRvt/vSUa99klxaFCOZ4v70JagQM/uTXIwnq8zUy/q/2cruX6nnqAJTGkRWbzdFtBHN4ag7PG
Il+xaQ0TSCXjurdEovheWbWZIJyqzQ2DwmaJGxV49One5pjH7xGEnnCsPwK3AS7ZalZH8toVJDY5
EAIKfEevndWIGOahez23xgcY+t0wjR7Q6dYDsfJSJquh8YQ+rku9rKubUAyRal7d4mA387oScvBe
CDGgtYSxFRaWRcGfo2KvMBjL3l4vaK7Qxom4rNu9OZWRZ9PwRsZLwFiGnD9rrT1q4nu+D30GaFCj
TeX28ptzZhmbnic3uTTl78Knvv3kMoSv4sMHHH4XIGCLZ452J92DsmzGOG4RUragfmbyGlnJQwTF
ss62lGEdzy0KMFLwEibQdlgT4ItOiMVnQ4AI5+NI29YqlfuZ49rCx7/zHs1F8ZssuykOCNV/yBG/
X8O0ngBuXQAG4bG6Jk4RT/Fye8h3wxZwtzL0Jb1Lu6mWxqQOxzjf2DzJ/vXR8f3MCECuOKFNPuMV
+Ibf83ZUFrQwgSmXU2eLSbwr5ygVc3RnJgiaJZFsk3CtZXAKRrJ6pKsozO6ld8g7BphGPsxFr8u1
FA0sDhMyzS/6q2Z0h2JP2HFn+FrN913fAv5KiWrOk52LQvDig/fF0kqE9C2/rig3yjoiSnn9jx5j
vTl0eB/hFv2f/U53jwbq0fl8AbqB3EZHlrRWk/2MxsUBFy0BaJkkqFEoSuxTZJujoXPyA8vo674U
j6v8X9nk7LC00BhgLBqiFgG2akHP4LqK/ykkI6sfJX6fQKbEnlsvL6Il05fS+7doPwONVSkfjIkw
X72Q+5Z01M2e/MEzYSY7poCSVmeJNzptLBnsqGp5P9b4GuLnRdOI3V/dV4VK+rkmB8K6YH7JoVqN
+HIdPS5VRRgVPOyE1dp8GL/gdBQPO5P/gZYSI6906kY50lnw61/4ehG/WtT5vX/dakIX4AOxjX/N
HF47P8YaLE6suaDfjHbmiKm1u77XeuPrO7AJtV/sQWoTU+wzsjh+wZCoy/lxDuLjr90W/pmdQmyT
RIxRrqVyBqiIw6OPRWnbQT6iglFP3hIKLY31EhSYpWcEjazG85nQvsVdovVPhbrs6GJn4VQIY2u6
3Kgxa91X2o1FHpdGrboCOwfejvrS1OhS++7giMS/lBCS/Pw5b4ZXnUwsl1yQ/j0DX0X9Be0Ad6Dm
ejKAxOIe68ABu6fe+VhnNSRytLqqbeQ+/YKzXndNG9MCLpNmjBcYxyP/tnqWmrV1HUcdyEaWXKGp
wqBUGxulXT/vdD9QhDUVx52JJv7ZYVnG6Z6jGLYdh4f6I2FR7jANSK3dAEuVw5eFQ1CRYqoqhaTq
4hgjezbY5NgRvqKndh75gIyOKXKeZT4UPQ3b+lb8tM1fhNAzosQ8QC+NDkNjkVsf6Pzz6mwWAipf
L3fKUaiqHbOMeovUP75j6wfTXfOVvIgBvBZdpc/B3PtvJadgKxLyDKhPaLtXi06lPLfv506UAobl
OS/gxVQVDcdZYp2SLA/Ne8sQ/5LuIfUCfjdE7SEfcul9CwCIZqtX+NNTfKPY5dOAkuAa1YA7kzox
CCwyS8EXX1GmAdI3MBTRNA3STs+IPl/eWG+Ms52G6YdAX3kPtWzn+L+Oy+KxYgsdPe699kbt1CkX
5sJaMMUcjTn4Iw3iMroh1gBx6a+Z5s9jRctC7WrT3saZTAo9HdFBCumrCyNpV8xvEqWaid73i5IL
8bKWR88j72/c6pYEIa6XXedTQlSxLiF8C2ohFVHrX1W6y3sC1ePhWGJ50r979sqxMUeh7fYlz7K8
jDacucRChtxCkA51Nh2XFL1Wp7E+39aJj+eEopbcb4t61PQrLlbFa036SHH4Fiasa4RJOrcpfGEu
HhYItrMPI5BWt5cCdPmex4OFzZUEoTjBeaHvajcoQSNWbMnjtXhwpmD5PRISJP/PbN6ztrj1Y8k8
msMHyD2MGJ4+B9g/v8WanXWiMyPf2mdIlcD1HaP1HGeg2xawZO7HUScPjoJVFdBBvh0Jy3Z/SH+7
LfIaWVKz3y1xbCtPc9Yjb9hhwb42mawhZZ+StpY+4Ahhn5gHiwk5FEqhOQlUwvewQrdDUwDfbQGH
CKlO/6t1idlexhvxPsMeCzTpGxvSt1tF8dm+Ie5rN6Pd2qvMFpNdSyNcu42VRS8U86FWQXAmxADs
AGsESw9T1l44m/WQngtVcgvPTdFYcbuyQTVJHjy6uPjqYxjABTop9rYW5fdcFKqqJP32FhQh5qq7
jrXP0ncC+YFKDTggffRoHHngeurG/nXcKsZlVbcWHysuSlI5IjCm2pcM0e7Ce4kphp/RfbqFRs6P
kSckkpuhzt2eCFGXSeU58wHHKg9eoifXfC6XMRc/qoNxKF+eru+gmEt8Xv2d5hNrl7rv+a+DdbJG
GBtfUFq5YQkFUu5lAuQYBmq2tuZhR3Cyq3lPNevlav2hE5SM9zPvpUHLlXyKwhnL0oYnZeWtf2at
TzUpAliIQEK1mofGEWe1trBPy8UqnShaIV9pRJ4OcyAZix8CRn2nO/jEqIMmI77sxjhy/qquQw7u
6D42OaKISY85haRcw5OL/QlBkWauD+mOPzITtnreM3iBd2EcUl53ChE0dzEEfFr/1tukv61wWh7m
wDXFXOYL0UqM5nw7v5zal4IYrGWu1aFd3/jLqvCEKe5GG80OrYpO91azzqxV4bTcOg7jpJOhnB+m
hzNlYxqJinYXId8XstS2IGv+VGyVgYfJBD2rGCH5JlIde8Bu43IYE/rGiEZ0KNQf1CFtXN1mFhh+
0a6eUm6OxR6aiyMN/fFk0ndLbDpYmmiE2AzLCg9yM6aMayka5DOz9BK6yvRtFP2UwXNICPmlOTZS
0U1jSCX5cufceS4kzSC6CeH/L5WIgw7XqhELWTesnIrPPB6E1IHVsfMt8xp8a4p10sRlCBeCb/q9
tO/5fviCnoSsY/4KJkVfVqh29D7+weUNJHndA2oKBLCmyQcI76zi5IZFKJlkRqP95AYH3D6me/nl
Ogjxallyxjcyb7uS/M753BqxPU7aACL+rHZ4+BtIYHjwTU2OSkzj+4rDci3j+fw0BV61q2vbC7Zc
IGbvj7E+Sbs5DRa2GcOm+FbFDcgvwmJti9l/S+vq9HYtKAJme7NyM/CIDT6FQpt9UBszjp8JnQLe
ZYo+1KE9/I99Uvtzj4HNQV73WJnueyek6+Zk9W9nTd6jgsnjRzPDibN0FLuLZt0DAGNci1xVCv4S
5vRWL8VFx9eUO1/wGTisJUeoWF7eA9lwl6IiyErb4BLuSxBg81O9IIOe6AeXgemJC/gL1TXJiA3X
nrXTP3bOKrpHtv+QRT6BBSyuZekdxu5+4I+HM7AMi1KhtU00Yk2GFj/HWvW+XYZrsboFql+F6pGQ
908ml5e0buUqIhgHcZc0g6jHb6/XeWz/FqNdTkXTW9Sf/knX2+FJsIjo2niSaIYr841kIHGDNxek
33Zs6mQ7zTNb+2XnZiQpQgi2jMUNpemm2X6RDFQNAXkWOUTdp4MoZXABc5ZocUxWGwc1dHbX90U1
0kfB7s4QUjNcXhtSa7zfZTat9mZeyGunr9/gL3WQTsXfWH41rVtZwVJRgOzSC/ReyAQe3Q1SBSzW
JbgkOBVBLMZpMihVfSwQCzEYu/qCo6hh7sG/791f73ZvH8Upsj+i0fiqaqWMLPGhY70weaH21yHD
b91nolpn20BXUKskJd5i1aB+347p2wH8dgesArzj5LvS5YcVhgn5KIteIeYbxS2th8myHqbw8+lX
jDibOyDU8cpspYsVaBAL4KhSy8TS1BBJB7X0md7TYNXNhd+Jk8T/y1DrV9k3NJJlX7JMarGkrNdm
7G87X2+wToMEJO6p0KjypsDoN+H4zVdXGGuUk4xbOKtVJkVXgKsRjvxoAbEVqbsAUYacY7WlRvFH
8xpda1DCJeAX8ChWTSVfbW7zxh339dFK+qYZvvb88RLFkExe7plo/K3yHRyeGpxPCUcEGJYW8ZRc
x6gO/s5wCQP9Pk0y2+PIFvH3JOa4weTkb1T3CGIg3yAmEokjBdSendnrtQfiuEWYJrzfZXhl3RDE
kNCxz0dmvmyToWuHVbdIrEPVqRynxZVhbVlATNobziy/Sw2r2z8Y9o3U8WKW3x66s6Dj2Aannsrx
4EOjwg5sob+FBLMZU8bdXhVHaKjTIgUtieBM0gF2X1Qzjz9GGa1WaPPdgP677bmvfYAUIUlpsoKK
Z0eeyfrE1nLMpJsh+YP2F9XWDazMwmD1biOFfKjZTCVwu1UET0vBuvCUu6U+JR+fFrlQC6wpmplt
iqt2baYMCkbxflSy7LrSdPEb+FqWrc8KT7F+qqpi49j1MS/G5J28h14DUYDzhPffkRFE2LSkhrAG
KOoiP9jEZsLLtI+32kvxyvXuN4BNtHcJyFViB/lBcteOmmGqF+QIjTilllbtt9mos1AecJQdOzgJ
trS7gMuJEcqPIx6uzyKm/Xbiym5nPO91yCdL2hTTwKqDmy2dcIiuAgPWmpp3djuEiHh9PJUmSQlS
TPNy7xpsAHYUMIw6lifZuzjMJ3/JqX+f5vg1l26ssVJF85A4AjUGxiGpu6Y9AiNeBVCAVx3WjpaA
RDzYjpvlC3Al1n6xAAtzQYQ4tbDdf6U72W4Z98ZT7IylrPKPOe+T/BUotbHnn06Z3P1lQwPyjAPn
zvbN/5ztgFaAsOE5mUZYVU9xJFvUnBwF5GcqjOCN+mA28mvBUxtCE81TJ1gNMf4NBpPCiZbk0E4F
FQarO9PVKEUaadcimpgOAqL9ORBrWtFkLFnxeEgPaP+a8QbezQFZ6klO3IXqOEbUsffrWSU4t5m6
IAwMDbt9H+dFW9xALZah7D8EMoEjT4g/rJ8HKeQ0VhItIYJdDHw/pBRTardIJ8dIvb37BW1ualNR
B4HEYUTNpbysSjybzPCoFDlL+mBCsepd2sL3EEcjgKFE5Kdu+RoSNl8TeI7BUzolXpM+1ZzRLnUK
vJ1dAbX/t0igMez+XJuk3bvPUqGvA5HSHJQoH3RcKwAjnqV1JfuG8BmbAHncnltovfdvEIJW7jek
5kPDm2eiKbUJZzw33zK539yjq1nl3NjEnPOpFrhoaKjFjSupr2zKiy/7CtEBWH4ywRkMB9u2+Mfk
Mv6eFVkQLd2nFL66K9RrYhta1p69RwM0x1MOe9w1Meo7hqYdC8ZVpjYxXMzekTC18/dP1hxO2Q7Q
ig6XMxkVCOPtvY5EQ2yXvbjyi/r6hpoGe7XF3f6l8dfbBjui+t1eko+SPkiz8C5ZpI1E2VoZZWvh
4CnyAr7evJRbn8wHxDoW+Zlt7UFNA53RSwR1aMGCkfiKMTip9rTuGzkdORoNbdwzMffqCZmvXAbz
plFLCA3hTVuZGVjBvxmzskbQDD8GYJMXEqPSbVOvWEAa6m//rXNWXOP++2sI85e3C/7yOGQIVp8x
p0iWP4KKEOvLCbICpoo5rmZxQuFUEYL6cL832Gp506MoEOQxyKAOy2K5tTrCGrTWe50XPZORRtM3
xRajJ2C3TSYjx2j3rLCeI2xlGyGf+h46HhlBXK4IsLz2MmhN/2gR8hpMrmWtCPp1NLeh3U/mzERB
2uQfoQDI8EvfPf258w68i9O65Hud1QOERjVE7EPxgBCWkEso8d2RfVu+aEw45beFahbGkuBkfDYw
1WE2KbQYkZGLam9uMxnwoMH/niRTn/hfse+tfAVgX9Bs4Hxf1jKbQTuK51RZ0sTpn2A0Ae4hYg6x
uxZk5H/ruN6eLj+dpWJb7oAwEynl8+L01+89v9uQ7YneeV8AJNxpREgf7X/E54oclZt+TqTvGwtO
vuG5clYJxumrgF0kmLr+AC7Xe7qj4+pJ27ByCmPp7ryW2PvCYGM3TZFCwTGDmVCv35YZSs0Ru20H
6+0mveQ64tMrvC6YcAc5tHkoBHi35KQnvU4cD7+Ah75Sa8Pebj1X2L1DhM50CsClEHkSDzL1fGu8
8bZXrQM36dd88LLDs6kgdd5AgrrfNsFWTwK0v2pJ1FSieZ7zUnUSiTpTrA+GjBuGmlCsGdtQvu/F
ppPpYzJmhTEi+GoT+ODgv9YESkZqh3Da8dWoRs+8Fkea/OpRkwE/MDb35U91EjEv3y7VsEHliitD
8EVHsekwXZNTvuq46MpT/FxX3Dazzh6HLYCmkTa75rHDZivB2KpUfaXli2+cUBcOzcUNgdE78lCj
nOWY5s1TXiy07y7cShguJbGoTMqDGiq0rMf6IJryueN2OHAzs6ddY+TlCODM/92TZr6fFcgraAEQ
sA78nc1R1n2T9+WzOn0rqdOG87yfIBrJWy8XoZlae4nEM2P7d0rpANe5Dp/dw/Yq4HXmgHacqCZP
ZI0fV6/jPGrS9ti+/cAEyAKHeDavrBhNSVp5zgU/w1ouWXbUoPRqkyYd3Wky3BvIstVPsEXlBcWm
DYsa5ir0F5CL8+M+GOilCUm4/PKRXy2wE5TSjUrJlM6/xWa8yMsg4CJMipOjUaszv9H7yOF97Iu7
lH1fhCgZ9rrjyFWEKNG70z98XMXqIMD+nAIVowg4MBDbtyZg+sMLbS/Jk7fn4JMiVjbDXJVDxofL
oHamcTLk/Z8NQXjs/vAQIdPNqxonzF7fiz7teOs8pnceVyKeFQvbON6PKfoWKD6lP6fDqPklYPHg
mtNtyR7oOaH2b5qxviOZs1ISbKmwJq+dBUQ21GQuJI/o+HfcJMysKiqOcNS3RjItk0YovrQ0NAn+
sS/fLZ8c88qpmRwfmFhJkTK799pYgaKHkgsWqy2PBSN82GvkABjZbV6NHZLRUw5wOCwHz3fURzks
3TwD2R45e3hCP1fEmLlH0DODp2quwUz7CKOz2aIhh/20AFIz0jvbB0ASCtig+6VfwRQbLzkLbOom
5hnJNmhkDmDzMJX3ZG0VFINME/Lem0l62fdHBCCJ6oXyt78SHhOwMCyEKwVf6evBsetiyIO5Uwlw
fdochYSDDkSTsfbXmobYD9fa+ibjV7f/oaNn/wukmxdn78v7hkEqxF1I0jmwSdnf38yzpPEaeVV8
6nDKp9EtQHN4Z2ZZGtVs+g4WHpma8Lw+wsqXY11Z8lhxUPSXBAeuj3h59U2zTuZyvOEBecW0PZGK
+Db/K92Afq/0pEhkOHJAWJffhFKLf9C1lglg6b6cd2u64DbJQUSP6ifwmeL0fyu2Pk7HuIS2Insd
UuvxS6r45n8cXx1+YLjWQKiK4j9sOsSdgegToDQj8YTb7dXlxj0ZjUkhbnv52w26HTHd4Pu1Q6eI
NPZyE6Gmi1t+Z83BUtbZgqn2CzkCJ54ErDVNk+uD2LARFdFYS5AnI5x4a6J1gNmx1xyJWZMwr/bW
3mjrJLIQ6JhIVGnjabFcJagP+XM8kWrWqluEQmWmeUe5hX/+7nsj95HBrR4LF0f33rD+n5IbnIn4
rf48DfIlr7+YTLxzFEzHQql4zdqIZCih0SiqvBFwVPruqU8sM4Yo+DwB6N/ytf34xjeY+8cs7nAS
IZLGY2WB/ao+S7sul5sE+70C777NXGstaV4sQwId9IvCGjrUlNv+YWHhY7nqjusH4iKDMd3n1XmQ
qMztuSlEKd7Cvz145/WDUjw2wteTasY2sfM+5G58QqhNLjuxGQyOmQVS1AiUdT1ZIgexu4JfQrMz
woyT+9qYKyjRVM8JYFcKNq6vpBkHOg3w+QSEPCtF/D73U0O7SvDPhbEd5FfUCJc7Jri0BC8K0+N7
zAZ4Y4/VNjq2hhWN9iGraE+tR7P28CFLo+suxbZanijOT3NmmwyFlSVRnLL4Mvm19Pk0XQpAiB0C
A0VNG1LTQ6esFnMtnUzrUHSHsC1OLaY4e3ghv+ekl3rAXUNu+UB/fWnIxDu7jyVmkvwjL41UBD/D
R3wnROEG8Yu+DDony3YJ3gUwW5NTwqqWEbuDlFj709+xNrX04ktE1r3MjQfLhD5LamRRTqeuVZlg
wKvnkJjvURTomUhqvd/ZIK8gJz0OVjmS3JZFPtXdWomSZj4FkzyMN42nnrAi9pj456D3I2Bhsvv6
g0KuP8X+/hghWSg7xf+efjWhLYpn9jnmvVEgB5vR2/d/OLaf65DpmDZDFEr3DJ0Yk2nYb8vbPBUW
kX4NCyXYXxn5jw1LkAs1s1ZGXyuqXxmLlcOZD+oufVGyk5g5DgF/eyK3ZIm1TsooUE5vz5h7lgTw
yyw8CFwloWnzgs4FrjdWFOgX4QMURggFz2YdqyB99noc/FBC6uzqD+dHDN7Z2DdosPlst7XCHQ8C
Q4xH6yu7R0dncaXPpxzWj2CIdlL0Ctr0idsMcVrE0Su9aa9w2XkBC/yJEkNXhDcSoILou+/R/JOS
UKocYax2iFCD98/gQHnAipoNXqzUybzgYzw51gRhhBjcIog3DSZ/aRNuAHF+qwSoQhsyrxhBjF7V
dpt6gF2xzM1WmJBdWzG8WBuHws9q99ZJIytiySX5pzyEv2MCSaenaiMFyDcvBjbw2+y7DXuRQFhf
ZSn7FonP+KZTwSyyFoZs7XaaFsrtfbRkiplJxBzG6CtHcD5R8j99CyfSs/4bgdphPUbyY6tpXh6w
LP0MnQrYOeIGnIvgmUT9g+9WiegaAsW2NAKUJmYsCOuz2UlOMRQiV0a30qbzzHph8SWTILC2UZ6X
yRGbjHtDH3KqTXsqY+Yf/KFlw1NFXJQmCxpNhhZCE5nYa8i3yEEtd0faRGdmFBn/BrxOdv+eJkD1
y5kTwMF+BTdCYhoAHPtQMG5vK6IrVc2cideTXBuLPaLQgtdxXhvk245uECY4I8nmuRJo7gLylFyX
5NcqSc97Qh+jwcN7NfqpVbuD4lWfFiN37z/+f4KDL6b3kbxNYHtV223vBPQbqRcpbNDU5NY5ahBz
tGEPnBlh9oG7TXjxO4LGCljwUd76GOh2HbE1d45c8sLBp1KKGg/9/pFbwpd9jXUlo1Q6TFtU1Q/n
g/a5sbO0ODfRFRlGBIfdRItUfu0xgmWfTbQMjB74L2LYUemF9CTnxpLv9+nwgkC8EiFK/K5u+Oe7
Gca/xzZB35Ixf8IoRREWCAgU9AbSiYQY2f+jzG8Ox1itNotZ6a7cqQEd6dC6H3fOeN1Ijzb7hJTp
ObL26lbQ8Vfhv+mkuBMtF2Os2wjdrnHqeZ/mZRBXf2dGNCYCKGyQWC1LYbEOaz99EI7ULaWIELuT
QaliUFBk0rsfS1nh1UEdCC0Nhlb6bHe5i8Hm4UPItzro+x/jssAR/P0NCea3Z57i41vqNzsgYCpO
UoUI8ANyagChaccCQDLTDO4PAEPImBfAnAjCrWrxkaQpl4/OcWxWCYOdFV3NJVY7ELvAvjD1QHFF
jsch2d3PDa+YzdbZ6Kid4D77LlnSZ3pdSBeD/rLh920Ca2he+tAzZhdgKW7eL4ht3QT2doaZ/qmB
Nxl4YfipqsJoKg+e1P+cFfvNAndsEw746A5YH95OtnwrfhNwR3SK30kWdsySksa1yZCJ80g4qU8L
Z2rsmhXMo3/Bf7EXhJmOxGBs/GqN9wtKLylGEONB3iPhiL2lkZMXo5WeKIGyUjs5HIRMqzL9oEL3
1C+ZtKIMgisGUWQ6DmoxBRyVvdJrpmVDiPBrDeoEuMyWIIQ2c+d3ecKHW1QQtnytgSYMUmgc9aMW
WPtEt/qf3Z1pEnLk6kLthsO6gh5Y/soLbgd1nKw0p+QVM/Ql8YOlD5NV5zqRIZh8UiIrTqmoHSg+
g+vItc6dDIMK3UzlWDMhhwZBvmti3H7NlIb0u0cVR/VwYoOPRC/CRNNDz4Ix243aXieVXQUPl9kO
lKLkOwhGN62iNaXxREQHklHxw5zwP60A6xl6g7Q52wfqk/j1Vz7DdfYkW3jxt2Jl+sVCpbw0mpU6
GMgBas95olMXyXS2Zh1ciu0vdgNY/iniAhgcARRirYdCJh9nVA2iYoiojFxl/ljawJfMGMFNj8IP
WNIP+peAlDuNf4oWyafL/n/CERFvVcjVeKHSdHWgRkKOQREH/Hvg22RgmgC8mqRg4fhIyBRcbL9x
XKIyGfqmzeQQLPEqt8j3KOQDGcUlb5NGQLC07Wsv8IXu36M1bm1tMXxHoZBewazyaeMAkJpZ8nFy
meoN3EWVUyEk3y9HIYJVqp11o4Oh9vKXdeKcyj1/ATHg+IHC6TwrE7VlYzzU6c5wVFj7MopeBBRL
gegNjMPpxMGsZgkz+nmNFCN4vytr+HU0zNRRP/D3Gg5FqLd2HHgtakuRtcHXwricUHjYZqIpleg7
CZTcboibV1DpkNd0Uei7lb1fvf5kbd1cqwYPJ7fOKliyWtxfREdjK3I+S0ESkgNYI8aF0Ybw44ra
kpydx8LOTT11fLEZzbQuqCBjtgLcJwa3Wu+tNvXZfUKTluXEBBZNX5HRZDug/0PFhxv+rMYvTG/C
5kRlBoTTSOfDLV78Z/vwXi1+KfnM8X/2biDqAascr51GRKnI748qr1Tvi/H+1t20gw47ioBGaxpk
BGH10Q9I2AwuCADyXDNK512zJ1h7CxGkjWHsLT7AMREyEBXIhUfg1qAaS8arfFyqrLvRVWJjRUgt
yoNOy6vzutV4n9BM9mhyzqrR0h72ubycuoazX8y5BTbJQXNcI0Cl8HAWbqU2fiUoCsuyvboqJpzA
IHCbq2QVcz5zwJ9oYeHviWddNkFdaDZbDHva42BYXh4PRwaDQAcMBzNaq/Q/iIVL7YT246oxKj6Q
gOrZKIr26ISLbXEty4omE9gVPXfCt7yRBteqJiK3uVma3X+ClLhZ9RkAXFG0qRNqmTmWIuuB7lN7
39p+BMEQTnBo7WH7VRk6jhXge1fhm1NxO73QCOjbhccq7yAogoBpd7Szr61jT0WD4QF4vHkjXxJY
+2ph0voSQZNW7lM36g8tTvOo/X/L3OQuxEwSip+fADdheQ1j7fjdIonSzacg1UM+dKjaDsICAEL7
sxn4PcFQYw7Lqeh0suxjWFGEstyoOO3oqCQLeMEmo5uupoLNVOKsaoSvUSFQDfYyLLgk6fH2yJ65
UrFggoV0UbWa9Eak6T2TArBk91soIolbqbCDFUFeYSOtrNtiutUss1cL5j2vRwF7Ip6u2bZ54MpS
LjdhLO8835qBRpHsuzzZaLeszKoZxr9epAkuzsxYo3LDqdJMdL2tgi4pA3zS/9HrF3wwxsK4sQ7m
LS9wPD0LrTVKdZowqh9mZKla1HuDWxoC/qXD8iyCPWUNsIfY2CLWR6jbntbzFg3P3iSkLJ1vksOr
ZgoqIo5Q+t9pnP2jfx24M+jUmRVMNWj1yjSG3fqK85CXrbX0q5UMfwZni0/OaSkvpBJKhrTMP3Pe
4YlnamWRdchocmefl2eBA7EqdEPTx852jFekLzAewZP9oRQtWi4RDI1BnJfnf3G6jOPOdnoFmhDW
avx9GZuEcjSySVKxTPQSnoE/8DHAbNt2UPh24Ovw7TrqqIIzzcbCN/7qUHfSVPkSwlBnBpyQdPY7
BmJMGkAZf4rqOJD/JGlAimwea8fpkvyiVcGYqn8QE+zRW4BMuPTLMAFnnBXR6avD+SUps+mxCBvg
PGkGTSr+gIaiZsq1a27saOD+eMnWDhHn/7GVMiHJWV2ctsJgvazamPv6G7VczMqAxwRWDdPMxJxD
401AvMW9mf6pNWK58YHVLiW/GngjErQ53qMg0J7Dq7VF/3HyuEHhclrvjkIpSOJ0D7FmOCz49frt
Q+/iEE1W/14luhLCCZ8EatXNF7VvG3Bt9/6b/l8iwe65tVx2rylxcwRQSLBE7vcpZNHBFLOnKywu
npVyCZ2LkgVCgIIVoGNSAaC8UJrDWKRyUgi0olbGGUiKkxLazxuoHQQ7QSj8lcaJBPdjs/WY6fYt
cPJWVOBO/wS1/WCmantuzxmp00Zgel7vBFh6sfImHIy0ZkD1+4Ih3W8gCzTn+19HXw65yawfMvhR
uOUvg0T0KrhuFRvOI9oV3+60yl8fQyae/RRsTnhhJtktoknQBniySwG2XKlS5IazIKZ0ftfgrnfC
avKYwL3IvkTjifwJmvTiYGEZbENyWeDIAeb09I6RCD+WKSCJM8MGlf/cdjQs1BYN/HmX884FyWJd
kP17fs6U2yMuFj8o6RvCMoVeOyAWcnkJyRIGOr+/3q+oHrGmxo+A1rDvnl7+8jbeC5AbFL82XQfe
fwI+wv/ON3JaqCfZ97jC6DWHsFS4Yg9kBnS7cOf4Ium4H2ydwIa8MgpsARf0aLHQ9mm4REcZHrLF
Ifip6kwAGyIzQAsjCgJ0h65O9aWapjwyrcQjilZn4fAHA5tmbL0U8fCugBcVFuNUw6v2Nq1HzGDw
66vGfctYHhA5GGkEOnEYHRLXUu2prJKSXYCbkvdlufLJ7+E2BmeTI1hXgu49OkgkiEMb6MbQZIIf
0O0Db23mnmlatB16IJM/WBHF3YaOAh4/RZ+GbDkC+xEuxCbxYyCrLD/9nZaB8lyh1FwM0/YR6SGW
wJmaTzq4VyZ1oWdp6IP8hMBXZqTPDimwBqTUZWO6vVjp6s5zJ4sRUBlglRBD6ms3UVybUdCWEWwW
pNkpOuJeIgHqP/3ALtP5qs613KnPn7cSCVl2uB6r7ory0XTnvpfdd7Muw6gNso6ze3y9yBGhRYjg
dhth2tx/z2+5ilfEvcY4c5XzqUPNmarZ6jiLu1+OhK6rKihdVVcvBIbHkwJJdFzuj7ePjcYNEVOu
n65BzMxPiyz4ijO0NpQgsnzWhwVLUfLXmRxKmw2Lq+uLXalgijswZU/aDqDhK9FZMif7PNNj3Ol+
8lCemG/oBvG5FCgT/WuhRMTRFxECCPRVqL8O1gS8bnyiyqCl44yeEtQb3DheObW4GRwrXtK7ImWX
M0QpxRcO45vPRxsvEBJaVgZJmmbQygq9he9ldF+tNYQRXDZw5PxYhSMy9KnzLREZzapWFqqN4Jgx
nudiRP4Ahl62O7rcO4aqArWZLivj3RRvah1AAWgXpq0riErxYiPkfN7XeF9hsGkXtOfN5CygsQ9N
MhDFVcsP8Ovhkt6eqnPJO2kE+flp5HUM4c+eWL+lDo5WLT/sH+NyeRlDXTwGSomLyK0m9IX+P7r3
/SeEWIEcLWlNvWaQQvHNqE5Bz5gzEjiG858bB+gLacifrgDpipo1gFCrSJRRH9W7jnOCQHOJnvPZ
DMcEosqqNBD8T8IgXES2MFCfTl4TJ2CccVL/budKTe2MlVwcPynmuINdDQhS39tt4ZGH7g7a7BVE
tUv+BtKhOxyzGzcHwC/ynZDP8Nk+vEg4cKesZ11CBkAo1pzGEhqrSZhMi9PMz03Vg0uf9pzQOdDb
RZ87jeqDE/akqZ6INqdz7vv6Xxod0hEnzOCCohmMO7flUtsvmiiFweiVQykmlTELAdZCRlfltMRE
Nd8Y9DBZOeo5HJxYjWcdgwpq2WmIVsOtR6blGZ4v0jRK+LahZe+LcSnePzo7r42S6HMoaSdfA5dV
UckfKjH+WjwxTtRrgrJ4RKPKlBJ2bSU2jqyfGe0YBDRDC3T4tVLh0aIkaFlc427Yd1sOr6+FNyDd
Te0kuw40c6D2tPfTRIkso2QEXtI5/68QO9q3AZYUVg5dhhTGu+jJp9f5z3gyXlE9fn0eR+flqYm3
DxteeW6aeLBB3GXSmbS2Jq0FHzLB23SPkxqrs3Q4Y8UPF9/z8AZVUxegTpBYBEmu7/fEv0J8XgGR
0z3QR+NhFt9aIbmP06uA+Vvz7+fqKqDd4XsXasnJoyQfv0mWKvq+vd9oD8pgaTsFdexIEZBtlL/r
Ga26ihL6UACMgx7jlXlJWpq4fZJ24nLEM051YgCUA+I0Gu+8gvZUtu6bso3vkIUEGj7aYe5sjgkX
KQ6WrlfFRbBqP0lVZ4Eby2ixhmypP6J4ZuAsgnS2GWSqWCFpJhS3A2WN1ilP7/R9iBFiDBwXNuQe
xMQfJQMmwxRQLHFTjC+G9avlb8Bdc/yN1lD/H68Jjpj1zqOlCvDEkA1sW79ezsCTb/QuhMIXD+U7
woIQ+qWRNJHGIGCKmG7BwRnd7B6cujThlR80cT+Fr6Vr758XEvCPh+RzGrqWVuoq3DxqYkaMEBQx
Rh+4iuHajxIY76cSgRVKXUydkZHLMnYYw6Y6zV4Md5mdLZZG5NSpwUd2WbV8qCnkZ0TcQOysg3V9
JwZFd8Mj3xHqxv+mxywhdbZGRp40oD3zzYfLUZqqiChEpR+c75WS/gV3jexqId5etJLXfw5EfkvP
2szyL9/2Jh3V4u0z3vDPlyUpDlUPVGqkypVWPSqaZLe8w0bhSqHPbPGtuFE+Yld8tsrmCzKJiGBJ
a2fe2sc2XH0RZ0Uj9r1NRa8G6cOawEKQDch81VjiMSAna6xU7rxacvdxoxsUmllsmbeyuwuEhXdE
SmD8IGqyEJ+DhcBURrnrIB5YspPy2202kKxvy11feEqM2PvQRmwp1Cf0uDzfTfbOphXE4XksBfKV
KWLMqAzQ2GhSLfs51rmxNeGPOBKb21j8oEU7eBvzfpNKhKJHi7Y915Fvg+0NnYZDlqpHVh/Yv3/l
bbTWxXDZYzRQI/Y9PF7OvKpot9FGszjpjC+Z5GPPzc4lu94b7SIB29VOQHLPipwJ+GgG5wg8sBgM
bQzrsGTpiHn1qmVktngmVFjBNeUPKKwp0xFLg9Zym5SDD7k2zwovHj9OfMpalSvwQDm0bXBOMg5P
WS+TwPyhZD8xPVA86aJxF7WYkOUJaCgcyIoJCXVsGd+yQsgoNMvLbCWqBicF9PlwZ7Mw1YvFYe7t
wEJGw2n50RkP+meQbrZ58D8ZURXyJehKFZdJWyomlvd8E7sPs0yeF98Cg8w5xAfRhSOq2W6lOhQk
eO1AC3t3h11AYlkJvPR/hgR69DF2YFYj/QrEeGox8LjXJBHySFI11jOfR7hUwspTloP/1G3FF9fd
jFQkUHpDofEaGUYzaDJPKTjTvBVNms4CFVkZWLDyCXguLA1EzV9cb2rXOulUA7x/IzRBXgJlJug1
c9tYXsrf7N89r/alghL8IzzWwJhgMoSaI0hgzuIKzMw6urAIFrMv7gheh+AruZRfarCDNgtrcJ6T
UGeoS6Bi2Hq6loeS65Ywy7B6TBrNvNt4TiCsDaTb8r0pKoUBt6RRob7t9Ej5rFVWYkOxeVvjSx0y
m2SzJSgctocp1K/cqPU3sTjaSFGYLlCEFmuOnTICI6x/bFoaLZwsih08T6YbehRxdIRVOKevKw6z
NEmar7Tp0TaEmIZTH0Tj1z5ApoAoQL5OpJAGnCnfRmugmRxw4GRmIq/lGHT0lDyzHyqkObikMnUd
bIh9awWiVjnPY7HIZJ8iYMCFi5ErbhePVzUCpVxyYp0G125wVu6bhd7VVOzOYvKAdiSad360cgmC
Scgw31sRKjYSzLl6dUidVIQOzKo0PvVrKECZATixA+VSm/dLlJH7W0WU8UU9x58XnrN6lDeKedP3
GtPZB8MvqLJ+6FkH55IlqrPXj/cGQ8hq1TVuUBDZtg7UBP+tqa8S0lxVyiQZLxzAYscxII6efDs6
8J+suIDG4iSzjI3eq+uskzOT2ESVH7G6F7eO2apz9XwjjihyHXDsEziMB8pEZF6Y+h+A1okr9BDL
CnNbNyxQodAui0suoYLr02PNSvyORvq/oUrtG9dFedZiaocfPr4PW84tppdqTDl6gn0lZnGSlE3S
1OoJAFZY07djUKZgY/jXQReXgcp2z1Cj0tCHiX459qXvsPxCCqyieblJdnMwPP/8cukhEJb88L2/
dlZ4JJH6WzgGKbF6eH3QfBv5j1rrkUCoh27CduPysOHrpYQ30jXBjjuYS317MrGlmFTWwrxdQZ1G
62XpWSUE+5Apd57NBS0c8N9rtRbkbwuB4jbAXNxMZQO6WMoeHFvHyuCecoIhzI/2+6TuEL0Hcezs
/wUavmSZ/RncbkmpoYYDw7nojKswQ3D1f81PC5ik+LfdRYhp+xYaw8056+mftVdlwjv78AmEfyvV
AiNJWhRq5jYpvEBTYUfpL6CHqE2sZJb4ALQfulaKu10Ld9lJ0cpH7Xo2AFiQZ43hTQX+S+prb4t6
ZhQH4PF9QpJFwq2GahCISWmqSftV1BEyhJf18NS1FvUPM634jl9Zp5vGIC/04Ah4w5M8Z+Tm+QXC
59PPASJAtw5ifzvFKBrzkaemrKwm6RCdSRKFugNd5206dEeh6lzuXQSUXmYBd0w3OGecYisL4dWO
5Vmuutvh52AArmMQfQbWG5y80CBJIBRf9JKtGsbl4wwEtOFuB1leULrO2Q/6F+HFdgk2/YzJ5wP+
VkaRSzMuZf8yCpFwDFje68vxhhzu1ca8qtcnWlJQ/agIS4styOoTsfhJBv9ufGSIZiUuz0T8Dk+V
Rm718Gwjvm1GznVC6Qt4ipUs9kqn5p4J/EDOag5fA8ak5lBct9w5e4xapKLuiCKjH6roVnCUUbes
Dx2ufLPCQ6YeS3txCyd4V0k8eZA3+k6QODDjkkE+hYNCTiO7R9Wy4ZjNZ0SE5IWzeA3bhsZOxN0x
+I0Jenif6EHPwrL6GfhK54gaMAZrqX/0I0MiR/Np5hYYSVc6kBg2ed4W/YnCjXO+zyOrkH0JhHfh
mLQfCtYQFl/Hb+EaQi1zQ/SvZC0zr2QY1wwLzLhcz42T3yCZ2gk+jYu3jKAvruIKAEZkIV0IEc92
869Lhs2aX8SA32/flB9EP1JNM7mYAzKjpBVBc8JnYnaSnc62882ygr5/1lwXhQTtEeaU2svp9MAA
HiVziLs2ER+CprVs1hQ35VNiOyjEY83i0oKPU2JR9n5vV5FQ/k/SgLysT4BQ4JPB5qmxI5cIxa6X
7629fSnxxTXwm8Zo6Qi7Cr95I6+xX+TOSC2ry5PNNdT1dHpjyBmS4AKTQ3ivTe8uJPojA+AMI9ko
PSyHxzyIFmH+8GFllINjKJpqAgHrWEfV/AGyIN8aunbxlL9D6BZI7ngA266w4guuFPXbLjhx65uM
DroVRVdkTKCvhBTRriNc4Tg3l9KWtCizs4qmio9OKevSQWV50hST/BXZ/2UrIayeKPayA1bYa8rG
xT4ZtTHSQWBQqO8yGKMZAZwzqb16+wkESstbVBeBOd14w2byV8a4Xq6l8o9TeB70Yi8a35y0PXON
csnAa28NTDa/JZ5fnuPSUxAI6c9E6HmmHDrrQVSRtxctIJxq2nBhGLkpAQFn+pEhWrzHZ0yqFhyE
elcdT1RsRHqb5f04ELKYYfWxWF+/fvYeAVAuog7zHnSZ6YiPQCE3lbsHDbyXmD/xAy/shfkF4MSd
2pVrKCnbAMZXxBR2TdzOsG666JfiG4rdyJn0UgAYID+5NwiWKtqTFWQ4DNLOpnMlV3UJMpsAybis
rqQeOMrubhpfj77ClVTV3YDmVWhQJDjCwwk4PdAZe9kSjBwBiCpt5wKo9aJrfs9JQ3eimNWRQP02
HQLIkiHV+OrXlqltr/sdIX/O8iJ6vjURPLNHakVeUjzz6yz8MxvglRPKBQeQyHqIeGNtYYaCFFzt
MrKCWy8Jo+CJb7WUsHAnr9kF52ddlOXCCZYRW2XpnRjy6xeaKtWY8OKgNyVZ3bt0em/06CMQflTO
0p+VZAIDeFfBXQkwYozIkHE2oOzTB00ynFjTG2Izz9TNer6if9l7Tqfr8d2K2gn66S8VLlDSEwKg
e105dXrqbezEbrXjgVj5IFP9nm9/gALJ9UufswVvHw09mTazXaOekJVyy3w1vxx6Lii2b7rL88LF
n8wjxx3OzRWa7LUUxjhXcMm26XiFLyiGIRYdCv59LZWrVUwLpbLQv8KPh0c7bzc/pdnSriH8XtQP
oPTbWASSFcaPKHFaTdLdTEv0eqToTO1MhA1o8e+GPxt2wjjQrmnB03HlawRd1u6HaCJ29MOYQkwH
YYe0A/JKCGSruRpREnZF895uq9ZLcmhcrlFPBWCKTiuqh1lJhC1Cg67JUYxjl8VBLpFNV1gFP7F5
dc9AnwdKTY9uR284Oqafa3gLjfBsyC0051c1Lty83EkyGXDjf/9twIT5OQRzp2ZtayKHqRv9kD+m
TXYHb75c/1NuppU5ECYUhIm/gKhbkc9OcqvhdE7pLLRiiJR+sj9HhgLyGYeHpi+VS200nWPFwOI+
Ue74KGOHfT7rh+vXafD5VkSsRi5wlEaJyt/oT/Sav6gF7epW+9YRxee8aj0X4wK2O9Yf5AXJBxgt
deviezLmzPxejxngxTgWXlDs7KuRF8OD9YgA+5EOqeuGx051GjE0D29+jUFTewaZaCPj6dLxAOHr
Mx976tQQWk4jXrHCEqKf9jVHAN36jxoPKpgdAm4FfwVg/0b5UYlaA+aoyyIa4G/A/nRjyC2+GawO
ab4/BzvMvQsLKrrXvTiYAICfAU+bHX02V7JuItpW/bqlBxs+kyDA8LYfLZizksZrxvxX21NzU75r
q0PrHoj4YIj4BsmY1yxjtY5ZIfVXsqRbj8HB1gFcbuMLJ4Q5kd6Qwp5H/imcRaXWHprLPBkICCgp
ril+t6RfYEvyTMemFzpDnlnGOoDWJahtVy7SW0kpskF0qsyW6qnEcq/4VmwRUPGh1tL53qBKirh2
/Nv8edBnxvfYu1Bji/pv2i0VuPtwz2btkyPR8OcrFzXa3OFwcjoaIwDdAhpHStZ9YHCwFfs5cvbL
k6rnygKBdA95HrKSdxqtv8IqcCo3SzSlqi7caOqWRmyQVpvoebmB2jorrwoTmu9CNmnavuji0Xo8
4xLPyJANw13Hy43D2bJgxpvlLfHP6xIBHSTLqTCAom20YxLmzCjnIYHbBKm107qai44iidy9j1ZP
ndp5wfj7TqFTy9q/MhWjaHCl8VdqXLguJnqerCe6hj1WUj3AdtbuWzlOWMFER6oYErkAOYsbUOWd
oypdouOsw4pfXt0RtTmfKX6UJ9Lw4hMWwC2EmJ2wVM2a2I+loo9Hi2UtinOA0mQcYA0ZIi65v7N1
j4kIeRQdgrmkFBTW791i2KCxqjJ5sdEWwQG7K3nbnajPJSZWAtDT7oZ7/e2mgRC6L0Fmss8ECKAW
WnqrpxU9/A8C7y18s/z/BoamYDO+6n93lq3OAKVRkASTUFD7N/3zPeKLtm/IVIMXHSWd5VhbS382
HdZztoQ10mufbY+8ebLIiHXM+eR0Fl9968Rw081AaDaXqhAw5vP+XyrwYHXzRyro+svc1VjSHB82
LM9ufOVBYuFQprsqVn8uFVd6i10qcPwVIZDpCBEpcnJGmCzQg2Kolk0B3o5go7pTdAcoNbC0lZNS
M6e9Z5+5RH+MUgRkhmPVXdy2GA1+ZupQVrMWvKXYzrTl7QImavyCY2o8p60Pf3k+2+oSo1OJcMfO
GFALMDzM3E6Mv7soJmn9yHhsA+klJ28eL9kOchgrKg6GbaQL78vuKdZwSepwt8+6K8wJka9+R5sj
Xc4QYOmJfjS1Ekp2ZJQ3ohPfOaN8BETHCZNvKKTzik5Q/+G0UMYWxK2Fquzi4cEWwYBh7mDUDu/O
x/65Sne7H7u/e9jZmTHPs09+Bwev3nH0cyD+1kjrj2IQ+abyf25KyZqh8t7Yk/44sp1/LLRhr2hw
M9eMqV5AvcNB7bybwIw42xdpN4XbppGzGkkDtj7ib04mN1gWGIOdJUg7o7lcZzxFDTB/m74SKNmS
2DatQIp4j8HfH5SsdDtqIHWQiKK2CgBSk32qEH1y2NvXfE3zRZ3MZyW8MwScSoX5VG2yKG4N9Qtq
C9OowKNdNN7ezk48T5ZuzHNzvR5bzuN/DV30krHD102C9JI8RgVxOTkE7PX7RdBPnK6sZOiHJzu3
3yfUzdQzDFHhKrwv6XAriHpfY5s3sL0l72m/CS3n98x+8EEDWPfH5NfQceHJxbysOpW5hz9eHktg
L35E8N+40WxtUCVOVAyO1954z4d/dhSfh2PlLIJkOjrLuyQ6i4KJWB4lD8bD6FJzDjPbAESpJyZl
cdhuReYqaO2g6pHcD951ZydF8A6dlwtQtEXmGhUk4/gNPatZKHN6llQzhfm36uosntIR/MoKsy50
tUlBjiZAwLxm0vxFj5BlgVolTxDzh4Jy2I7B0pAPhNAG2HRHdzy9RINV1iq4kdShEIj6hyfJWKDH
0TGVuZHfI9Fc0IuJnezbrfOKkzOEahggGXkjCHXmvUV56JmsvzypYSSJXhaOjT0ugRcHnNV4NO2C
agQMEQizlqh9/MQoU7bfxosOJNPqZMkHWm+De7UfEHMNBA8JNYEB3Ohvwipdrgm+jV9vqEsy34SK
FMLzQAEWRxB4xOBaLjwNQe3cM82VKzY6CsCiO2yMW4B+dJYcXhAGqhEn1vltiZYRKUfglzwKA2MP
EZHarJPKinOq3UZw+3l9vQAgQKaSi412Gs2e9S/htL6/TpCBdVThTBREex49DJqEZtcyIhGKVVxJ
fdJv4ONeJpgcuFFlrnyL3SrmP1YADcR0uCilul4MH+bCO16bzzYmBSqqnflH2bsEsNiQs1LL2HdH
9vgsBIcwVsoE87WwI+BC4wU5cB1WVD7IeDJ77671VJgzxLzmJXjWSU6afE8mgTbSUBvzspgZ3wkh
wVDxoe5yUnxJdXdJqd4Tjrw83L9Sh9ZFfFDzToSq1S7pcBUQAqouJhqFSPJEOZ5AEtsBNIPC2T+4
Ga0Mh4TpbtOopfOQqGw5+iGw0QQkdo6E3tdAz6oA1Kf0yYVZq6vYrJZCi3/NHU+oGJu5FMZdttXq
2/RyWh2+WmL+EjY3iEk2KIZUgaZsxQg/Y2bjq+/Ul4muwOOgNb34/W51z8L7gFSGmBpc3S64Gdpv
qQHmKA+SdCI+nhu3E4whXG0lLy868sp+jNZNLgG7/1l2l8npvxHwr9PBzZOpfiqWnX/HbyA3bsgG
IA8e4yZiLNc3VKhLDrcVq7fwLlLBZmBjuW7NJU8Q2TfcHzwk/9Hc4Pz2ldBu5N4dlHCy+rwfIwB5
G8SExBAJwBCAyG1q5SxEIOriqGJ4j7kUo9Jm8NkR3fNjzH8PAMZc7XhPxKgB2eDQeZHjwXLXPCO9
2Gj3ryL/Rq7Vay24/XEVwqVVeUpdZiic/ddgHKJIPD04Rqw3PGiJL2OZ5h1sXOoIuYcAYzHVoP5z
EcDt326qO7iudQ1vTf+Ff2cHgZNZP1iIme8wjEPfOr0cLj4RvweP8GUIvVbH2yG2N3vJWIfNVGf7
H6XegMqILwsA0scXRCz3t/g3DApEmN1cv7JtDBppw45NBOEk+mkFPL6rfEMJzW0TANsMOml+Nb/C
kMjg2UDX9sbvuMm7EqaKEK9YtPfuMq25bDwyZfkMR1ELTxeHgWDUsR1sVG3Mc4dcUIc8dfyL4KK/
x3nS+xWBi06RpQFdj1gejh2LVj/EcgIsJs9hFk7gOBxHOCGIUsjE0klm3jAH2WWsA+MHv6yhznx2
6B/IIkYuwjOsAVsdYuKJuHBdP3pbC/zb++xTXEsxsK4p/2Pm2wTDv7ABzaUcDxqiiri4XaSGI4oA
Rk8I74Rzeph6oKt6liAW1TWc8tn7QqP3HRxv4ijaRVHZe3Syl8AM0v+Xrfv6Qs1qct/2hYB9q6kv
49D66baLBRSOxdqFd/pstFnp0n9JKJJfPfT443rcVCYAXBZGxmgCnwMh2Cgg/j13Xu1/DeVaFM4D
Ot9ztjwOaGcwe1mkePXEYfo4vANm6DtwOzsBkwqcsUgm3aUNhQ6r+ZnxOGXy66KYnWYtU9sjwyE2
tqJj6E/gZf/3WatNGenFGjfkFzYWR7U1QSH8VsKnNJ4fbABgrZy4/baW5UB8TvG8SvcJIeJmjBeW
Fmsm1YMOFGe4Rw3ucqpX+J2ePnU0ZawkBj1ZNjYteVwPOnjwHJuWBomYvpJr0EaO3Wlvc/WULUS4
/Upl9QSxeptB2e0KDET+ZYZqHgRwaSK4za+eu8BVWlDqfNNS+4HCtb8GfvjbEl4+2wARqCsynanv
WsFX+q0I0xo6dRTuWCDSXC0SBFLrpBbO83ILC7wnxOOWFn7Wd5t0LaTtQSKOFXUshc4972L78J+W
7Rj9+4sln70tEIBKneNqN1Uuiz6V9GRN1JSxMPpQDJH/nUCQIwkQgTbpci7tJFoerV8CTMgPj4Td
jRHczrRGgqZ8KQefflMrfRmoTwq3njWlpHpJhSzsbdxBK4MBnOJEnp5ZQUwsPElcqat21rK+/U68
Bs5Ei/PJAvixiIOIDuU9rwaiDNBVjYM1ClxciDL0TQC0W3DhcZUl6+Khjm3zlhs+2O1/tJ0r+oJp
Sen+Zti2Eri1iDnRpB844YekDO7B9ioLfFdXrYTqp8gLb89RMOQyEYFzIidBOdD5ybxV1E8rF+k8
uhsUcc8CbfbxW/Io1Cad+toxv/JJi5pX0Lsiuvy1wXXcgRYcQJilEaS0UDRnJt8XTD99qIN+BrO5
ZRqa3kV0tgp1Vdlcep+bMmFB8p6rOESVPx7iioVfrtm/dFL0/qjApW3A0mL0mzhwbYj1JJlBZEZA
1TPSArZJxP7/QgxA2kucLwIFVyML/zjW7vLlm5WaxDfslfZTibxmBSSXLHBW6yqijXtriMwif9vO
/j8p/1Hhri5U1e66nPEVBdnkbe1QKtzkxvldiQ4xCAXTlLPOkB5GpaVXdvd7FsvEY3T0908Irhsj
VBcGAtvCgrQgMg8nmb9NP7W5XfXmVPe6cVl/U6rGz/qrFfUn7CtY10y0My7FbLqU9iu8rpt+q2Ai
uuwtfyu4hy/UdG68A4lu7CPCVj3W1MuH1T3fsavs3L4NaPH56ekPtun8dAryE1D1H+cP8cd5TMZs
P5yBAUaFjr/uTH4STqggA7bUwGBvEoWExyItqb++99wKZbfqLJJYRnxg0cl1dBww054i0zYGEL/f
lcU2PrpsxnR9smkkWlLPct5lmnmMzP6FuuXWvEu2b2+GfufPVWcjSEUX7qS6qltw/4YhA6w033DY
BZgw7SMxUq72nd0qeztqx4HMP2WnQR7+YXUH2Ec3RQNAp81d4nL2sDLAFexZshfuxAkz/5Wznil0
0lsF5sbvC3c+7pamuzGlfi2YYH+EtQtzurfqiFuLhCloD0hkHclMztvph1dKUXPK7aDj5z8WmeRP
rm3PJa7L+HqyRO5RMb4Pnlt7a572hxCZ787r5bpgIbY8pmpcncSgLSaoonF72n/kznEM0K5i1l+V
PyKEOXnizMM3Zkg9RYeAB6YcAKl4CMZz0Y9wclsPbgvfrV58ixvPRXPF4M6+Tjtgg8bvjfKOQdNe
P8zZ2KJS43DmT8SUKd6wr9czziFCT7a96M/aW6slMVOUKEVUfLgWQ5a7d7/8yBlsTXyyWb0dUuQJ
hH04DjXpxN+4iCB5QTl7mu2k7SyK+fU5fGHqM3PDmWGsK99V/1jzRRrB7rWIONglQ2mFQKEVTlWW
lZ7mLYpBCI/QHVT+rCTe/DKNEC50FNxlfIrxqfaxT5/F+Ioh/WdCYQNiCN5yplslmjavevaREGJe
DWUITZrUvAPKSQSOq0zkH7VMhzTqnOjat4F0JdxlvoaKwwXElGZ9tf+lRfAMxV8hdWysQ1+UTCs0
oUPtrobP1HXt7jsU/Ob12pzDEPLfLF76mZI/xnqO8MWb+VrZvCX7CaQXQuyhfENllZApEW9Pr+fG
pkTb2ZL89ZOSCqR3OxkX05wU/GyzrQstNQlTn7V3Rmz2ZoLcB1cNEYKYjs/kAlbzr1oP/En03rx0
1mQEcDTB7mQZQiAeizzMx0N10L5YcxUc6dbv3FMGSU6zHXbUZ7/5DYNAQKipeLZXbdzusq3ykjZt
6LZCOdVIR7vFwS1ou64CLHV01NVcAErB+NdfPcwMyNU+ZHQoaIu5OoCwnNAIkpNPa7mfWNJ89JwY
JULwa0GAxNQme+0NgS6rcfEsa78SB3lKH6YI+UxCKBaURwTsLOLqUmPYL8C55d5XU97DkZm16I4t
iGvOgBfyBlf9wiPIGfRosfYQcEmUP7JTyClwos5I6lPjEwoHPmj57cBEATkky30ca/w5BL3NEAjJ
RdZg5kaErsXqWiDy8p9VbxuBThskrTXs5IHEp5d8DdjdWwIg+n77p/1Nfo763n1lq2Rz1Lf+cok4
QZpj1uftgu0IlF9j9hhJWsbi/X3hEKklqFk49gQ/av4WLNLy33uustqbzRjipu5AVBUz0G6FW5mJ
m/iaaJw9oH4ElKxqtIa0W/9RixEePeX34Z6ezxv26ODpflXO9mSqP81gCn0TUK3mVaII4GQHu4Rl
Ef+VLyZPzET11WoNLb4C0aKuHA0gjfcf2pqVXD0oZ3r9Mgdlbt4I5YhEOIJORU4pdmjgBcSp1hZ3
etqOo9209krMLCzcgV75unMPMtQDXaxGcjVQLgJhECxsjgotecTfp/ONGuWwe0W1zuKLCYgX04at
QQt6sO+mTZg0oTRVSHqk9ByqWtUibalnoYDHpkLKQOwqj4rbZoTkmfF2S22n+zVs0JOj78pcAS5g
OxivZM0U7a2AVOdUuluJeTaYDwbuOIHPiZGLIjmyx0N+k/RLrseXhELiE3Npg59bqj+LsbhZUHCG
nlmmhuBA3F19nkbI03zrG/js7g84W6DII7fuJPzXazvDo1AwmMu3bexX/kli2Ufw+vN5zyzLVeEC
YuJqqlm8UVJIKianNI/ytBD+uusYMCVMPK85Vd6Jrqb4MJ5YHgE/4uGjy4OttSnEutk9lOqD0C6U
uE47Mc3hQstSTM6mENxLVXH3DUNycH+rSog97tJiyfeOPx7UwzrzqtnaMg7+ECi68xY9tPuAAI1Z
Jz/wGWTBHrd0BT0Nw0CNU8C/20VpQMHVaAWjmJlLm/fyaWqBQ3FAGutjenYswx3fmDMWT3SQScJG
7OzYR0Te1M9L00Kdedc3bMqJk5zlwccNUXXEiZo82k3zUG0ZRpru7DljmCUuQZTpfP7EaHHxHsKY
zZ0kX5Sb/QTKPNYHaAIU5E8I1aS6BNmEe4Pg6n4SncIXV55gIG5q9Jja8ApcQdTpOsbva1i2P2Gw
aiT2yJGgNM93Dr2NKrZYDhHfzfphCTeCCYaWrztQOPf1wDIWevgizz3Vm0iAE8Mrg4V1QKMGZZWb
Fq5vp4oPVJ7RospcV0RNaTifPc2x/nZvFK74ijHAMLO9xzCrFxHjFY3xqmMhOnRkaMF3mjFOZd75
n9CgQYS+LeowGX2T+QUVCJie+KP9vgSb8KPm5pT59CjI8ZiQY/uk0D8G4f1UWY3Blpav/aVY0l/d
YVThei45IffhEPGWXBsfpYEfdup/oR0WBIUIMdMecOH2t+JI52voBCNhbPnv5RUcsmq2VtWr2v8Y
Hzjr3hnxBOIRxAM9M+Mpah/KQR1J+Rai9ob56IfU0gcR48vvF6ite/cLfhbRIi40ad3eRgi34UqL
13vDrqXTHPhmO5iXWhied61GWwuuIitIwPiMZpqPMKLoCImt1LElaah4h1pfMcthvNQkcDGnD2Is
knY25bOIf57ypxIOdBRw5sI5eN5fNoAq5afg4owFco10qlT130R4tuBQO/vZr23mBPH6dkpaBjKB
NWitEc6kmHdb7vcIU0iNjBn/4EeT4hTIdjTM7Z7nDif0dQboY8qP5VYAfl/uQAU6MxzvRlgy7xdu
FWgB+X4dEpIiy+AI4J93aH2g1z4r/pci1NY9pT7KwyYVigBw2Jwwf0xwX4u3Nn58rrj+uhE/S1Ds
20MBiCWGdBkU/ay6G4kJLJhR9h2Rqc7NlzdyPhp2jgVFjJ1ejBOQsGt+Gr0pTkl12j1r1HfOyi4U
4yw9Qm8T2LV9Kb6C+JvGz3EzeePVioFAGlVmu0QnXNJl2xeKN06ghC7XnrOUAlzH4HmJm4E9ZDFo
08uKP1gv8vvAZDIiehiyunbP5Atva0PF9kkB0+vE4XXQYAok99SO/h4iTQPScdhAU3AlC69bJsrM
GijbdO/A3+YyNJU+A9uSo8UL3tuV+v0vChRH+PwrH1U89YE+6qBnyoqNRUagsE2+8Ktu5Yw14PMJ
T+ZHAbjGYm7r2+k42td3FpS8XUWFSV+cctCjKe+X1FKs6/ktdqJWsh14XqFHbXwBO7zPOObAPj3M
cUpIGKM6V+qX0V1BiqbxujzV5X5iwvPz60NDcQCK3cUAYiC9aqWPRta/e6kH1G3ZDwmDsEVextAh
UwmNC59olz9Hsi8Gf2+KCAYos0Yb7XF1KDsa6pqvpRaZL910ItQKJwh5vezE/47JrR3bHoSE/JMO
w0IlYlQb/FS2zNrlkkhJECek34nNIp+/19QSACQSlGQ71nDMYAIiPSOz4GBob9NOG/R4GPDNxdQc
ghbocpdvaExh6WUwm9T1vrTdWLoj8eCVZxxtRhNYRqvPasevG9gNoX/oQiKR8F2RJDhuBJJjvVyD
xv+H5TrX9P91l4zZycLHn8xN/97/xhp+faV4qBe9mkN5JeAJ8Bh4mToxmAkdk60okJDfirsAFPey
VRNHdYKIzjhD6Em1gX8Mfxhq4wpM0ZMQAAGma2M/l9IgNvGcZv3T3g2iRXMzmXIRrhN7olLFFX6S
K7E0x7qWQ+Rqyf69TWLKXGxqIutwYwQbfBnoc65r1KSyuBs289JMTrORa5wC1R3yjoDQM0NSguJW
Xc4zx2Qso6ZHYmPY3JDg8/qbRxa2J9McpWW7hTNfnCX7aGb3Q/MzCjwvZU+ZyuppWRWJHZzt8z/X
mARpLh3FwD+pARlJbRR8Hfz/cvY9ECnjt1TvoNdK3FjzDJX3u/W6Fi4kEo4qRXgAk95I8VGnw45z
ZYkPan0MI6BFrsjYrlrpEq60ffy+8qYzvC5/h42jzbkL3lRJ30OGmeAriqr1JLgtYn4xCtlZPeKq
+FlftlVakaVJF8tRA8ny7l8FMoS4Y+GtW3TX3lJ+eZBxPu6Cw1u0zw0Mm5Iona84UhPFj/OrpOBh
1TKsaWwIYh1RgjsE3M9gg10OEtT1AdHlz3HOSkyzyj70FjuuI2dzRTGcQekQhodG1XIe9I5C3//k
NeedNbXvHzxkfWEtGyYGLCI5H/8vaTqmFdV1wT7NB8rwxuIVWIhT+svUx/RPMBqtADIh9gEltr96
UL6yyzulDE1RSkAx1rFqYxUM9SJ3RpqIrZlhsai3jSnY4SDZ/x4DZzZMtSuuu1lykoO6wynG6xaj
Jv/9Kzf60Cy79ObtmC4md79zF+GsVuUo68ZRC8OPsIiN8vzHyADa9sZw7CHrJubahliyYecaqRFs
UJxIF9z54kL74imlvqwYwvxrbmGTBXOyA5uiU9IGZsrg31rphAN22mR/L9ww45zkA+fpkDM66CgK
lAsqhSnYMYX1zE9W/1Fp+9zL1wC9IsVCTlcfVKl821xwBhvNcDF+HymtjwrC8y7wTYflAvTHlXWl
U+7fF2brkUysoobxLVejjnVNMLsKJPVTJdLtc1l+Fh4MdkzcXmcjpuqpxoskM72+4GlbhjT/B92D
e0reFIR5cdFagohDsdT78vQaVEHVKIlr0XoI9UdH5kcJFEEef0J2lnjz1FQqIkpmUXzP+K0zLUR9
N+S8AQjB3f36JwkEL4nsZKhGU7a95vor9TmNIE2zkyXBkV4Lb7rOg47k7NvypxTc7FJMpL/yuBiX
pZ8vBQbceSNnxAY/8PYXwWGdJEpawlNmB39DYDulYgVzun6erWyyCnnwy8x56ivH0R7pP45SCsS3
41SoNCPfi9o2bGXp9ycsTpKI5Sznm7I6zSki8nYL5CX+L69ZFmMWa0U2qTM2h/5DAyECD/9uUs1/
HKIcilZyq6kyummcaIIsa5+HiP6ehGaw9Edy60pmI+1/PdaCHQKLHMST6gjt5QidKMnXHTu+xmcK
pBfdHl80mYUEU2tt+KfAoLWZg9YhcyLPJ7vzHX92a+JlMe7EypA1pW7dSdO3r8AOYAr2xA525MM1
FM+akN++q0ZVcG44Hgv9vwR6u0Rk9rEamsz2L9U3gI8mV6N5I766bwsq7MR9QaB8AKgvo3MWFAmC
gQKTNrwkXmtV0bS5vHO75eVzkayHWuDn+fIWURsuZJBbva/QR1VEqTOoXBHGRzkdPu1i5N2MDep8
cgv2k/FMe+br/ef/ZtUPTxgNPF6y1/kfUyuLoDc26icjN1elCuZOjzWWsjAJrF6irp43Zi+wYWzj
RhWTkI8JhnShbsqg17osBnb7kPieRZaJlZB8cVexYVV9NgY/ctLnArBOluHb4JifEjeyW++3L48X
1b2vr4ulgTdb7ivSHWwd123j+0oI45zKo5MyxKDpf7QTZLFxhhXHuA7RvA6opgVBLCimrAUjquo6
d/2dUylBmA/BgzFpZ0Bgnly+npzfplokJW+WG6SwMtKRNY89WWyiqFdVTNwH5kOj/pi5xgViQNe6
RGvgAbCUDfmCXzzReX+LaSZWzL6J+kfv8cqFi84zBLnOeaq18hE7Gm89cNOcuFrpRYwImZCoKefk
GHmu3ekw90yM4GWtZauoMpSIb2Np5SN53aS0PC9BKd4aU8fN6pf+jh0ntQkqhqJjBZERw2gXVHQf
ELZ2xht4Vc7S83osdBEnaY2BY7pzhdYivTe46xk8KBvkwufPj0MjYcu/mPURZFRV0jqD20Ns5bPV
YOGEAJZ0S6mGWoHgBSXf9sSJi722hcuIto7ohpt8YBvVIcfCalVcphV4+U2U+1vZg53QXK/PTvWl
/6+1wQjjuIgDn4qaAgHRdxVdoAsnqlLGWa4KLxdHLTdlV27aCW/iTgY784gSTJPymV+vBbycdro4
hOu7+8YsYp3a6bwPZf90o5k3TEv2piXISgxBp3abQDEb6ppow6Ttm74TTpjZ9fvjPvWPIXljxCuC
CXzD+cBar9vBnNPZ/sXVaF9k3Siimoxn4JEnG8gVn8UaDn20YFiM18R9pZrFUx05VilqgyhDxg3Z
kKlcVgvAEPx6HZiCefUwrl6K21T7HzhbJ4wOPiFCgaNV3gi9K2WwKp5hqnJQSI6NmlpEd4U9l7gc
0OHcPXZ7hYRbIdTSOiqTCjyNH77Cf5mxnHAtiWn03sTIdnpGmF3U7CC7JIDzK5npbKsfpTk1DyQ4
d/Fa0jnIWz4wDv9+2K/KNiNAJYEyMhTwe0Q54gusDCjhO9gKked5QXYMmSvbHygQpXNi64gJzFSr
zTj6zpZdXzrodt+UPDb+4Ut/38gKbI7p0REMK7Z/dfOe+BXKQ0gEpe4IZQHLfVNd5kkIQgOr0dOn
OpHld9hfUghS9mLxKuKV/jeepPtVnE4chqO8Miq8+knIjjhElMTS1HLlh4rCH1uqayYPQDnk1Q88
akDHRJyg1N3kbkdL2aULDYDToj66NH+FX3+s0P0gfM25WQMJQ0q5rXXExZqMosJhR79k41Bopwke
YozLyna/oiGZK8t4CG28IexM07oBVseyinR7dq9qrpImlWb2wN7p4waqg8aar9LZy2K8onOdJp09
qkfho2ZxKaA7ICD+GNe029JoJnvh4sfIytW9C8mdgLVMD1xnGw49lj2L8reILBeSSG2HRiSFb8T3
gCJnjaENdg2RmOJAeVq2N6DmaqBeoFs+GeHmQqEK30YPm+fm7uWiXam1LvR50cZ76/bTYf4c1B8z
DwQJKEK/wd1J0jsg/lUJFRfFwmjOs8HLAVLlyK0zES3oTSaPV7YeuYX2d6MND5ckbki+mDLuOy+e
s7Y4jubG3JpRBlURWyR/8s2sjlSYntYZ///OaMmo5COaWjaXxJpAp84Y8UliLy1UxcJQe8i+B3zd
OeYrApb+KPaQyR8Sr1HBrmKkMVlEc8GH7zcZLMRh/x+JPSeLINOv6TYcnB7hxWcgyxkgQIpSt42h
RXJeLs/hH4R2ZPgwI9Y9IMkNg3oaSFvpiqv2DyzP73akGx411ZUKKJpPRQe+lb4OE4LOYZ0VSA3p
WtwyhRJnvvepGDqPXZlXWeeXX8g1URke1CioYNM2osKudiiNcnj+6SC0n/irP4OeJiDgEM/Vuj+Y
6PmRqb4Ohtvydo8dX30tUEN6d9aTPwzoO6hUHjViCcERYB22dWOlD0w/54n7yn+U67AP963XikPm
s1LstUvC3d3iq5PDkwfiHeBG1SC0JjNwFX5WkRd+joUQuNU2OJ5y/8/oz8puCFbcYIhZETnzH6O+
fqXTfnVFVRI/E7WxS6mHndn6OKXmLqmnatDzP+6YHwWjuuaAQbMvDHSuCjD+BIAl9YxLGl0DSWwW
vZ+Fu0jPiaOEwB14a0ylmPOInX6LbfdGtq32ov2Cmd4MvTtEvflAIqTK449+WGquGLY/W5feBbWH
8xz6DPYVQIWDTByC/+jShcXpQVy4Ytdg8JSRjiP4GbHWi5QGECuaBTro3/7ZYoqioccS6WDAWoWS
RMysFEW0tOLVCT3Rp3OBiV+AmGsCnv/+L+pqEXDynjt1Ceim53M7J7qo35rE/tb77JaqCnVNQgCz
6RKrEjriH4JL0gEcchsz/ulhdTSaWaEr8DmaffFqwn9rrTV7FswTYlyTix5cXeOAd9lspdEnGpTj
wQ79njeq+yLM5CU/FV2E+BqJEyK0a+BOjEQNc0/xq71ljRpoOnph1C2d2iHjmo7K7nQyprP0qPW9
o+smhcGw8mXKwpLdAFwv1cDIY45LdXIqVDDDr9wo1+0603PQ9ijWCYdnUeaF7pbc+CoDv9MRWDA2
HhtJT1W9J/qPsQWB2qdu3SVzbMtbjUofP+JMFg1A2bHEscmjhIbKKQmZEHS+VCYDvHDqI4YmzTqp
gvwCGGL9xXMs6O3Yh04Co+IxrWJobEzRGeVLfyNpgufZf1u+IhM0Qq+n64a5DM2VMDHhdhAeH8CL
t9wvgnxnmMmmIdjSElJKoxgT8J/qW05lEyer9GQs2nroEGtp3KUzDPhcW82K8jFVAkVmJhKIV9oN
ABPkuq+mGu70uch4ZzvtfqhxVjBDOk581xiqkCwO1Xq4lv5rA5PgbU/mUZ2kKLjOfGZAgYo/u+uM
qbo/WqJINOx6fDeCm/DpOcAY4O2XIs1jo5AwxezuaTWhshZ6haKOQGdwmjduJ4g5iM2348tBTZl9
13y9wPAeVJ0NkpaL/5GUeU7olS4AigN2lLfpynAfkeS1k5jJjyfgYAkZqbK1XjNDMRJPvQqYkDmd
e45U2aW95B+6petfrAocbGuJKxK94QcJvSTJCQ5jf/28dt1GxXxGVPAtGTpQaxWqNqmS85pyl96E
eNHGqbKLHpvDJaTBtGsedVdbqx96W3K2l0iFEPJTeRu3FN1K4watHUSwzjQLW8u/2vGbKq64ANt0
3e/dfueVEqub9OUu9VG2VHGXbrd1c9H46vxYHXXoql+YB0iipvhjqpxQzHeQv3dw8z2b3w7OM3BR
SMJDGSdee0JdpCy5E2D5SFjx6Pl4t+OBxCFlY+UdG+Y41kpV0BEOfFLr0Hegs4tYbRd2jEapLl+S
caUgBEQTLqOybqrecI/w0pLdcO2NnnsUX7I04i+JfdvwyZI3LTxt+3bFJKRhAS9L2MGeawzSXAMB
Au9kh5yfw6UjdVoOMmyfhe0lFEO++sEPKfoyY4Gdj0dG5oTGbAWIJOnFfgL6gART44gSOiL10Vva
rpTf4OvwVLGqbcsHkcUmiSzt8Fu3ik9UI934vyo5FRI57sCllVLWaSgt7wamwOIpyu7hbmOc9gEn
wMNyTr+MsWVQyWW9bKrIO8wNLWgHk6epi7YKc8xa79QBkZICYVtW8lBXGKMHNC2nfgIJCENZ1Bnx
ktqO//Ff3t4evBpQq+93EULlrIybT2qQOnYEpzxFQVKL1HGLpr2pETULBS/pdlB7bIbUVNwwlbJ1
QOOjEe4rSnZn2B1N9MdBhDZjLFbdSx0+mwcsyrtq47+bhwkwIOLhRhRy5qrdWb2yFXJLJJltNp92
2xRbJwDNAIojYQwl+Nmj7VCge/5oRtrtqTnpc/gwifTztBWvYz6r+hLa6tLPraVS2XL/zR6NUKU8
pj/zHFQdPclFtH21Y4WzH6pTiWFOKV9SYrdpCguZZavomOo3cE5FBE6PAh7UOxhUefxNAW5jqcnB
SWTN/gIelSILOm9r4kusFnntJMhFtDliaZD6T+xKeNp5sFrW6CxGSxLeNSU4O6Zlw1XWUx4YCSrO
Lm5rikiMqrxDV11ARSswSLxL/a9uhGlXNV+0kTc2UKTf3Nq9W+4k/M8KQb0VIyfiA4Swl4w7VDgX
uCrywdO99csqxxVSXHt8VJy85PFXSJw4ORakx1S63qVqFTSbTkjTRZaADLszRDJ/jbIqInfg0osg
sEJLupxYwqMJgzWFkdbeBAziHZisZV4GMVh4yvrIB0AC3UeyD9SGrYltEQs1ZdomTmMg0J314dR8
2pFFSsgiAvxDFDb0nTpwufU+mCpKm+5qym59D3LObaGAN1xguq86IMXo7Bqs021UdHdxHXKO2quR
SmMa/0moc7F16eZ/zpfJSEL7c3NrKYtBn5gWC+7ceB6QuuHyu5MHV2WAchve6zl8G+K9Ptk+poWe
mYom4+/44IUm2JJSlKBZiqXzPZGOlk01i08R6PvYG7Ao38A8dQqJbXiVuaZPSlS3WUkVMWghpZKn
tyUumJk4Rq46uThFsZqhDW+vitkV4R6W6Ao7he/zDNfAoDRw2sfktt+V1huqLbRyBAINg0lzXG1s
fRl+Cyqhb0FoEa5kydFPipEQg/VwjJCd3s6Vgp+sozzSuLvP9VVLcJEH8YmMImlyiwrkoPrd0ZHF
klzBiOwjeXDoO+Hjb55kPN4aU9SZXz696bdA+225hMbBK7SymlPMoA25GezLHN6V1cyoihQHX3/u
j8dJKqa+jp0Y6XylQuSNxtUMUb9ZpWx++VA9FvpzM7ZW73TcEaYNoUjhMDL6+4mr+Hd/XTJG7bgR
8oa+n6xM1GkVSlwgOzxxEo8adzmnFUwtuNSISkCEg6JydrwIp5VZU42nA0JsNdjEgVK+fPJH7q59
PNOMR8DEWVu35grRoouDDElgUosBVfjHM5R0umlK22BuGaHTps5dyjUH8mPUSUGRwFWb7DbUCMxx
hIIqq6nyCPOjq0VeXOevd3Km9fKHZDkg1Z2KUAoEYWjbSf8DImJf5GcQfsg3q2hW+oOg1Z8zMuGk
uymeSwkz+3E1kNFW4R0uNaiEKjBF+YZcz3wJ1pZpV4+TGZEcBKG6c3QzUE4wSR9FFCdL7ZLuAupj
GrsuXcio3mXFY5sez+mV0zDR6Z/dwrDwKFs/wh9giuE6Bu5PlxXeP1QWCfWwrUs8ZqVnuFqIps3R
q3ikRtD09NMC0bveC2tNPDYtSjfU3RKNhGs8Kw3h0hBvt+9eCSBpNiSk45PmWsayxhcmRl5aUo8p
sXDpRrddthU3x8g//UdyfaFvCNqKzKdaYP0GveN0wJwCvh9JKHHfxdDdK7p/Y3442oACLU89Ctaa
qKmhBM54u3fX3nHpPOPo/7a4xNiAE0hmUvyzKv2bZ+ImUI9F3YdEcypr4sUm2iqlvwXj72PX3mwV
EAQjS/DPmsygClDuCtkiYbm2eNSlo8jv+3FFExWs6SI+ALkbGxgiXEVWTycttD06oyEuOZIjfcw3
nqgZckPJDvkXZ5HqwokbvhD6QpTp8iRdQSD7ogLtXC39uLhDZXzZTOLYaQytFRZ/1Haabc/Yp8/w
YwnehICfbqgRBXWVxJpQm8uglT43BY6luGZMf73SILYQlL2xH1+sFB6WlTQKCpF4L5TwDw7Pfdfy
9nDKqIZQcJqNFvLClYuQVmWSwsnVzX8cH8GBGNoYyfuzT3X88resFc4OJnXFt9MLrAmAtoLz7Cho
4z8Nfrv/L+lMZQDCrMuRlRdbt0lbaGvbsG/SoF2C8F0UXlOhhCk/WDM8Vhew+9CMbnoYUiZNM89x
PUgqSxHkH+nu8vXmaoskumiQpWf06rcmx/Mj0B7jxDFI+z9K7hgPXXLDDZ3H59nm1sPp9ael0gkU
laEC/x9x9GWsFCpUSguGkvpUBXzKq8Br8Qxwh88ukZyy0+yhDEnOEJqVR3IyjOBhldFBsnSHQNI3
XPHVIsJhLpRfUHBFCCAvdiyPOeFVKKB9W+DMbIHIETXEISzI1VgGx+GSg5l/7e1N9XoUn97KtJJf
bWeIAaY2uYNS5fEjOO+a5FCjv9ynIWBM78hMTgXVCOAOu5WUPSCntkFlceEOfystJrOVUC4N9s25
zDVmAKIHztgk5zi2kBsSvG1OoCpUc2lzNjy5VbYurnZXIqYZEpK7LQP0uMY9RUVH1CpbjpRxw8b5
/XWUCE0Wp7HqTttl1DNsfTlpjHOR0vuIQTr6ZydFyrBDGI70tRkG78Q+h3Naota6ZEvJlpm/D/Iq
WdP51iO4/nKfBFUkciIojIFE6fn7441gINzld2pUIoMMy3Q8mRgIVjSLzffYz5MHO9vHKU6fN2+r
YiDLf6N4Qgxe1aEbqaS/IZRhUoAap84viXQJ/OYIBu9GvaLX8pCgjqgUtWe4LIxuJ3yC8Zplc+9m
sLL4c6tEsCcJtUD/rOdBvLmHtqkFbAsJSdjrMVcUoKcqBsGTrNhgRJdXyB8k0AwM2BIsXN5QQUJq
8L+BWY2lF9i1v4dOq3vI/VJCeJd1y1DP2LzVNhSrL5TIr7Q10m27vpUH0K7xw/i3aPIVPeKVNYsi
6Hp/X382pFH8+O1NAMbHeOTxd/F9IBAUorZ2vOib1AfUCwWAa39KB8K+mA6OQguyOt5WoDMNoEbC
6Aq2W774VRhwDME/sE159l52CtgW6hRo0AsFXUxH4OLJyxs8UabFKSFQYZ/ha7930d34RX79xPVy
CbtpjBt7B4J3jexcrQdbpST9/iP408Cm4KipwO6VuSLKLGJkzAJfn41vIEzujDMOj8QFCKLEHQfL
W1hwyClhYPw618cHls9HZbpjOMvGpIzwgz0QdQzPbGpiofuP0/Hxjtv4zkQRHJMpyEaiiMaKS3+8
E0bbhkpqvKLucyOSW97YIMHXDLw6Ls7jEQOr/3DUocJc8J60R4snfzGtulKOH/5W/kjDW3z/A3v2
7766iCify+Kx1rYl67CEElf/q/OMHf+LUdA00Da46KtOT0vU2gOSiSAEVic4O4rhNCVlDp2kbSdb
yGSwDz8JiBDVENlD/LWLirqDzQV6F6eY74JfDWbWb3ifXsBZ9RbHktcsbJdWN3axnqW74v9SzG4a
STAwpZM+NkU41ekExOtJfMG/Uz/L7IRvUo4N2HSJVotrwPzRYEV9IPZu0sfvoZ5T3YJNSZqI/jRb
ZmIP30a5QcEElP4z0xVjuPS5tQrpt28VIWe/t7M5pDsuvlOfzffi8/ndH4iRNVRyH1TJavMxYXeG
zxK58SfYHIK+sRYNZJQPDNzppdYblUxpCBQxwTYcXTfq19s01RzKDoiny5Y2qEk2xARFCNddqqFd
wbGTmh+jxKNCKx8RFwGQtdT7MCtg0Ilyz5sz+8LhhmlE/Pr2+kTs7e2nUBzeqRCYo0AGFXy8ej2h
P6A1m+iMtPNv3OHj5n02WZeOqHVtrsbQX2Z4fyi+xTM76crH+Ai8cIr7rbB77JXJKeExtls6fqxh
+G/nvV1sDL49F+UxXqNJDuqxwEvdf2PoRhVeyKFSuyok1JWTxzhoC6vv9QHRvmEYWmalI0gXpX64
8/YwCKjueOEax8f1fmjAVFStpzyqXOkLd1pxEMD8zGVYlyILHJYXYTs4OsTtrEsICoBkuXgcx922
T+dRPQEYBiQmNkp4Nsd8W8QkKujfoXQ7jGTVJPhCLgljnQO9JXAMT/OH7tzxqMh9roYk0VMSRra5
90Vghm+b/btE9MXe7ARelydPEEQaqLrUE0MofUh3aaaslZyPUrPdpZeITKL8BCGGFASuhb8OucFj
RwXq7FVR3RNjfTp4cg/17bb9r0FYgRotye/OPaRi25Tqk9nYt5DrxzC6YW7cKsH9VooKHQftLk1F
TTzjpkeJIZZeXwNQeAQatnN8Y0bf94bAU7sRgx/ABSYeKwHMzlupH8pK/XF7o46SL2Ju8PZYuP6v
7yigI31vso8b5gcH3V2uVemOf80qT5EaYkBkrBGNV8wmNMNsl99plkX5b9O5PuLLU0OJiLlRewlF
k9wJjcN9ywM9L+G4wYBAFp9Gk6tk2ncBOyZNXflKa3RIYHFfhjzeIKf9Jt+Y+TwheuCvd9ciNjxl
1Cr4/0RFwqWFtWU6h0IcPgYb6QmuCkh+U9MJMDECHlOksK1jFChdKaHJjJwoZ7+uC9CMYKeryuwR
vBA6xVQX9ckZ0sYFnB1HurDY4qOI6exqEj+l2R4WrMR2BhUop1BTgi+meupT3oyPRhKQOp7sI+yS
kwH1asA7+AuJa33G30X+eLzbquOZj4vdmk99xad3gof02t8KdmUPqC4ppprD396P8uDlZw1JIRwU
r6SFJb8hTWpIimLOBh0IuEqtbkwvnyFzvLHSsF60RLTqGP+krW82MgxU6i/hmUcbW/mxEOPoqyzn
xxrJTM+LUEgSdNmx4rMzUGXrPka7eq3YZz83o2PdB88gnM5mrTobBcNJCkfCrbn/8yp8IeEcWWFG
ccQ+C6Gs5qCH2InNpebWas/0elJQI39kDMpIR2VmBfl6Tt9tO/5lq4GRia+owcYoQyFAsczsUDvR
c2ZQ6zBACBQTZx4FO25Zz8+RBBNaw1E5N4MwXsXHLQi/R79pAWtTz248YgklwjRvp24EJBQpN0B7
vs+fwf6Ljt5szZ6iXG2CL4cysIYDOFscQHPgsgP0usbhg20K0lX/onRcubiVh93LkV1AJbxGA1dy
rw3EJBqDinStmn6gjcjv7IX1CURem3TyFkNX1UzMhPMFDiVGN+l0bA8mMtN3yGYtn0Sy/JqONmhz
shTWgKzSukO1kUykfPq6UidEm8aABf+iBiaMz7ZnL3w8gGEYQWOlXSUX9i3x6/CL+MbB0ULvovFJ
KlOSzdDZf2+UjjZhuLsMLGOzuFGoHOTN/1sjfEJSiSFwL9kS53tmqF12sijjB5JYnEZYki7Uh4oA
GCzqSlzpFKgJEtRM4QWIQ4EguKcQ6BkeAnQjkx807t7eF+WJ4DBHmtVJZqTneZswX6aB90qA+f6A
VFIdGBudDwaEed9HyHiK4GgxnwoRpj12ZHPn7o2Oc9TGD1C+3hY1cgycB/dhaTd8iXgXTatEdrEE
gAn9TzF9P0ufB0ymjXhJKClQhzJqsn81pGiNEobuqe7lsjucQwTq6mzS1ceGQZwSVEcRNXyr0kO3
josX67TrTc3HPSTh7NSEFrgX9tGxBAQHbQI1R8g+Uapv8Nx9CAzFLw7qDmiI3KJlz8T6avHdWouZ
J59UBFlHSrvz8bbifCTqmigCTEk0y8LBZC+vqF3Ol0suQFR5MXecIJQEENx5X63i88v+zULbAvfO
IVsi+btNGBBbHOA5axwckLrlRuy37JrZA0rszqOrhlF7Nsq/RUBhEOVE50IukeUUoDEO2bJ7XHXC
XkSTHgkBBx8RFwqXh+VnmnOfGBHypfThflxnBxFk0Ai2K4MoOMBgUiyK6eZEGZDLFXD2v2MuA63d
uenAZB7XZrTllTmr5lu6DUzQTLhTb2Oe9D12TyE0L3P8UgUgLmsXowsaHo7hQJ0owOWKc97wKQ3Z
c2kHB3Dud5g/cTzdH9JAbUoD38DCuWQYbCCrJFG8BAlPYyBdXGR3fg/ah0gY8hVvXI10jHJ14/bL
eSPdbuhFX4cPkZF1MuvGyjTNohd1/o6hBI7s75YuN6eoLum72Br8YsX/N6rFYzqPKuTRGys+NX3R
sZ/j0qZmH6zKcrF4hhjuTg9KBDiEX1TinwymTDnQZSpC0/0qM/2dZxSuzVYP/7UwDuWzzsFh830n
jkQmJxaewrVPihBloU6ruWSAON6QHrgStFyHcnU4CYM/zjogEdE/pXY04aHTbdoBKlLFNTbT7IxD
7P4sqrQk5Ba1d4T5iEKIkYYPqV8TlF4jjuONsIdg5osemwL38pTAoNgMBQfQ4mCFqLHjaIpGro+M
SnIuKJ9XkYhXYmLI2APeKaCQfFVbKkhpbR6Y+PR4GFStMBRR+VHMQ6H6U16OTUgxqisma4SmySo0
YagA/mH1U+THHDK1HCRTwyYgW4iLwtsebKtqzUX7TU5pQ+iIJTOlRFhYRmUUnlq4Y6/soxah+C1v
ERTLHZ3bNcvb+hihbbto28WYhOQIao47Bxo4nJRtKG24dHKXrLFUFcfenEiu6W1MD072xDi86v+F
M0SmWJZSzFn3zojjj/mxxP8GFZXG9jFtFHgMQuJ7iUzjMdJETyB/wqwjAcppvoAqNyIbLqqgl2OZ
g2uu1Ip/qoqcKjL9Q6kF4DRK0cIDbRS7uvN9XUpsqBog7VWTU0Ew0JmftNACIHdlW0U9oQeE2jR3
AXjt/pec2jMOKhqXNvZj5WkZCtk2S4yTpFPvxjSsKCZOA4d+z9vnPz9BSk1TfiSEW2636zNhxNEP
eC8VZ/o4EHcDFZigG5oPaLHSdbzaS7Bxdv6V6kGQWtnipI9F62zspoxRc80PiSg+dt9fj2eZVvVd
m8Tk3zIMeyJVnojPmzIA0JzgS5nFfjthv0oVi9D4xl4yFmsHN/lUf/yiB49cB4aiQyUcgs+s9Azs
3SndbBZYqfmuy8XSmJcUmHavU56JIID3UYgeFuRcQ5TSdsm229RJa4DSVz2f2xphnWT123FkgBmn
Zgewwsl2xV4L4XqNOWT5zwCAnbUaLgp+9FFdMEd2iJpNSqp/FP4U1gEjepW6PbgWK9pGPcDTEQpk
ppjlgMxaOIVxF+seaRHCwUchNN6nXLdb1qIL5xAk4yS6bWm1RPI4FcoMMdb6hMgoEVuqQII2Pmbf
FBVwLxivnaJvPn5bpXbxq4nngRIlszdim8BMcQjOsySN+525tI8skMUKG0c1YzvyG6twP4Kfxtpw
LXlp8oInEU7JOLz0x1O/Vk/CfcoGode769IJ6UiIVG9H+Lw+4r4wHR8Zzi1DPFiQIP7ogktyNLUI
Cg22tYUNFqzxqkWsDiGDTjE2Yhk77rcns24NUP3fppMudE9Mts6LzwCJi+8gpxH1gUdrhwUpbw4C
NgoEh+XPdhRIdNpjfi+QXfQeslMhfjuST5JGUB0SPxtMnEHP1VV0OgQQgsizdOuteSSI/TIOfwCc
7QYm7GaFDvwFTpRoQA3+D4bp/qhuM3Nl84xiw+LnQcw8sj48+ie2wm/bgVC8QIVjo9Sw1TrcsMdi
zXjWq6iAIE02ucKaX1/NjBVpKZgl1z9AY1APk58IEd7wqfCUi9k5zp9BexwCoCPvEWyy7Mdq9DGp
qnNVxdIsqMX3lDmLH0g9ouKP3jiFyFGVg1d9UhYwwUB1sxeWv12PcRGDHKyl0cbF6Aj9EwyLdD3b
QiqhFUEkprrT+VBQWuiiNO8PxeMznTdWL5V5pCGuY7T+UF7bBVgsWZs4ZE3kRxmfpx2opeozDGUo
tNHCiAdQPu7oH4v8F4TX8yXH5ZILGNzhuI+fw2aKRC3tLaNl1bu2jTpzXCpq04FEbKunSJH/+v3E
y73Lsf29G4CQAjViMKClzY0golj9NZ2TBsNJM5vHASi2jrm/rZcLX71KNHKXtyYtR/67kIiOW/jS
jHUgs3rFJLBEvJe7xDA0KAoH8l3otOA0OiVpRK9R3Tn3CU6ilS/tGV69ITXHbfjn2VRMA7vUBYTK
9Nm+E+WDQHJBljk4MUDRA6ehuY9cIAL1Cfcc3ZgytXre1gmAgyJmsHbeVIL53WBqkONd7ugvVAtH
gGxY5ZNRwzn/IDCdaXHnb9Sx0+flIiIyEYWx7KAFqHuGziV8WGBduWXLYr/l2xgJneNPZ8SUcASa
VlsYETcV4Dj+41b19toP01IVckYRgMkCpsL/x84bENfrzRkDo+fIq8hUuv4PWzAntgygLFyp3GcC
4GkkQNMwfuU7bTm+LGm50kLUwE+aBmAOJkYk2IqAhOJ892XPgCU0U5Dzpog6zzgqGcXIEamQgfzb
G+vV7l4uuHeDvyI9CszEdDuEjfxk2p/Tx2/YNT88xmheGDjz6LBbuMVAB6qDKp0O5yrg377E1pVe
zwQEHVQa6a3fYPgfNJq/YpjLeaDNPjWHkT7prgAs3ZBV3zmokXCjxxdt5GfnF4qj8+UjlV2gde1u
kqT8Ar42n6XjnBrFeIYASQ6HNRIje+3VgXyXdb+ls5iH5J6OhSU4UEKOQu6G0eyPisTC7H7FYYqL
5eGJCSkthkBJlut9tD761YbIxSybPPmj22gDi5tFbLa6PGwkQ45blf/+q74H9UuZSEEST/b3p/bX
cjA43r3/9BaKdP53SKrw2zunujj+yDlSPruv2m48n51qWN468KFR2j5rpnoXMYKXxcjCWBqwhcSS
28QSuGSoRVSYzUyVTgRcGsUYR6oTf+PlX9jJ/qVuk26sjvITXcqbspPDDRIHONbgUaF+Q1VxwXfP
g+a4m3ALuN6Wa1/PcAsG+/yySeleojThbVy6WmcJ51MC0lYVWUgrdt2VdLICA4zqVKbEk+obhWN7
S7tnzcBflbT6HLq9JvFuXafWOA3dsJmKbEyPzlHM/7FuFlW3oVAsuF4GculCYWZy6AyO6kEnOB+R
zdQ89jkAI7hkz9288YE/yEXuAi+EAYJn5l3c+OEdgJ/KkQhKwNsXdKdNyQfJGiXiqOPv9tOa6Lc1
jCkHyoMw35j6WRPv3vcfN4HxElfgeLhvgpGOJSC+DGT9mM7yleJgUlVSb+GdgBjCGyyRy5Qhw2HR
O1uU1tsfNU0ZWmrPpUhq1czHBHKk54Sd59e6OaPr7gpEObCmeBpJIAFYNuEvYoHw71Y/W/ISUL7u
4/DOM33oHa0lK+xq+7R/XJu2s8ZWSrQeyVIWcEz1yUASMaaTxwDbsEaElV1pTrSA+iEak6urXFwe
5qbBNHSmEuvffWKfPrnK8zAYqX52BiYTRHxyzFGSJzFnyo0MnInbw2Qczn8BTX/MU+u9NYsR4RsS
jz+2qEviwzokrqafNL794RYjVb8YyKNoM2qLfOr5zKTreIwsQl9ENUXBqK04yK0mzJlvFS4LCLO8
pRMrCpK4AbCPxD071MKdFRJQK9GAhcW6BKpfhRnuFWUNAGR4CzOK9rrDaLwCNOt6UCH4NMtLYQ6o
W+bdJKulZdagKnlw5UwDmWiBSiq2tt+fHZ0ZmWhmRJHLM13plCCM0tSbYg6trWv2jxPOsf4e4SzW
t9Vt/QMME2InsgaGOggFXIJGQA5xqCnuPgFAuUzrtt2r8AhLUzHSBNb0f6FEZ1iB1VEhIkmY7lHq
8O1SiFj3EcSkYA4tdFGTqupGnLoGmdD9bcvHR9aQFkHsdcLmqtWoSfGZSI7xPTmqnEtun5B7Yi5W
GD4bFPBDpVOIGczPReRXCvpMaCxv8/mTxf3FoWgvlbjEh+6Aui9i1Jvw4vTqKajxxEpgIQskt8oh
0vZsSEOVKs2bImSA0mq18KixUhcUzIhU7pmo2oSDPahV3ipfk/qrSHXV0D6teT40sM83Ykhun+Uu
4WXvU5ccv1XG3N/RUQUYqosdOSxY1sDNCFQjgWFqPeD0Pi/+a7I18XEELk/7Nq6qp0Vn49ptqqsl
TZi7lRsS55+moz1bHRMSvA9Cvbyalr9VTyBwTT6vy+e8CwfW9g60M4ZgRRQ7XeAa7Q+o27Z/xGHQ
r5UyO6pjGoPpz0NBQEhKdYOvAuYu2CpfgPZODWqGpcROT8wDXIz2jiIJfpct6J0fG317ij/Wwd+m
e8b4hsyLhcbLMmVc6JiSzGw9efplMg298bdFUfhmfDD4P96IPzkXBcziZsTjU3rFW7l9KRhCtxMi
Zl9ZbDoWdSD6O6kt0vp4h1KLmHN7vWYc1IXUyp+fJfkE3rILD3+KqhzfF6hmpBN+Yu3QT210m+63
xI07qsUINxvgs5lWT1rIArAuAr/L3jBXFAY+40YPnHN1GwSpl4bcqaaNunmiXj+pnE60g/dFXesj
UVRbgeMhhmXE2p3jS3HBb2WhjqB8UGyeUB/OPdEI0a3eFYVtmT9MxmjmQy5u1rk3kg+X98ZP2cO6
neq3FgkGg49UAvQ1p9paAUA5/lDmbgEWBtPpxpYHqRkJ1C224rn1NeDppTQ4u6RREohfBNBgnF+2
FkZTyg54cWAozbfw2lU8SDiPxlNgybxuo8PX/VhsBBbBHpBsS+FGfdWlshSa7XDPiPAztauDGoSc
6zDeUxPDaa+ga3Sn+KOYB0m9D2kUKKQPk7o/N5mw4yaSxUjyFl3wIm9WtptKxsu8kB5bFY14vSp7
zT+Vt1tMgIoDyLCa3/VXzsJvlpa+l52r0CIWM8gOa3fVvYMUZ4JG6mAZWeBu+P2c/WcGO2SIrhSq
xJCFCF2BdkWJtro620R9Z7eypinNeo0Bm9hqMb2a/YlrhDAbrBCa3lGgYUTu5uibwCHkT8bFWwIU
WekvNLLuWZiz2nG8YDIJCaL64m91SEAP9v4e+ld/8swKWUEenXbMNGPAAkh/69gZN0su4OGgOJ5L
NKsqsJ2sasHwM1zTOnTJEVRAExwziRHiYUy09CPxBQq8V2x9+HFECPH3OF2lcsqHfwLF8BcuxMwg
ZVPUuMhjKLsyEMGBSPGkXYhhNo46aW+c5rTwW7e2yl+bT45rLnRHn4oTn4cdKiZ+1OSDRfzrAZsw
IVEd2w3yuNscgLMzqmltJi/3e9oEYrtF7c4wXnP0vTyXmY3ctljmkY2bUWK/4+eYaf6AdMf1lCU8
t7Cexqlyg21FZCCf/KRKk2qe7PexlvYZRlIhY0Ytx6oXtUlwjXG3SNhaFbbGeEgwKSBlYHIJRoSo
S9RqZCK2+CtQ+WCmp8NgzVLWniB72iqWZgTnasLZL9Ymyri4VVEeeAEkIV6JbTLfFVISwvIkVrzd
ByRWpBt1G9VR0yr+SxmjMpkHxAF50rRwGH2dHP0/8vqUIJI6eQhzKILuiQX4IASnDIXzuE1HHvXI
ORiP6no/1/vrTfmKNY0jMePjksS+cad6VoY2CDRRUbBgN5CLHkTif8sND5XRyfIGt6qdV15ahz6f
H87nuyErDyScBrAN6vN4/z4WgssFdY5oOcABUa9vb/1Y9l0MoBL0gnid/6YEGAogIJheZgBE7hla
0+ybotudW2IeqW1HqlYQ50+qxFWWdc5l3MQ7dm3Z6gIkpJeQPRMsIgOgoB8dRKDRvSVLMeLl3WOH
bc32O9fk1Zdpp+YX+5eaiti+Cn0LZl2OH9Q2MkIrCa2wcB7HtX78476SFoPSRYX+BPQE5MZrEf3Y
xxowgsBbf0D9S/DLKbYPnJ60Y/Mf7+DFUnXTrInDmCeAyOkfu7hITDUD+uyzu6uvjqfmN3Icr+JD
S+sE2t0bppU0avXdW0Sf3PXj0P4Ho3y+N/7ivUa2+i2rn2IDMz375TmHVDczUJ4Cr9wngH6JEZs/
TXkZ2FzpH2pnosS3vj4vVjdUZlIWqNQVBqmhB+ro6K02K8s67J5YQrJeGmIpud6krW6dD1lLKxkv
jGtT6a/7vRmiLK60McN8GL9KuWQ5iQ8RiZyTdrxokNhsGKoLWbARYiFr1Uoz3lDww3uHHhmtF+/F
7aUv5Wtj4LajlzlJwR1pSGmjNNRmGD+DYGmXJdb1eAkxEntbBAPLKoCAp+M0jwqdCo3+CdDEDx7m
hWg1WqaKHmQkr/BYjVdxL3Xr2bbZqte4ZdHcl8J6nqDtRcJeNjlCeRgcXb6oF/cstdgUvrEfHnd0
6KhEcI6d7bbMN9EvylimvTxuhxBCgrv+j9HHphXtB06Ozl5qzMH50EJ4ER1nKGQn+GsMdpxeHD8b
Ied5p6rz1uGCDZyAYkMwwUvDTyzEwqTkeAJtPZs7EqDfAwcN9e6v4iW/w2+B2jQv1BeZY9/E7FG1
baqw1xLdQqaLDgEKqLcY4AM/B+fuoQVg3yVf4wd4omD1Pm/c+VFE9A1Fxnbr2jJdRwQ0LFG/vtyA
RSKpcM4o+bOnzW4GxBnDUYdCiTJIZ3tsjbbD4Q3fnFQ1c+K7On7N5GCdrUw3b9XaRFK5YlNIJj0B
EqaXKaWawAX7Svb485T0k0a1oDzB/sAX+/aptbcFZMoz/m2qOkJSd5iI8/LbP6JMu62FKedsbMrr
dtkKhYTDl4BfSpPy0ELXv5/ZywmLhKIJGk5zItdTPFXyptGDh9UXGDTT/dThANFlaiI8eQmKM2Xl
wOPqQ8eRWr7vRXb0glr8b3TKUuoSFWQn4uHAWPxPH2FPArUaLRDTpNrzfJDppcm6fKCfRno/MNuz
dEBIIwgVWWlHxTf5JoIlB9LcQV0VTPX77Eeu2WpyF8QgBDfV3S4nMJ48vQfFY6g80ABuSZi6feD/
HFOhv8hDgspS54b/3q88tTaGJTsUMFzL5mBb/WS4hcTvc4ZYV90ZwlsSSqz3KWN5ps5N9vr+Q86F
L25HS+wnA5SEtdLmCXrX2lY29lKWgPcEYrlnDozgMiurVY8dx5osvdqNjISc6M8ZnA1x+gGJsPIj
a0BlU9+3KrA0TVywgIcYGVZGfD6VGB5ZvoG69w0r/IhLnuqGRRIgbvRULlWC3YxeUmRhhpsr5QgY
Y1R6ElxEodxZEopFPd+UNRh3itg0hFEELqOO977Ch+3jKHTbqjqhYsJIWiVPIuBSZshvm47z+2u1
eSDaNHhbRzfAfybnEcH9V+C4UHzD3FR8WrtNNkAeCKnK/XH3f1dx19JC4GFfPNG+1Pwy6siGCQ4i
VwSY1E3IACJ56DEyN02sgiyt5K0Ch8Nkbe3ope4GZLeQDX1rOI/MPJw43IlTC5h2RTQt01cYlcxz
pGSeMqoOd5o1NA+wlbxqhmKuMTbdlV5AqxbFEot8IsxMuk4OlUSPvQ+wLyA5snwOvtVdc6+fDRJV
BLtl7qoiYcToCEXTDbXVQ47ierZDcTN/iw+nfY+eNA5Qkr8SHrPt/zoRRV+FPo8hHTnMlG6EpfvO
oPDbKGXPupeJYErvC9tJU6ZI/uaHB81Cop1XmyDqXcBM1nkXs0c0yoiAzLFdDjWIG9USFxmhUh5w
tZ/ijiHPNc+d7pxCF52TzjY7d1Ub3dux9FS0RGEQkumbqcSewLXCPEvIEkl0tXyPgf9e0L4Fb2Tp
hmvlJbP0yT3T1r28itKpy4NXclHGvSiqNDRqTjSmimx/DrNMih+B6YoUUADdIZTyfJ7jhPNSKgoB
o0K8HT5RcnXd5dtigYZpnoR4wriCB9oQlPy39x/IJMQWNbrZ8ClwEl5/IMgkIwNxPiTNPg2YqqnL
4/3/aoNhAL02H+ploSCtW76/0OOZRvFfCmCqiGi0KNLfG0eCBgNjWLRxpQXIIumYU5swkBkPpfEJ
A8TD+7d6dencKk3p8fbak9MnT1P7ZCoUn/VO9lU0j2m7H+x+bCkXYKzqYWfcKYFT8UBx4nZAEls+
YacZOAKlN7DVK/wbLrqaQnXi+upem5XFYmLIQRbVR5njLAoUzitCnijf/nUo0dj6fe3XTrNQJav9
yIZEtXi0smOoZenrdJeaUxnGQJ2gMwsRzOtskl/Sbyb9ihfAvcr9LwUK50HFVP1VDKQ3LpkcFZ6z
AaV+JHhKFZGy3m3zX6aTGgCHqDVEC44UeF1RJpn327Tu0NRf372mIr7RLpuL8MpyK6cbHX/HafVb
mvU8K1lJusx7SgoycmMS7znEBdWvvZc110qm4GtqAseAK30OJJI7tkXpskWTOkVj7OS31rYZ2K1Z
QW7zHRCBPAA2GVWKbH0FnGLZg1xIXtx0vqFRx5BEE6kMpxXlwRBZeiYuLQu8knyas8/ypgWs3MnM
nOn98xySWkjGTeKfNBZjhU1y/zdxIg8PWLKW6oDcwfqtN/BUFqGlFi/x/0B+05f58UTFuVb3S4lI
Bya4za0oOEwGKRtOa6RHkjVe+py09jQPU1qUh/nxpjbdxzRuIIYobVuDgWhvgVxmEe+H9ao45QS0
cgRA7Awkg4NQgczYEQKG29c1skm5Y5OqQIDRJgnDpzm9IeUcUUPLKoL16l3bYvKYBOJ3b1tHVhoU
C7bvh4sAEQlfz21oA93m+grRcfPoAN8T2plyUoLCdEItoFLgKeXA/JY70JbUQu0qmWM1tt8YFCZw
VHTcUmAOKizE5CS6iNqjBJz7rh0ek5sSwc9gnXDe59rcOPgw9HiAZE84l3fcGBoRghZx3s5bxLny
6x8y0m1Eo0P7J9ILD7vrIxiwneOI3NX0gIYnhCANy1uy0LNTUIJkN5ZgosvdWIPoYCxFJ3CitDSZ
CohzezkOB2BiZhAe9mCPVb7g8uHnvi30qxEPZvSBGb4du3cmW8GtO8rgwfKKO2aoLD+nYBk9LKtl
075h2AdASgXaNpouPQP+tivO8I/CaYdMburkCR10wVs+o5YTqOZVMFDFSFg75Vn2Z4+Eq8PJoona
g9nivlF3FKXK6y6oStZ6ino4AXkOHRPtO3+y9veD77+9sMvGc2RZUdPufZVlJBmEb/qTpxGsJNvY
wYRKZWZvXFE0xzG+aU7uynEIvlRQcXEz/MSGCJDPxOCSotoi1vFv16P7wFlITdRtMCpCCyleCQvN
XHLnyhpyWMnZFv7sezs4GsHf/wM8/phd/XvfI0uKCpyf6IAGE0px3kmiHtntap529acgglrKbgRR
aP16qVTn4lp3cLIotokNNGsXtt6tgRYu6oYry5pZw7dCzDc2Wz1uYPmKfDl1IRTGNvwTYyV9/cEu
bm0sdYGGDSHsI3Ebi7E63hT08JCzxKh3nm6Pgs49ezrxF/4oGCMFMEbrtQ5asZHmdvVbMfoxXAlm
F/dkp3/mBaSHI0LuF5SFtSiP9GGUwKXr3Qp7XguFtynIkGMH/1e7XGZ0MCyzmXQuG5S/U9loQLxQ
qCSlrACiazzKL4dWyicJyLfo7ShkAy5b8HIgB6KJ0ldJNJ15OWl6gdoCcxaJFX+Q2wpiFcqWazP4
EyQrY6g30+UkwyFamqHfBkZ4/JQxXBeS6nY8+peEjbEMRNwp+wJsllmJNnEkJrBGuzCtnp3xAoHt
lIGMspfXbvKuXw03PF7fUQWul7WE1N7OaKrywY9t35Leny0IuVNKPfzC9egBrmsT0nMn6IrHefZd
CFvK+gNJRkbwV2/DXdueRmqHG9iStU9f8px1Zye0Owl/TXly5FiHfPGKrFDNlGS3NNo7+iMChn5Y
GVaND8F9GTmt5xxsKhvuRDLeo6fENMSaqjLyD10spaDlXKEqixBgoUiDnRQYMH/f7eap6OFRHNBY
MIsM34T+eGsWYKroAMFtjU/Cug1GZdWR/vW1E/lQ4FKI0ycG/TCyyRF/OWAEeWJ07LoN7Ojm33O0
CzS25VuslxQECAynEyitFQQOixmxveblbWx/Y7fqNwkkI/6QsKYnJSP33tq0p3dNIrysSC4N0rrQ
b/kIL80KKsVKMuQpigd2eKJmOZX6Kc1N6L9rnt69BMHag3DIilWx/lQnv3H+FhPjJFQo2liCqW1X
/UIvGIuUXzBZEfcmjMj9Vse4AAb9QHmpw9pdQp0eJgU9RILUJPGi/uJ49puvusgm0H+oE8o2mkBk
VaHfR/MhiZlbJQS0kOITwsMqrYm1o2LfMeWN0AMK0SIRovZQsLHwMXm31q0DaAMpR/GWGI4ltBum
58TI7LCXYSW5kuKBv6tVuC73HRhNPzCqsokvLYfhwNfiE8w0uPITOUd/Tz70yNeBzbXSlbb7P7da
GjWGJATkgRz96Ll71pEPTaeiJXY8HumdOEzQ05zAIiqHTvp7Q5oCO+xBCwMYtgumLkad/O9jbyns
hjSOuIUTYWO941O+FiuuuYWBYQmublWXKplIlkaqf1yMyx+7WS2Vp6Krroo4OETumZY67TY/Naz4
zawDYwziaaXEyuCQ5JIRV9OEzZ8vmrivTGFP+iOi3Vp4arTJXR7hLbi77yJkTiOlrwX/aiBkw1OP
hzmxrnDeyZ0HGxXI6SIVw0SU8b/5PRxcDsCFYH8nShVllKXyzJXYqsMo5pnSB0CaJfenHY5q2T3x
roISDhpb9hpX0Xmvv8vD6Ml/0DDhoiyuzMXUd8y2sZLpopmOiFBE0Qp5VYjOD1uyVDL7JuMt2nBT
x0YuhQ+RL5QLy2o0DFZF0zmG2U4TB1X4RCq5fquBfcB833j1+Nqg8YxQhpAcMucRKizQPDJZQAPn
xRzAEp+eaFn4nOwW/B6s59xlWj+za9PnAcPrjtAKvNfYunvaGnVCXnhrnQexy4/47i7XqIRh5Q8T
CIPEQNuQkUxKRGgvbcW62ttH5eGUkQHYP/FwiW+MciVXKW479hN67trGVVht6soqnljhIsGgKR1S
VrwOdCN3pJKCvsKty3JgpAx759HxNkJ+nWI8sk7MZ0ReDqkg87wZDz7MjRxXFbGkaLGLVVCO9o3n
UAWEOBHO8iyKKOS0vvRTOAiEgvLAfLgfRQDASivSiTyMhPoObj46cVA7ncBqmOG4EBKz+VZ4hth1
BjNadriWnnAIlUWtZ2Ovw4l2fK09fCBjC6WQdXcIdeM8JEXgsMiu0XWlXKYHyJqpMYUN9M/JSBij
NmoniZhij5OZ39NHuHLkRGEpLQOh6dRsRJCtO3uOjPPaL7l+BPMFgJCZAPAapFEluUhWnNYmqZyb
4hVSjAJRDAvmohmwBfKpE5Zt4Nb2K5FpSTnDcgf150m4rtW9dC5cXT4RdS8FZ36qUc3pyhIMh1ZV
yhIXqG0GoPtQEvXb4OqlIbvzKuuIi4uWWB/klv311yZz38GOnzeQT6Qele8Si3advfTGmZnjlesr
b8HVUkl3Nwz59+/z2F9ZBJ723sMjvxhbXyIXVRYRrQ2XFSkyhwWrvCvsCGQMbco7LdfdTuV3vQOA
gyp419HArO/qY7Dyv2Sck0TrTXcCjh+Cf387QcvDbSPiCilYYtTq9xgZe+RKqC8pNtu046K7jfdC
lMl4dizk/XM6VWsQRmSsmfLy2njSX11wYNlv7GvsLOglzd8giMjd1JgJ3T6FdFYzADDSW2Hp1v0z
QEC3GPIe+TMkE09XEy9w06CaSJxzIJAy3AoCN/yRUXM1G3rFutmqj+4QYWHPUtmbUYMgTVIckzDc
1U0SCJl9953pNqiAyjrlJs6rPKwCGmnHCqOzu5xOAHqmNZhluSA23G71BcFot31tosxZCfK4ip+n
S73ipZDKIN0AXsSTL5TTF9q2yExEbArSXpZfyef+OorsSzYQt0KHNFYqelsCzdCazhlSvj2jqkhO
jBg2hVD5XOy/EGdgjN87frxYEgUjmg6H4v+XMv1bd6Rys72yvXqZEZOAXspx6Oad9lK/JEbH60HQ
oZ97rMnZWbRN5Rj8S9Q3XLJwktQMs/1cGt73PYRUPXqUH345BPjlKDQckfxOfiuv+A3Zz2vJOWDc
oqYfgkGA7zEA255OMaFvPxRioJkxvUMvB4SbkJuRzrG+M1OL9nRAj1pBIUBLaVFFJvnp1OxWvMNI
OZqlVBOHg33SPnVnGU/qS62JhUp4K4Da+5cJg+FwSb/FPEpHEQeGDmZBrnria8yMkL9AurixabYx
20GXtSQoUJxLyeLO7HD4k87/Fi3YkYYijrCuqPMlilOmZumh4u9UnJ0VCJ4B4y0pirD3KXYIL+HC
IomJQ1N36wG642MBLiLaUshJCXAcaM/yaqxZ5k+lmAlcEku3GvT+cA1SaS7D/PQeMmhI4He1QarN
uHcny/x+IpAFhFEsFcRJHGkRKcaINONSxGIGxN+d9qhgPTd0xU+Dul9TYKay1x3Q2C8wlr6XcpRi
pn6Ka9FERP2UzUsTV1IhMVo3Cr0/x4yY8N6KlCma6PHxfdW/ys7Int/TWXJVap4Ry4lNR0MoOQgz
t3Z8E1efe4nuWUfseyapEylCMZuKYu2FQ1GoH2M+/rD9qdUurdhLX5n+C+kL3ALOZOIieeL7kMvS
JcFzWhYTiw8pgJIsx/3h3HrszQC0tgnWeGFWx4ejK539W5PvRXsyH+dot3QcbL/A5ceQkgN+ZV6R
xeD9QRPXerf+8YqOnWwOtOhqelBXahUWTbCwQeU1JsNl56yeVPrPoALNr6y9HJkZwBpIyspuRLDJ
0l8IqH0qTVDYskIeIXZeNMqKSxOe8vhJm6kxDNtdyt3q2g5F2SpFttjkJIJu2jG+A0k6jxZ7HJ/2
PjvX06rKWr00sWrFpM+vtm1Eg/HAn2l52Mp8eHJJBia7pPSvL/dmrM6wfi/mw8ScLksLOpTcj/q2
F8dFQEeVsCg6+TDPpmihDvQff7DJ47Hi2fVmd8M+f0vxT3wOYaWv7dgo33TJpMvHiG9ucxsoEdU6
U3f/llv27l7FBL8vWDicScscgL0D/99ItrQ0LU1Xd6v3Dgxx8TB8CkgR3IP7Tv4SVHkbzc7HPNCd
QANXZYJkdRyRYvldJFC4XRTcePRM7f61kGt7hYp6yE8jgdbqzOxVeaUwSykZG+vmImp0U61PjwIX
mKLbQpowfGH9O9pKQFEFQ4kuMalv7d4tHvtaETSGcB2O5AG/MkxIs5zbJ3wvUMRBzId2bh3/o9qK
dHv9hU6yrURowAMTkiTyTPVjPEEE/tnLEfg/30Jlk6uIxHMVzQFefm4kDue4kqQayHlTKLM10zAo
CfDQbO0Y2RGt0zjVJwq5IZ6b95VSfvqliggA8PMrfPRsZa8V4TK32LduOcc/4hfJ5ccGT6aJAOu9
8nSgYEDL9YXbrh2TKrYWSWcrgxPjlZ1ySk/qSNCxXbqOZcTB5U1Nzpm86P4y/hSfDpb1+FsWNoa1
XvoPs6ew7QlwLLuWqBtXQlPlSXyMIP/LqAwsDVV1c7fhh3gjhLkSd+4QxaMEalvHYRXB2T7GbQgT
nKzseTzBE0r7JYHNUUmUnQ+0hgexpGHDYoCjfDId5yA7mFFH53xPqth40hn16FKUQhzsux98Cc74
JXigjOo9lwuElJIFgHkiKB/4J4rFcxrQI6fu6/Li37Azbbqbj7i15ev2jdJ9SYfKfSDStn5uJg/V
q2nJ+xs7KiietBQamRjUd3Y49usBhqs7qfDJ2mA1mQBYT+hjKr18FNLQqLMoz5uJUj6/C43vMfl/
jSzgiS1gj9BBUyVL0Z1q8xyTe3JLN9QoVAVHNnEV8wCIf6jXh/nmTr+8CZCxjfMVUIKrF1MCa6y6
aAtLMbX2ZzG2FwQHhJDakJpFv4Yq2p8wad0PyfGl5LWxnkJhYGemi6vgJlm4xIGrzfJ3yq3sgTek
1IAiUmhxK1rAKW4PSIvijJ+mNU4TuifzTc3qzG53ssnlw8cMuG/HsYEXj4c1/PTR01JhOHrKKGOs
NwwnEMxaqVMrea3+/O0I06kmi9ECsNmS/RjRySsyECjWuN0jKC5EwUnMZP+XD69Tzhqr6pp39RBv
mRi3AhYZCQRiBNLE46kwPZ1UFMrv8hgJsX6XmUoHq8vS/Y9pKz+WLkR+EZcZow0J0zmDRb0SWiZJ
q6spOSBQzFZTRlAc7+vaKc4tNkHX4z6nYsP0eWr/Gv9SMAKkn0EW+AGFQVDg68FELWncqeo5QMTE
uXrt6rPhNxJApK4A7kgmkChaX+t/iWWhUYDIzf1wcZUeX/9nf1DIQy43ROl2LUIqdUAkM8uH9CBl
fOl+QdGsIk818G6b97Z4xTpk6d8veGR5LKvgFv2uIz4R6jRxFfYHFe/7oOboslu0Lit7M51StyLt
TXMQquIrX3HVMbtXWHWAPERSOfCklmpC4HLYExlBJ0Oni5mowDh94iNZ5pwxWOv4OPTtKeAxEtQF
HUYlhJNct3XIPo3HB3lLAtSDrn+Xa48V6a6TJWmP3InC7vH8pJiixfLhbsOLsEwF5gZgiIR2TuKz
t/ikFrsYt2tP/8YLL9IsSPOBDxoXwOEzbX5a/VAvuinfiMGTzWkQUtllImxsMRLU7WipReheHl7b
VxIfp3/dKY+mkDFB4AwbjRLQeI1lJo2CYmpQy3J4P1r4gI4l6B9Uy220HW5mcZ3S1qclGScuhDw8
QWmzNhrEa8hgbb0vFof5jv0xtRenpz4YyLJx3Jf2r5ZR9YyyfAG/bqniMvpmJKQs+L5YSzzMV+GP
7PzzzZMB46ZUSQGWpEl6rJOAvg/uxV7FY+CW5tKpMPX5vs4M2v0OsSi51vnJAd5974a+UPsL1H9X
wkDSf5P2iurdcFhRaIPO7gJ63HLY5YSeO/0C/+MOwS5av+wT6rDUtKKTYS5K8YviJsAoxkRc1AUK
n6vD064jQ5UTfZl3apGxbAG6x6kGeQbmsUzbi7MThm7P376p/eZabKjSfuDGMMJO3DHvYtdrYIjg
V/KHL2i+SonIkQ5GBQBM/4ssZOiY+1mwdLhW4f6xQ2fww+Z6BFccyYDKJeE64r+NybXUUPawTrYh
I0Rr/SjvHxiqKqGYpxUz4ocTpUO+9vSgnsF2TNh+4o59Q09mLvQx9IDJyHN6GbGk5HRFfBe2cP+8
8vWItwX4tsciFZD5DMGsMFwoBu/IWkERB4TJ6KMdFFOp3Kz6H8tguXq41ms48KzkYJa65dZPzLpE
f8nWbTbRvVyWQ/U4P8yks8NDy37c8qLhMPok/wyEu1x2/8b0e/CyaCNORHMzpRFfjyOoSD5m6dal
11RP/FF75vTSVSRrMX1GM54fCCCAeiMNkXQXwL+xo6VU/SmaxaKerNt2ihiUfBdUmO72NH3K8xFK
BZlFVggvtvQfvjGk2w1Lop0tLWPWSjKUAH/QNo7PnQQJWw7WdYBbTVDeKjgHa45g4k1u6yTnmA+2
CWjmhRZusyunxLEamCrT/Z37QScMXSnOq+B0+8By/llvRoOb61nMzJYhZdAPELuGc9riVnvuesCJ
LJhhC4mkVOwFxZ5UWJ553rGyEQ+CR/J+BDjxRauJ9fkyC+OzrWmDpIomIDuciZEIm3XB5MaAySvv
F7FgUkg21lXODQUWgkm5K4jHpkW8vBEQc+POPzl7a6CoXSIc5iWHTHw3DtFjzylJERLBdNwlon3u
SKgL8OdmBcIKKQGU/lsXb5++9prdIRIE/skeqZrfTVyqE3nEMXUQRdXPYlR5hmjybgbCnWsYRFED
sUDJcEPJyV9gtzMeM1afVC/VWtjwRC1JyacOd+MJl3RvjttwF2Fu4LA5VzPpIlmTLicRLqDnxVkM
boTH8c2LAsGkHMH020UUl6yG2iBv0+4Z/sqYDoUYQ0VpmAJkYOMqS8pt1begYFjRwkbOBhbYsdWY
arXhoKr4JY5e0eDWeESlbwL2RXz7AasPvlqd4akUpYrBgEeNThCHkAIvEIOkq/UYiBsmb09myMdp
lkYa2tzF1369lPOPfB/4+Ny1Xi1+ISg3R83S1Xb5X5XeWKRsR8BukUClA7c5xoQ/n0TVYKft9J9l
Pb6vpXNUEiFT3mZ2YMRziLVEJ3KV9oXGGnM6pqy2i+S3RA/Kbj6me1k8/WXUI6W7HTCCEmGK7SDz
ZrSvsXSwni8pIWj/o6ebxEeflfcamuUx3bYyFIZojiHVrAi9ECh4XWG2IRZkuHGRLg87JBImRmkt
SkXEqfbubngd3OL053288b5zeIaNFoUdDGnAb1F6xqN1n1W8kf+oht8HPBoThk47LORltrh96dr1
1NK5JM2TAQspwF2gFnKfEbBEPktEygg6vLUNSyloB91aLcBJCjqjx+vHZAcy7DyA4b9YU1sUtijM
TT0Jlre9xa7LBtZoAkGOXkzJVR5SLigruha9fM8y/PUU+WCrfu3LYobN01Ik8E6P0T/wBOQxKE1H
U3vSGYJh5WjA+0YrKQnK6z/A1qI3TI0xlWW+UrLIyp61mnrbwRt6Wc3uf1eNdt+C8XLIM4zkMsUI
vDC7L/wmFu0h66QDlqdqV7yvoYoXVBd4uMR3YrEh7WUHa7mf/p2iN55kRLHPYpQIdluQInjsHZ6P
lBf73SqpMgvQqbifcq92BMncUB5ZX18SVJbFNHmeUQpnD4ZwKpOMYvCsta33+BYDEV9ZmQb3cgoo
9kf6HkocC7NQ0esgVBDiHgwKiUf3jY68yElwz1LulY+xb9sy2bGTqD/TocoDQX/ntfVbZWobQg8D
JYOEhbEs5EqDnNbJ/wPST16vFRysZqWyXyqfh9PzHHbeav0kD5zPijtU0Sc3b0jRVvsOvZyt/MKz
+wKVeldpO8zg22D6pjL82Y2q5QjnlOS6wzAVjjWyDUnVpIlS2hCjoBV+AssknbdjFgMatU9m3znz
yB96Jxi1vUOOZ4SaYo8zZvwEJj55pgmkYphLJ4KUxjeadAaPkW+AEOofjLvnuj/Zf/qlWQznpuh9
3ozZ9rOP55KG/qTXvsDviJtDjZ2kfV5vIuuEwo9hwxEqr5Q1jGCm3MiZZawpr7yUagOqFO+ZYRnv
70psQ5Kdk1zsXWw34HbFivk3OUT6Tj9kHMqOmhXfSrvkIocVFcFMm6EXH1liXqZV86acwPWQ3/ep
E8gwkfXce+2pg/Nxe8SXI277y9Ffrl+KTtoHKOMcTKXOKCLhOBf50lO7PdBqWAJ6woRi6OGGkiAh
lFOdS2eSgZZ501lAVPWM548uyLguTkQfF63HJJooTpwJ4SO+YWbCdXVLoOf39ua1CDYWRlCea19n
5EonxOCHfhnoA4cCVyhyEtWOLqqIMzxs1wDWGvJwSt+NDmFU8X/2gJcEDqe8fPrrsodKJBIw4Y2m
Q4uKoO9FMY+3PMV1W3sz0uHC3luVAPpJMIaCcH7fk+4WwlzrOl7tlxf2bYL8LGLJN8aWPl/duWU7
ZOgu6s2r63QtomLrMGl5kz5OpxtKTb2EivHJSAEzIpPDmpgy8pOUGyMrO3sYus+atj/9hahcFNhU
g6/GlYPOKXyzKaJY/vHJMIG5Pls5e8AKoYuj9ObeLZkcdcHvpBkFn0d6XELNwijPvx9B7ntpIo+U
QtaXFF6Fb8/95arLpnkTD8YCDuJuVDuw5vXZFaY+DwWHt9qV/R9fQRG/Fxp7cG+XNzRKPkyACAX0
jWiusNMfy1ouwtIpAMyTEi78cWAXPtsS3w36tYNQEyQyLjicjwQGMIu6CWrzVljQTiMFOhAv/a0n
SGOiVHle/hRGfse0SuoRnVZgR4BKFwCC2qcEwyaZ5lWibl8xaEGsmR3BNNyyHEwYM3XRpG2XtDdF
knTdoYG8aIgB/93u2dkosC3SuPec1PXCT7ax/OrGQKO3SGcFSuD/Q1iMG7wvlTrT5qNpCUwRyjBm
W0Tkvsb8p4XgqdiX7cqXl017r3aJnJph3VACqJYFJJiZmBiQH5/g4F0ZqA9wyZaEdRBjBgygqH7L
C4cZO9uGVRPgGjHW6Qs918nvtGttqNJPy0kSBRyaOlLZEbTlkIHZqBT1gLcHbFj69ky2afNfcTAu
l+TE6y9rKcKGMvD4Vyt0qEh1d8IcvxAea56paKYsyk0UULeInoprTmWdS/uMHNUZAub2BX1CU12f
fI6PF18aXo8KZU8Je+wU3JuuwAQz0tZOK3rd9dIf/iGyJkPBvqTcXVnN4N14UT531UVOOECRc576
pbgoL0EymtQiWp7xhdSaRsLWXDSL59j/dIxIuTzemlMrtoRWWSVDojmtTbSU/IAO3KkpTkyZDlAi
dgv8TfuFQC/Y1gXxlZKZXLCDo72fqXN4SF1+mAjMg9A9cwCp4zBuAyuIXBUlmQHxEXzbHebB2yDr
pfeeByal7msAq8IP/2tEitsxVr4hnAgWgkm8XlM0R2TlTpbTSa4rsbnhl24P0mXOjMLAsKOwwANe
TjWc8pAlcJThoXTDC2Bg0e9YMqqYTUCI+9LYai7ajRg6nE2/MFzygi2drWMfLrTkz14VlcvJBWue
W/FZbAZYEMUvWqhllEYeVN7BtG8QsdXP/TrGxbwwejO8tUJH5wMR1HtrW+wmDQB9rz52FHxa7JRs
GzHiaqhUavN6IT25b2zRb7u8pXb1OYkjPEf27DCTT5SqGmm0FKAHFOYFJtmXxao9EQUyAF1kzECZ
RcPJ/t1vqf90Q6+cYgr/jQYWFxoufUpwyh4dEOH73sKbUDLcUixxum1cPViZsvbOc2uCUrG4pLf3
Fxs/BiZu5MxuUV0N/CjJJF3hoivSb73ZTDE9SaquRoTRxzHrs/yBoCneZ2nYXaJz5Llukkp19pas
dx/pZx8Desz8sNH3gr45tKJNNx7S/sa3wRQskBHvgQ/gLyega7cBHFuJmM4J5s5hyuZ5auyIZfuA
HVok3SVEppoFp5+uPxPMbhmfndbClwPNzGaa6gplR3iTIEASj0IJNeKuWeQnwo83tYxoC+ZH7q0e
7dL1T44FK395PCkL2tfpIr+FNaggI6A44aoa2APlgapTFvOdiJ/+uFDaqpZTnP5QvCTToBiUQz5h
TzBWhzssTooT/Q0dQ9CfVFssp3z0PFKNOR9KsEexUdwdP8HllJU90W+nRFPB+qBUDkPIgRVz3fTr
LudqTvEVUObt8094PLvI0aaym8YknnIrens7xu8n9fYOlXDgnLb7EkPFYa26QRzdUqSqZr2FzRGn
XWlQBFaZ1XfDGpO3a+vpBj8Yna/5GxAudD/Swpy9hyaauA0l60EhNjVbgTyT8sTMFZLbnLE7JMa1
cjmZTZYe2V4zS7Qk20HUUjlunJACXDvIyHdyk4aIpI7uUGd9Vwuk/gOwtk5zOuxCpMzJe5NNxHo8
JdYXx49y70rJviZLhy8lujKKZrKUYQZHA9nXiXuMsS4LCPo5tBBlYG6+1KeK1UyxQ7HxaKUMEAeB
FzSSkfxQLdSuIYghXFdMFuilg0zU8P+kxKnZzmCiE4koLe6GqL6fA+WJpzib37AgUhViZqWJPm43
CrLbZumqWvy5T2LaMYz3wpUFwlDtQTHVn5b4162JShwMOHywHZw4qrIlyc43T594NxJmhOF4B376
tFoOF5VfQaorTDQPPVEgkwBOMp9FiiRTmu/yukqceWbo5lisouXaOVJCqkRCt3B9u9q12Ns8zJB7
OFVQQszK//+MKQx+NileOTifTwN6HH7lAoJfDp2ONVtZX2vshS6DVZwnCb0uFySMoRYEnjSKkzEf
A5gbLx5+KfXvyLx3/McXrSqszcXV4hsY8tJn8PG0f3we/OOOCjd/Bt5WaZ4Vt+GXb1BIlvZbqfQB
7CapYpFQGgnT0bsrQkl1v3Ha/4AOHu6xPoJd8eHP7u3VIz5u741HDMqfk/F7a2PwReigi1Dwbh4q
UyAmg/o036GZCrxGGWECI1oAJ8ZvIzIQ6WCNlrT2imPQ9zrrJH39gb9c6GzDSdReQgu4kGPruue+
63AHu+exvGv1d3HEYmgyLDmJoIeX+/TNDJnpvGka/hzNVAS1RAUSMqYWUX14Xr8caUbWLw+0mDvl
i3j+vwk35CWfWQrhz9cP4MR7L5n7vgQwL4N5NEdqHzkcLt+RBLQfFhKgFvEQ4spJMI/6UolqjHzb
BSRzeR4zN6xQD9qR3GCTtuFd9G9/kiiLoRQUy2tOeOqju6A83P4KTYSKhFJTRM7LrgwvHELB3STF
f02ZE/kjWirKcrqVZxcN5aYEp/4epfYye6IhA+auTQhOKqUg+ZNG8C02W16sWZHD2v7eFLJZb9RC
8iFNqRmXHCBV1FdYKn9sAT6MFigQsxRU/aoknix524mMixr5zuyUSwJ9LJ1WlToitZkuhxxx90k3
zxppDeYeC4KB9qhkHO0cxqU6eeGGMlLBxGipZM+I36+QA+uTj8O63eS9VqONo51tOkKIjrm5cP8k
/Ea03hdDfn50RloqKrkhUNryzckRZ0K6tD/166ucCNg0Nd7ilvhFkpLW9WjDDCVOFyNzJ8n+4hJ+
FYHwpe6/PI6iAbI3JFSHZw+tmw8my2OYkIej+Lul8HUP337AiJZgFg4xIpZT1BEEVDy7dlmfIlZi
sx+lV94cxS6BvlVzfYnI4Vfb+Gu8RD2O3KX/h6fwcrQqr/nskY7dTdo1CYotrf64WNSJpmARrkCt
AbLNxPzqOTIeF6dfsBrngDkN0V1jrc0LzrDRhGskNEZLBgmw5iw7bfFSWEXpDJe3rCfEYLp+iA5H
goTtoAJTOkVYAZLjCFHkA7niwicVCuSBo+cbJlnJr+DrPgnoUaI44rFm7YcQ2AskHF9PfzYfCrRN
sajjBirWn5Diy/9ZetsXeMXpkT//EwaShrKXd2vO1pgo3r9FKM6I7o2snrySxx1GJxTVSBfHHPgb
8ZeSi5Mfc9ISGk0uyT++YQuj4XgDJzDMhlH4EVa56OHwmHJhqU483q8qu6WR6QK0uEO4eoRdCTGi
f7A09+7hbuNDpDizb2kVYd0gTVj2gdNRxHOTL/rdsHfHL9jE+isJbLYrkorXnwEI+Khl1kmynnjO
m82WPAmo48vW9eZUW+m7uxEVYqBfEtOzTaubxgq153C/dtdOap1I/Kff3QiSYv5bGNLWV//pfmen
B7auYQlqX60R0UKutMuouj6gZobDGskSyypuWq/wMylK8xP76WdgTftZDle9mvSsZ10K44+Gtb52
pKK+8n8/VI9RCagQSJkXh3Ap20cB1r8J23Ocub+AOrT+ZA+EVpAxEgCTGaF7PigDXC0XAV3tdZHp
dng3wp03CuT+jySIUYrKbFkjMVBPn4gYVzKsxZwHulLPI5kh3UtBJBfPu1JmJ6M6JPaDKXbGC/rW
ZGpcZaEapr9KZcb6buofbEwnjdgKQ6xAsFAmQOdVTo7bZxiQHoGYB+J62SjSECtPGEnbGvRFDEPF
kpGRfnkGtJEjIUcV+aeFDPGomCIWGz5Txi7Au+3GPGyBfy9oIVDFuv66Aro1IpCiGPvuKCwwzzaD
HKNg55jeRndYWvu1JqfRuOwu0uwRNErPHmqg5m3vK1ehJssLzT8l2W1cPUBqQtuES4tvM1QyRAk4
bZsEybDSLCoHHwvzGRfuDisg3pyQnKp2J3RnEhJJcdFhaQOzMkM69zBBj7DHE7O1tDvrFPwuqGEv
ltJi4+4BIL/6NN9pck/WtjNwk3NB/WgO6bqEm0wB0gswKXHzLjHx9X7/gq9fh1uK43r/VWw/Yggx
a5KM+6ckxo4wGWsNMBQJjwWFuIdEPV0uEhkpzxEPOB/zVKFQRdCABWxEet7wzEENEdVtX5tom38u
ayoReYMsczN1bbh1Hxz6A6wb+Rgf2m3husqW2+WoGWb4sBo1x/VMpPS395PrJBCdP7agNS9nL5Bn
QN1KnR6piV4joWfjyS536vMXcSgzvx18M4TFTlwrhUWy+b5WRH/6jbaaIVdukPSrqA+8YrM2jocO
S+A4Zih0YKlbAugUfHRERPlgB/mQaiNSMu+haxPlHWEvMIx+1iEm1ShvW1I468WUIGsH59MGusCc
jULULAAamOmwqWqhnfhIal51HlG0G4MtRC4kvaHCXdArOfnbmlVTS+xxc4QHepnOG0qYHBrz25Ca
P5/CGeYr6GWmzdnMKTN0tbrihMCkiPGUwmTiCDvQfwJMKHSjY2cEFZ9uLLqNRMA79Ui7CTtZxu+0
r20o/jKs/NNK2izMXCwB/Mheko64Q8ba85fSy4MFrPyHSe3TDkzilvhRm1Kva3BARXWDfsDwwisc
2RAHIdRieZwIHSQjg6JRdd2n9YBzcTDEBKmU8IrKsCOhky7vu6dAsEPqAQ4XGYrcMccxjRn/UNwR
Vq1MacdTuzvUT3g1LXhDsZgXW+1bFHaj+vLgM+k0M939RqBxNr3AHXHIwdGH4GPrkaQ3nrB89qSb
HwThz3dLiTOrs3dCS1O5X1NMyHLoLMeZES3rXcKDQv3CG5TDTpXTiQ2BrLuyh1aRMSpBTDUm2Y7F
Top07Lar8pKCUrWhZKK2hw2fPf19VvsmJWY+3xUsUueZwWbL+M82mqTyZUmk3C68rEBDNEsM1KyK
yMg5OoabaX7pG51TjCTy/DiY89TDL/xWikRcY4l922LvN2MF97q+4nyXUY7YwUn1G3d4APGxEoLK
SF5dHPAPulhRjz17Nu3BZ1MYQbm8J35w/qlLvNJ2ZD9DF5KvsSaGapW+jqltIn8+I1P9lrRkGr2t
SZnQpDC30GV3ate/sNMfxlxXHLdbo4t8jzkk/d20Xg9fyGAUbbmbTnFr8u1fUaWw2qb+o4SjYdBf
WReBhhmIFLX1cH9++f4UAzcQRxTKRgy0X4Ke1E3uGXRmjuX4OK7OWp4O7oumKJNJfbyC6ZlU4N0Z
1IMjQy1Kl80AGbHb3CWIZUw3KgRp6ok5G0gw/HDPwkUV8C8+bV7CaRRlFwqUMaAyQ+CLej0ZOCdn
lMhr8RC1EzPX2M1s3JJQWZvGc27uMXNF5v8aFqROoOD6JO6fAYh4pTeJnCyyTzf5k6Q1DSJgunU0
+Le1bGGYZlsMRKStndL7sFvrtRuEf+7/aIg11JakVGmgCs3kpDpXvrPL9pHNdanEjzURvP5rPTkZ
tU10iKN96t7Tqy6KwyWRG0f2o0fhDDRYSbR4XccJyUP7qDEwwwCVsqh+euKkfuouCHPTZJxz6tPu
6EcBxMwDHONOsjij+WIDhBZFGqZUGYEpujhCOThuJlz+3/v+ch0W2glHnBT4Le4JO/jYy+2CZ11r
8s5L1kmxDFj76xpeIfdthLwgP7LOh14MLXSZ2rFQyk1WIleTqrGMdE6HaiJ9aEp79zhYeTBOpd9t
0jdhCI445jbMw6CZ24UVCXeV5RUeCVNQFJiuXdIgA0Al3/3YRaPDtuARAqdEC0d9x//9nF9AQq9t
hraBxByvJfNKkaYz5y8jjdsNzeeoTi0QSyPTpoJ42/r/rcupveI9IJ7ccl62frORaWWa7u7iaegP
5IRVSlYKFBiT4NwweDxLumCjmO3qgjDm7c9LEM55qRvY6ay7H+7+F/YKCcgaa5a9dzn5pYwvpTjI
tIpf0019c1FodrDNlwDIURpqliEVxTq9Kl2YnwB9WmJrPI2gVEBan/getH3UyZ77tNZV0g+grz0Y
8S3tjhGXimiM5WOua36X3jiG0v2uV9QxKHSc3vFbbbJkzYOFTIAijtIhDtWzm8XzW4X4q9ucPLbn
wCTK4H4Il/jdF93heDyPxgUQ+6HAhlVOVUL6Lmp/L2v3epKXI2GDM71W6nEvMitBI7gvbhD+ABsz
/n/7jTmag7eKDwu+Z3fKYoRt4/nD/2ArTW2rwwbxSXlwQOpE4++2mkf7YvokuEp8Xxls5Li/+TJi
9rnpOwVHXQrvycBtb6EIojZQtzeANQQjVL6qYpLp/dC2LrTQKeFV8w2ZmP3sdlx5VAkZP24/LtRT
BzeiSSYXfjI7P8ceieJKyC//le1IbzBpTsYtfqQyWUuA4gyJhs8o0Bgp/HlVEvKORt0pvskhZ3ip
1Y5LcXJ62vXd3L60z2G51YSuQUm4cenkyaAQIbWo/fpM56b2W1t73Yr/4nVP6W4qFL57KIbmo1Z7
fhgFV6y7uJzWJlTjCv/aj2X6jmho//O+dLGi3yRITnF/oOmjjv74cgrWLQt3oqQ3Rk9Q9jv0Tqwd
ewUsxtplNu+g8SAcVoGSXKCh1MOTA2fpkcNypkGUUDFUZk6ajOra2HWgQn1x9sVjzMa2QqHB3heC
5/o+04uzsr7SygUWpoiU3t6zecHXGeCkcAGIGqSNHv+4NBmT/xXxCjkWtayQ0yPjFU78MG9WWcD8
Vyih/FYJQtA7WApFOS96gqdfy6fx+KPEw8YpStOY03Hl2v3ldFCyBXZfES3VIO8aKjWOKe+s1BPC
DaWV+MPla506cJuRqdKuoh8yQj6sX89X2unmTslFcI01gXQuEQOE5b3i+koZ0XkZoAGckXkM2xRH
wy3qdQRdyXr+sLUKUHxHK3yd7N8dkG1siLQ+3XpfRSwaWwgw7qDBFgnzrOtDSTNwEt+ifT4a1mg4
2cp4zbIdf4R6029A4Q2LvOlkr6pymUeYwVF0BkVYFUgLpFw5HH4dSuvTwKaZNzmBZ/iB7ukTRK46
oJYodZIRFE6LOPTWvZYhH2SlF00dyg08/oWGM6d6XJz1ey782ooo52g/vuCZjO72oflPq9ewcOSz
EgT55NhwDtQQ05RgEr1gtBmCgSXee8IIiOPB85r65R0Gsoxccje79zO+icBWMEGymhK+NFDdcWDd
iopXCevlGtRj4fqtvAfY7wRyryMuTswxoEj9PiElzuChvSx9xqMAwNMrMFCb7Tj/bKLbeMF4uytv
fNNglEncz1CLe9lEIXqBOFfrcJDTNJCo+Jz2zibPJEEx5R35mXptvIANGb0IDfW2cjJUNcl5PgkD
XHV61Beh1t/f6PGxcKc9gskiiKpDCtjFThq6nnUMxbeXAYTnJCLpHdyX3nRmRqGrbn6gho3mCgVF
QIjV+leEcym6hjiZEhmS/xZ+5TnUCn/5KzUd19LIsAY4KyiYIPp6oEogSOl1mokHqmIA5s+SBJ2k
3yi10vK03R+jVDuXW04NotpbMe+hLwyUfTV3RGF6TPhM0n7VPY/VWb4nfuzCB3Gxa7c9GUdjGcE8
E0YPgiZrw7qCadP/zHRlDgQNKOSVCj7bnXAPJJL6E96b7RWvuH2sBNAAyO8auqkJxNZnMRAfEWla
g8dUPWeQquOSBphrZhGadIOTaWmpUYEmw3TVeTNsQKkUCD8xxckWz18FzY4Jc0KZ2FWK2/ICOM9e
AnGjxlyhglbAEMV5rJLA0fE7+SzCtJHfLnitwKCcIY4DBGzAyXUeRDqp5LXb1XM08yBU0+uu5Zio
+H+ip50044Zs5Ju84kg9hQPLgPv0EH0aI8vH7SdWdBT/2QyrXAhhZfXZuOBIOr0rti70/ByPPIJU
JfigCn/GiB2HnI8N3ZfjuKsREjZJU/qtx+o4sxsoDJuTvAKS4BcHnr2DM98v/VmjRbrImtZCX3YX
/nJCKGZX6bm2fDNrIGy/npoikPPzcz1DByBf8f1PvMqbNc7ftTUIaBSw36090SASbxImO61sCRjC
d/nunePN95IN8c/baJ019qeFn/2epj7EGMNf8FCqkXl8O99jQ6jDCw0gHgC9MsxM/9L9o73KcxsB
gwsMY9lFFcHWYURIJz7F1IOzcVsIfuXEc5+32CWRDEzB44cSBCjAYEyf9Lbkd64wlB+l5vumMlCo
PhuHV3TvOBU/I2exJ6NK6Vast76lF86khwJuxV5TCV3qAzfNsDHdlMpBFJEKpZbk4QfN6qSI3gJo
RfIdqMqSABrsUF9u6hRxTSMH1PZLMG1WI4gXjHHmnUE8qbd6VBDgVoWyh6rXKpkkFEca1ykZ/46t
FEus5ivS8/S2lIwc2i7S1sAxWvsnPoh5zXmJdafSxxwDJ4NBfs/Aan4l7cKQnS1b52h45savntr7
sPb4ykSIrekFE0CRbNXy/+PNdt4HObn2gvO7ouUctTu8CERQZ93zQcXge3kPqx+DvK6cVOsfwAiY
nlKFaaMmNo0V7tN7eP47Za31i7ka2waLR0Zw/IJzaZxNFuBmCdRyp4Dd69YSTzJs9HHdQ+fxvHnG
8328jBmPRbckC7n6llEmGmNRTK9JtgO53/nF6bb8AEammsQtuv6wxEN1ITfiv4/1Nxc86/EWPIGk
TMwOz10znLdXQ6fsJV2IE7nOn+DHyFedjoXE2PtrgLorA63y3O7+anr+2Di+LY0L3d2LObXghPgV
x5tz41J9HjXLGn/PNitxpzf2lIfcVqIsmmsDfS4mhQ3/O/AtEee0kssI6mfTtv4soeDpoMs/bvCP
xOAtY+j1BzHrGaP9i32uWMrs4RKDryaAJe9wajJtAXhJh87OVTZj2TAvFVIdCke1vszVJVSNzzJJ
GIqUUlX8deXKYQtvxzB7JtqAasKuINCqmWrs2P1sCBmiA6MQSnk0usXN+TXfUuANxtHbmPSuFSls
bWPmSEEWuM1uZlNpfMdYx98Fj5FfWd5Mj8iRR3ATSKxWFx/miXLtgmZT3edFKs3kJDJu0YfhacMM
ubA0sQT4nkHrSaeBUCGLE2QkBIvT4KoPoDEcLNDa6sCYWR6WvsHtKmmGWslCn7fdZ2GsD+CWoCdC
klpP+O7EAWT+R8eXjd1ra4+N8MFAv3K0QAyWNu3OYs4dbdFm4mUHRXeV7dK7SQ93RJpMKW7mOabv
j9YJ7d0q/IAxoR1RyevCnRNWeSOF/CRo3uu1oAspyO/sLFyFMbjxEaowS/VoRJ38gkxYxlSOD1uQ
9xENiXxWqW16Wr7leNy/HASZTk8ks2PkDQcIxP3LEzCn2XBFvHrsG9jVlxoq7TF+cocp1rYz9Y1C
Dj4BzdJISoq0tJBjXmmJFLj0biZhR7xWOZCwQu2PfF+ncR0CMwyF98wSA2NqewsjtsltwS51mBPJ
ZkuFogpNRz4po0M+SjgZFFCDv4fE38DohdzjWYj5ZUN5rGhfpgnOwzEwjWF9da9Fo51yXA1ujFmH
whY6rMIC0ycfbk3KAEqLF9sZkrhwMfGjXBKQoTQm97fjEVx1BS/RdMuNNhV4N7GQq3YbjHwkywaD
zYoE2r/xEAggXbQyI6Gbhhy2pCWVPmjxlIwUongcegyyCgecCz+I/A3nlCJGJm9rYoAfr4c31yTs
f550BZbElwx8qXl3JPralRgx7leAOxVgMbUXy16wanx2EHlZQbBphAMPis3WHk2FPAUyY6JAeEKJ
+90d7eA7Tz+IzagdhNmZzIJWUv5WB9A9oknnrigWyrPOuihk9fBMjmivJEcph5GMPXc68hLi0IXv
7OTDrRBWVxS/NUiKU8Uw+AhLTVIQhADgFUh/L/WHWjhyfbl/3IrTR0SosDLIfdDwpcGYRocPLUeO
1KY06d1CglH0WlPjtyy0sCYDQIGLl3esY0RAvBJ55nYukLf2rwRs4kAyhFX8NPgmBddSxCwrPKfH
CLlUXXlwExLZKFyt69bSqGSCg/Ur9JmKh9ODdTQseHrXKPODgPR5LK3gcfR0W8V1nIbfZpKSXaxl
98wyc1DRDIjTBw+jVYmoLJZ9IJwUnScBAli2vJ8AGFEAHUlOp24XzshespAY+jd/ogS5YH/8QPOt
xb0U47vCd8bkejyN6f/Rc/y9Hrn6zKMbvVcB5Gpdmlwe0/hw9uS8dUClwENF2k5liOG8bv+W+fuu
R2Sc5dEwYAt+5LqaZiYIharDBM7Eednj7eHfPE+d8cis/tZKwSM2V53L2rnUJ7fmZvkDNkrq9uOx
eNP3nW1+5Oc+Q9vLhpWZ4ei6SdhjtikhkJYMM9Ee4sQLfAVBD8EQ1hWqttVLJBkymXrX92/dslAq
nXJulnDLBY3xp7BdMnr7bg6BHZ036I/2gSKuEFUs471egNDmvL/Jz23nJJnZvQwb37vsZWIpA9xE
850qjejQBky0OlL0e9e+jCD9DmF2jePcLHOpmTeyISzTrwu/tOTmytryiBgqSOxo7uFRbj1hMIGZ
IDd7HVJkjrVQ6NkPpD9hkm4NkkgrCMZnfgbNtloS9Y4W0JyBQFB/UWH4uy/QrLu/UN6mJKMbO0Xa
UDKU3FLMZcTufauHGr61vICWUi1bAHDvC2C7d76WVHG0oHqim4/H5xPgECDDuijDJ1ftxcC7B4Hs
n1pRXmDHBMPevRuM0TYgDclZQ0dObGaGgykPNL6ssKLl779ohoxM4P/GPxrQmaUHlSyvKKr3z6Vw
UL0H/oN06/35YQrLKS3PDitNGYQ394YNljbAE6d80VK3eOmaAQaq0h0KXU35EWA4FYgb4JgdFA1P
hDHMAnvg5xgqMXIUzUb5ceJj0x6F2zAdJL8NxiZIf2SK31DH8DG+dTHh+twWjolGi5tzAwMcUMdX
KsVjUjDDxs2wLt3zYe0EQrJEjGjOZ0h2SvbZSPRr04bNM/GaHaoTGPDwnlVhkGWdRgU3n2X2/Hyq
kjikjDNApgDurLTLplVMK7xwLC4gpTL6gp7tQPbN9ab0k4LQ9rwtY8PmSfL8TiUnm2NTP9Hp30Vw
hck1MuB5lEYjWMwyOCg/hzStPAVswjObGf7meH/BwXgTsP6KrJSb/1PsiOq3NUsp0VTuq6RdsCe9
qHgbfITuUfdSKnQxZa5Hv57tjb6Og/Lhf3x5h7IIhIUM+U/itojvJ8jQXIAkL7PnVyKSQcYdU9uK
8bAShezyck6NemWhAIDrhzge1swvpVTJcPwhQZtZGMR5dMbwj+ood8jazDe/P2Buas87cJueIS59
9ILXeDKjYKEwn2H9XwrhROTJnu6oKuDk+T7e6jv7GQHXFxG083iosNmYJYPBLjXEmVr3/fWqi19U
fj6pcM4F/7hF/hQRDuoGv0yGOFT7CLGTIAWaCR+c5oEro3bMcA9pRVXAqZirWPaj75UFMIlcansO
aoQZP7Fd6sAswPI0Af+vEZXrlN3wIeA+oHxnNf50D1crqXxurxP1X9GmVjPaEPmXg14FE6UK9KKV
1+MDaB45DoymH7xguifFOLZGSuKfoLSh8zDqZiHlTZIebs7iDeB43A1LNPD+2D7G+SMTBg7CNPs4
5Z5uRG6Ghfp0dSA7rTPK9ZtZtjISlsyt+Ebu7v2kG10DhPvLahxiTqpewEgsOtqvAQ4xNe1/riRD
WqwbTUGrZQiLZ1yY5AdV9FMfnUGlH7V7th4iQ9lssftpSdxJkMmSe45Y8jvMPRim64VV9IcOYw8V
Fqg9ISpdFRRCRDhiBEzXKIjrOsfSjifxcK2DycEelor0Dn5C+V1QBh+HSS63Z4x7T6p9xE6YOVbM
Xag2bRJwn4ykg05Uxm8gDDpp+diKAuN34RiDysRJn2cDlO6CUdJFvUUnhhZ+iVeRiauk84fHocC/
jlpMVHHhH+gf1b98JQ4GGHi0g65bQ9tm265pSuUsTxNgzE6asp4imw6Npz90rb5A2l86hUkv69p7
5EjMNF6lkfYU67LNJ07bk65xctBv4Ule4tAsTwxIc1tu2kHfa0xd2PMX+M4xzo+RHCDaJU5EZYzN
LpADxptxvrGY8D7pRMk+6RqJ3xtm4hQQhI/lZbRCJzNjFQ3w0Qoeo0uVV7jaWibJ9FBZwPmLMRPs
om0PjDhMKNRmdNE0yN05rlIvEJAx3S+tKMkxNHVxiU3HqbOTIVAVETwDBsSanOEm88Uxm8cXecyi
7rovStSxzGVx1hGT9+nRYdjWDRuwuyVwuhOkS09mx6xsihgqvX6Pz+KyXW1V97mi0Z/0wsjDmh2i
8WBFe8zSip45C33d9xLtaFqQQIb+2NgB5kv9WsNZeCX6UZaGuy5fidU/YTvwy6vLlMlSC8dKD4f7
7ODPMbSZswaAHGvVPKGGVIkfOV9vMOdu1yHeeDj0xcO4y17JN4Ub9oDJCSTWR2cnlvAVoL8pM48b
FHGhpNvGeQII9rTJ7CnsBDLEaRHnnJbLth0uuVrNsBk8hDHtO+d6bWeDTs91yKrt+rAxV7V1DPGr
U4EMU2XDVQBrS6IldZYJIS7gycIU1JyIUVVZS+2qr+DhoKZL4DkBRyUu6ZS1+26fLch+SQgGT9Ft
AoPd5bfU6BFMytICDPK47FQNhLSccQWLSZHzaTVT9RoIJlSdce2TsXYXt7BlOgEWnTypTgT+pM+x
2E3gCI/fuJ4zszqTFN2znyUIMbUpIdaOvRIzDqH+Ui+5oPbUPDR/pboayrhSUS8Djs9it6trym/0
bhWG3bjSNE0ttPIvRPbSnZZuBXzhvgiVJ8tCZ9bJZTI0MWnfMrGzAAwPH+ciJ6fG+TuG7aYT8fUx
woNQOdJEt3saldJexyKUoK+xebByLy09t9dgDKjkcftD+jilJBdYKDz1iEMSsserdsxr50FCyQa0
vq9db6J+t80YbMAGSz2zJPXniTew7pBbe3PRwt1ZoBBfPMgs78MuOZs8KPCGoQHCqL3qZD7J/6sp
zgTEm/smMNcMa4ANsIT5wf1zWWBf7TPD3xdH6/ieT0JaY+QA0gkfnVNgq7NPaoohYLtzLJ5+pkny
V//FQs4j1lqIxSSbpqE9fr1iF163XhgLvgIEe/QrZ5IGEJlXF1Ae4TnPh80SQbfGBxbIOYexQdNR
7K+aX0BoWMJTyaMLXDzWWvhY6Dkx7sJ+b8gLKmsT4bz0GjOUPt8zOjkqnkzXIBqywxBf3TC5NBDC
OVvwgUokMF1pV/0gs5lH5I26ivvs/laqgORhzJYy0m/GQf+TJQCfrySTGZAGD5Cg3fe50JEpCCOA
EI1T4lZxP6/AN2kNHVj/yH/al/ByuoWVkvQ6sxVs5e361pS1YMFY1/LMR0b5IU+d2BPg6TijHsL5
1iX5AC1go/Lbuq3VfguYDjCu1C9Szlg9K+LrI8/ZMmC7OyfZnhVYfKZhjvsPSRBRs1/dJkO3DRtc
iCesa8YEP2jYKBDoGMwsgyalwvbqHU0MCq8QKQ92xODi/QjHNoZL9BblqwI94NMU2tl4JiKcsXJs
ctPGf23UUhwYPUImseW8PpEoL4q1QM7WRBhgxSoIStQKtiBVkFf5x5WwULr1DmvkGSvZhYFDfLz3
JgAAN3oURWf/6OYu1/LScU/jJU9eOeBIdyUbOSEA/RRAk0fh5PGNUkXUeMTlH7bCublpt7RHjetu
sX6A/G19mogqBfx4yxb0PBskErm6NTebhVf2FlD+ROa0I23bICKo8QYhgoYtaHBS1smDJtd6983D
kXQbFnP3gSPwKM5p7mcZC1y/iklqdOPMhNwaKoqze6fZa6kWCFjQSygf089Rhdy13BowAV9+xURG
g/Aim73G9MEPV49L9AgZQGj16xPCAhPN/VUR1uEBw/p+Jedhk6Y716nsoOBLE+ZUZBJu6vFE/ARw
LSl4lsIp5zV4ADTypRN3U5GXJHQe59XcPfGCyyTxT8vqsCAmd/rJBjcXLG/RQISs257EYpYu/9Zj
UUwZB++Tqbcf5ZUhrfB0DSLiOu8y3oa4dXG1RYax6y49/DY2fa3xk+dOfKaJpQvwE2+v0eKbAX/N
5GKDdZPDRbTXda+dY04wxu5CHlLgDMkoPtNlMTzKEIqDWlSIAB3md2PMYkr+tKarCjZ7OxKfWgiC
i3OlKVEHLpaiHXrVh/3yu761igM6WA070aJoYg7eQdRobIb7Vea1MkDXiTW+4PubxyaWqpAEQr7B
8mHeVpos9mz2qmAWxePc7/st/UhMnYB0ZRpyOwLeQ60QJ+BOPelrENQjzTPaPuAkznNcBVDddBp/
rSj5PahuxAfO3R45FXfjfjhJGjLBBtuLnx6M+7a+y4TJYKqZHdHUhXdr82sWYUftcivKUIE3K+TM
g+89P3XN3+IFxW816D/oB7pxr9tTeikYD44QdMz4rX7TQ257dnQrHiKrSbwT/saKNfkugGQAm2Jl
tGi0tj1RapQJbRtiQEcQaVzQ2BT/r5D4T3u9nVjuRtO37/GVl8mpHEXcBWUHOomhkcu4PDJfluJM
dVMS6TMYL9LOYr3HeAJZoToqJsg7uHj1QJMrMg6KaqjR1wvmLFr635txBKZ4le2vNsu9eMRmM/n0
MW9VMa0dcmbx3mwxMvOEeSIWsvyZkCMU0KX/ugBv87yTvH4x5/GQZ3xQ2e0aQ/DlR/ARdr2OXIiT
MV/UMvLev+pXEEjHxiiTIP+8/G7LPEHQHHOP8jLp72Z6dxjX1AXzMUe573YMI5eM4bCKhyN+OzA9
UesQ8B2tMwwjjPKkyVX1o+Zx3NBKttfpAn0T24BhbEe6nmOVrwL32ZvtZ0vqJIWhhVfdrWtJPize
51kXmiXhOM+ucaTFqa8w9xL00YuGWFcPXa6fTcii4h8E6S4t1pnvj/zRkG1BA/2SAkgC/yuTVBk3
7v/NZglvQuidpnMECe1ZJwbFa7EgGQHU4sCUHKNatnhkwmTolwKypy8Ia9QQGGyTsSBlb6V/zwo5
EcpoFKaWwgl61JxnlqGMo76OqQp80b8bg/fP1dVuHKtZsooDXNoXZfUdrdqcWk6f/KCHBdy+InQY
yJ9Kcu4JQjDngb35FlGWHUzsyERIgIo/kPkomSMt+9XTQFRholrkujrhlFeDBGTsQjuCiJmEG0SB
z6CMtiCSBhaiLclOWjNbm46eW60J3uFEIeCjjX5kkc/ST7VGbOvOSv5BEQyUDzInFxqnToT5Z1sd
sroqHyGsNRoU9pxws5X65iYeuGONV8PcMHYx64R4dd+yFxRd0qZLhgIiq6g8JnKXtB1KUPTBOo/R
wGW/5wgKRI9eB1T9H/+vjjQJeAI9wetrciSE/bacglNd/WmG/cV0YDA4bhtWCnCAASkD01prxDSY
Jgvw1YgkbP8z6ObPw64YcoaOLS8VjLwwAgC8cfrBkfUpeLeJwzBwHvCVnKxWVFySCJJogG4H2/gH
ph6pEflU0meAbcCvbUF5i0YVwRRPA3TVi/E/ZYaTx+VM3tYGd/A0qdPPVAM99CgEcsKmZLJeRGXG
r7WXVBHj2cJ0et5o+46zidSsDAN/+kdIYs/gOgDgms0VeOBCxoGrBXC+QKgBZNC3sonkZFnJ+POC
Y0i/F7j/8powXdulroM4SeBum2YZtMNa39xABZphZkmj3SAN5qkLAII6dtUFom2tQap/0QIX2aI6
2qB1ZqaIHfNSlTSCjVwb1xGgIcCmKEOdQt1VcnwQRKd6xhPotG/dZJAlRAFkFcI/aCOtvhjwvPeV
en2TyYRFOU4hP8I5oWooj6Yvt1ho92cFMQNa5MvbKPvSeluPfmcudc3+VjkcNLYX//HzC1dM5+RP
BipCc7NMCfPvpF8wlLQcMscwgi3DPmg/v99l1FWWiPBHAnYe7Q3THAwkPakzof4F3BIWJK5RwOtl
9Q4MsizJNrgGiZnnVF9rqDUWAUSkrt231AQYcMIQ3ZcTXiopPP9Zkd9M7f535ynJjY+0xsrIaakN
4FTzGEopp3clga42JVjfUbg2u7O/l2pwDKx5V7KkPDu46QnHI3jbEsjaPMzVpZTQ1Nvsi6yG9kbg
/fEadnfVvh4czy35EQ+Z6hwSss3YNWgobKevp+kCrThHQk9e/wqQGGxab5EhCmizN7Rt2CNegp2C
Q6qExw8+sHp4nKKPleodPNGX9rY04rzeA1pJIburFQVuEPWQ2EUuq+Vfi5THGg2WLPpSRNMfKwyN
xpnIVH9SuGReEcRw+Zirsy3bhOIXRI/1dDSF9wmssRgLmPbWyrJp5T4r0zRQu0Z27X5A+GJMWFDI
2nQRiElr7YmzY/08ySTAe06/s4aIbojcIbejf7bTZVYOFs7cpIHC+ncv94RPdsac2Rvx3R0Pfrwo
FhCCGSR0KIExQWKAv0GTQsXM/7IuniZRQ1AjvfA0qT4QOTZtlx+T7r0Awy3ZkZzP6RmWMqszvMQr
nNgeGxtfDpDp8Go+/Vb/7UV+fOv63jzlvJplNobs8zq49DAWNJbY96shM/82sJUh+UOMyBbuCCkG
HhnEbei/jmHx6lzZLXuQUF81dANkkD5hrd84tCmRQaNr9IS3nd3oUAScDParsrexSYM1xTQeVr93
IdBpN1Qd6Zw/lwyd+yv5SwbnGpmrx6C/QCJPKtcu3qXRFe70xR1G31j6sm6xolHwLmx43ttfFYMn
hdm4ZsDpv9SIATecWgep3W54QO1Diyjk5Ru9JNf/BhJn+puvMCZSlpyrq+OUFw0bUhBWyUfNvEgT
7VwGFhPioONZMCneaVSIqn8GnrxIr6VqAXGos4+p3r3bZnu/JUE5ooefx3y00dggnlogeRs8EZQ0
WSLGHEAUpBVdHeq9sl2FFDOfApc2THZVVnLIT6M19nxAt9/vwqHIC/ddnwfM9NkcXDbqtSFZxMUu
FDAPhIF3endWZLZG+xe1w6ngxjCLGA0vISFHgYv55erqSxR9DS99FBffqYq4uGOarygpi96GMOs+
CZe5wZcidwdHc6jRTlZijTBte0PBd2fVhGLMXVTqyuelnUblKrnkG4ImTqGRIdqTqOEiGQnt1F5O
z25xErBGvVGFS/7Mese/KZG907GObQymSpFYLoW3NSkZaYeuOSJ+og3xsZvBJ5ddF7a9HdV0EGIm
x2cG65A3J52hg0Uoiz0J1F1lz0jfSJZuFbFUQKaWhxho+tg40yhVJqedfc4CNcADd9sgUnFxDsMU
HsEIPO2kyuYXczZej1cTJYHjGmU32zojGZgHPa3GdItUNR6nJbhKo18QUJIiWFmF/wfLeVmHorw+
TcyMLMW3r0J0miy+XnI3ShcuSom+UgvLISXWy3O0N900i6OgLh/L1W3NT4Qfiz1LHoUy1AQ4mL5X
qpr4pT02LhLyT5nyQnO619Hw+sgs5eqmU/0AuZAPgFmZMWEOhLdbra8ENBwHcfgsACrhtyF/mKfy
SflqX8GlmwP+eBlYJuez1yXl9wwIJmd+Rw7n2vOf+/dRek996x9wUuw7YjNGPtfhr5PVTLtElDaj
oGpiYEbbd9NoeNBSTzvmlHECcrRl2MRt5DxIACnqWLATXETTN/xMcHiT8vZRTQ4VL9t7SPw2nZ3L
khohSs9+qUaTk3oYZrBxhFAiKx4W/kmmRerqFvPghNOjj1Nf+vp34/FnwJ+wRPZQRbyhEGTIdqXs
eFtx45Ffe97d95Idup0LwUUXFSJBzkRESPl4Miv9+6QsRykUaelVUXe5VuyRJie+zfFD6pUJW+f9
0xrRrdKE655DXS+0Cf5cX4KVXZSZ7cdYHmOJxJ9i2oF1j4akTjlAX7P7dGYDNJ/gNej22qzD+wWh
TEx8apo+ERM8++rkMZItd+eV97P+0S5CSBPFhNeTzE97t6Phsb8Rek0u5WqRxe5OuQWNSXdLZuax
spJ6jCUbb0OvBu0uM6kH2cXUGaTxAEKaQ4UoV5HCDYm1K7CWVdYYuLklV3Q745RBjEy5ByrBzByx
BXqJQhWzYorY4DwpkIWR97fuFF6hUIrJaR6/i3Fip+c6rH2JECTlnuW8zP40jLk9fUhqOYoC3/yy
KJ9osrCDp2ZV4hS9VsQB72ZklKcMTc0m5l/iV94CrKhEhc8S8M+V8StXAVvHBd8D7Kw20g1kwm0A
lJTDbLw3tgm/vQtjBtaEisIjDqNe5d3BtrAPYEHyyM3tw2zBN3QBSqJZ9GJRKD8Yt8EDqgM+4ct0
/LYk4U2Yazz2HcgG6DZ1fQKvyMVymgrl7GbCXjryJrJPHGMB+w7704AN1IWnIdJ7JFHbcZDFEsWN
6WcZM7648MJqSALBsACttl4cxoAIZpwLI65oYuXis3uQkvbx7sVGPaanbxXXzmg5RSlnzkMEwEpb
GhbLBG1vKAoikMF55t1uQ06zrh4ErWb4egs/FS1fmxZHJ6nP3qb01VqaDUsX4ZWW/bTfAYec1Htv
tWT8l7SY9yJD7+JPZynfeuOAH+MoO9NyCdncXwdVFXR7qq98Mt88xi1k8k5wEvPera23rVtOrneB
fdwWYLEquxwvC5+Kt9KwRf8ok0i3yRCf0AD61FdXJYwGTtqSuaD9LjXHV4ArM/UCd2P/I7p73eaz
H7sS89EB8FaN88teBOnXpbMvEAmroz3Jfk4JgE1ki8EUZxfmDcMWpZ0QgFRhagMWZseg9UQC7mL4
oZE0WCdzT/f0SO1RfmYv2kEZP0edSc6cx3wTm1AcIKpvLfLtsdTYeeyothYP/3GQOVHa26wvtx0x
qhpq4AhfNSARffEBt7dZViQhvzJB/vPuBzESm6/1xBY2VEXprbE/x82Py5aPpuDVuLGnIjUhBUH4
Ad6/2CMEIr7tYO94oaiT5Co6AT+jn4GEJdKHUBlPr/l27Gv9D+aCGJ9lhyXTlkosPucIf/ooCuAh
J5BpozvbDwqVS6xPLcND9y86WcWfEMIupIEeEJtPDNhzVxghi0elRYNSGuS03D39k5GPzwlGiM/B
r6x/bfbcZpjT5uDIyRS/GTwzJPt1hz9Ggk8net1a/yr1JvMrWECcW3d4Fjy78/V1ezcvzA0aw1oa
MzZh2fJpzvLUZioc1mnkBSk0k6xYp8JhjLCfMFzapn2IBThHsyUrjn93zGf/h+LL8k2zbw8mwiCc
9IV72l6xl/o4S+65Mn16vr6A9DamJX0i1xAXA97bS9EvEZiNhj13YKmd+PIfhtEEwP+TF2O0NVsd
xIKHNlihjKoZGaQs6HhGcYldJ6ttY6H506Y8Z0QTNKFrz0Kzuf1qqd/f2TZ3euGCkAtFOS54rxgx
7fW5MaFZV7w+OpRHJipkR04hx59lAEvmoH9YSTFTZPyohjzCM/QdzzM9xGBx4NoFZs7+MDmoyGU2
pkGlMqdKfN1tv5bF9272aD6fb2ZyI17VE+vkQy5q1W2EUCssMiuJx0foGp4wY1PcbGTzDIkwff6H
89nJ7gwRCuwq6asHAwarGiyxUghCAxBN+2+MOyLnqEqHFCMp8oQ018wLs1dAIl+dmXOcdKHQpf+W
AB6hFwG71Nr7IY8pkIRzeBI7YvaTcm6UGOihh+t80vxA4+EvE6ORLNKpY60/sbje49HceOdal7to
/CMf1UFuLlsfAKsyXb4DuHaq+6KtwJOljQwmjh0pcydShW1fhcYOEu7S/oHvjetu3UTH/Ngp2klI
0bW/b3q0PLfS7fIU5AzrhskydRkmCIKRFVkEZqe44rntz3uKr+cv+xgsjhnwOCvG3jEBai1sjmfU
JiJeQewqc+m3YOiYRdW9Qv5oCdkFGygh0ewbf9u7Zy9KTDbFsvtAoubtzt2M4c2dyTUcimMrjwZb
nsw+VTa5ZvrYMSi6i2yUTpBTE1MA4/vy6huZnehh26ZxMqWEq2MRVtXCngSpSGOKp3zIuY8+LTAb
x5xczT34BcJPFot4u4P6qsvfUKaNX3u/E8sicLM/b5N/1DVxmuY0EwgNRKVA3/9kO1gWhNSB/6b+
VMPvBntnW063qdRDD1kyhxvXm5ipbVb441ektCehjAgUI/hKIdRy8Mmh0C7xVaYR/bRXyb0sERV9
4h1eXz8GFaZfB4FSuR9EO6aymNDDjVddNAnitLVDUOjN8K69KYZd8rkkpdAPX/CtqMcQW//QOrZt
DSVYEJ9tzdJ+N5b1BCBJTJRW4t80R7UJaVo4AKyqbhps5U+n/A47K65PGPn4Aw8OMrTbfQq+EaO/
BXNbXeUAM1D14DHrwdEDdgt7KBDtGOTzpC7ldQwiPsgsPrXHTcgY0/rhN9ACcc0hTGpQMT8IgV/3
S6Xn+mVUz0h2e1thUFevyMTjBg87+wS8m0I48WNWwTjhvx3Oie9iZLEg9bJOmWQq9mEfskVjKyau
bcm+IdsIqgLL+McLNtvq1m2kOEuNdf02/+nyiVNb4zvVthZ9sV2RarT0iagrcc6ucS/liLu3kwtK
/2HVYv+p6teC20GR/cbyp3BA/gq4YX/WfGQSNYH0S5AYjtVlQfPibwEjaRKNkqDBoWL0aZdZQfvT
qBNaMyCJ+3Fn6C2axFlnGOJxM4UAKE1FmpDX6HWdhfiNYFD7PgCEx6oTCdPp5HRD9Ni38COj25Lu
i9egYMDpKJBw8WlZnrHtbcfmHrju6MvchG4WYu+JHW87q7b+bcMNyHa+HTwzjaIpJwxCJOI6bibo
wvsACRA8dANnpieFBc2jz4LgGP7FbAFXgZ3Pr+W1zl+oz0hCvmAO4wwFP+tx7gdjI8Xk4GD5Xazw
U99MZtUxgedZmq8Jcx/vuNaRGjrEw3UEIjq4jk7angkHTbHZUOiagd1sZfVNY8u2Lq3ikAN7/jES
MQVdJO9Y/6Cry3DRsyX3F5B8gkh/hC/Na9Sug8KRV89M/a/Oj69egXnTHix+CjZt5NpdEqJPjSeP
O9tb7yWo3lDIQkh39fRaKLzY68nNllbAzweK2o+Mh+UgcOLpycAiti+iTPR79o99bZr1BVyQjApL
A7XA9gtRyZc0Qm/HV9QiiAKKZRqMptjzznnLrwWiZG7G/z2xeo978TKcjzUnvAbTOozVvnasT+OM
mNrfbIX0nq9Za+1xY8dSdcmXT4jBQZfHEdMapcIQW5SpMK9KdrhvGJkc3zRXNy2mjbOCQT9nsOt/
IKb5h/8hJzm+AyxjXXeKUWqwP52paiPRtQQI9hNmsRhJXcJqFrX6yZPEifeGxIK/Pw2KAK5FCNBm
5kpc60UpwpMeZLDguKNMBnrwR5M9c3oDRJzYr4Mg90Tj5JY2GVkstha7LZj5bUuO5Gp0lisq2EM7
LmyQa8dR3GVH/4EgVIBdEkPom284VBsav04IPSIDvjqAxauhdICIltBOm96BdwdEfwdNpgl2zJNt
+vkBjPawiNK3RiyFttisLSbbMJ/19sivnEicIYY6v/DDG4vjw/6O00vRdNI4WRpBQWyvX4IxYRvb
0y5zmEM56IfSSpVw1lm7DISkUofmGL2grBLlolJMhfVHrF9+eqqndym4EmkHL4XtzoGb3d1qBLA0
eoizyijjkVcGQGhjZHTtFsarG5jZPKsm079fs3udKCpQSaDxkcIzhAQFB+42EsQRJWKeADT8Ft5h
ZhkBrhsGL+4+UO+clXldNiVrSADObgoqqdSkEm7pqWBF089dFCHOsDSSDlihsGMFjrRtawSkPNqA
d3O1styGms4hRV8+A9PpMGGhlfrI1txFb6U5TRrXFpCH6HHN+0qsQweMFgS248CfW9depWWV4mtv
ZXDz5Ja11H5+rx1UmBzKpf9Hw+YS26O2PQ6PhVnNTeMYNxTPxd4e0T4c1wnVVNapvhTrg463MevX
UGoFBQz048gHedgkrrVxlfPmoHFbe0bAanxKhpCPxn3eCuB0QWeVRoxJR6GMQlUzynjIWRv0iuZN
P7/+3AF5GfTPP6YbmOvks7Uzsmb4cjHMkivNJh3UddWxsvFFjn5zz6xYUYBktb4S+RmQqqmH+zGL
fZasVSUmWq3TgG9OPMd8qzWQ9EpRCb9IETOLcl8kbYFUCNO8NMPTlPQuzg8KTBXL3yDau55+vg6O
Zvp7wEr+AK5+1srZ+LTayaNxsxcevvULH8v5AwQngkW9AKQ+adURPCUlfKKiADyF5WOvZlR011WL
b3RisCL1fPFNVWo94Nu3Yl2MbI7BwbEGfAZUvb8Rhii6U7N/wEDmvlHP5A01Cm1di2ULui/kb4xD
2zAP1L+rlMOT2d9liBUbamasjZwt0hu6xfRZ6ha/iobr4Dry0SkhDJY9ZasL4mBGYox2YEzKSVRZ
vaeLQXDW3ilWfEaOgNtgu9TRXZWUjJld/OuxYVCf9ycFqhX8Qqd4Dao2NwHnQ59U95mZX6Ob6qga
i8/JVaaXJxj3bKsa5i5eoC/zHaDB3sfAzlQ+MPZ/LnJZeWOzhB3rRfnSiheJBfBF+ci50PPl2Kme
KViOG7JRMdwKh5ELlFvIhZDoKaWTAo19+eJ5CvFoxYy1IbjqeroCWIGOWeJt8Vx8KENdjYs1gK2A
0i1pabQJLY8wV3o2xiwChibq3bHFlHO9CmJE9dshGI0Ymdjc/X6fa0b3/Uf+dJZ2Ybd2NCoTSb1l
x82BTerhaynncP9oe+IAmOG+YCf3cMRQhbZQ0i4IAD/OqhIRJD1yWdl2tbRgpZ2K4TwY9OLCwDC9
PW47bi7YymZWtAiiVyK5943ji7HVT/H8IpdWd6uzUl94YOhETpPeoXvWTivhZkOcOJv5u81P5Hen
5ezd9Hgw5oss4iYnEEfAD6wY6O8V9KCqwlRCySp8t6NxdkUpt1u3fimSql8E5oO/dqwEV3z0XNb2
Ls+6J2dza0iCv+S8lHpUprjfx4vJPM4McicIGTr/IeL3e/xONKLjLvit3p97WPBkWh9uOOSi9goP
mSpLXYQIFwBBAbIhT0b73gfuiOm9akPHt8WWbGvKJpoJHY8JDo8Vcp9ltRlorWeGIKRXZePkNLne
4fQfabww8Z01o/N1ncx5Lo1rVeDtzs56WIiHNqllt99VdhRhGISp33OobOiD5PBLjVeN7rnnPIpv
18c9QbYNBQWqBWLLn+OBeYMXBqkxZYIlHfff6xQbx3hn9D6ornC8I+2GEPLQ/LikV5Icin+UD+4w
znvhyvriMXqjXbNf0ALWJlYDjBUdAq2OiO1Vki2n0EhOkgiGi5546hmnPj65Zlp9dEsK1uhJSjCV
V+itiDCdRodVMcAyUf8/BvHbPFo47Gk3Ueo7zveBckZZWwA7obpZgTaMopbKyVhhUOm15dXS8EnF
9mQCImthOYupH2xxG1T7SXUCFfmUKNksirx5aZF4cMxOeiz7Id95S+dnEKfyXLsco/YrHjOZcE8p
DkGS5yFpR2r0/0WXw1SJ0cURvky/di6Wo03jpmLZZhlkP5O4uxmmLM5ltKVal5yxkQgdv/HxZ7EP
1Z6DRD+FF88vzM94ls/nuQw8RBF7BY/X9KrMPLHrRoKJkA74WjKKSocq6MGe9X9dRo6Su20965Ko
8ok8GGZVbK1dnwPtybmqOPke8uhKMNVypRL7rkj78oalTRZtMzkn5qo1OD65cpaEdIUG+9BGFbof
ibkmKW2pKSo0Y+de3HwCoUuPiUtWAQ8Pi4XnMnTFJYE4v2a7hPRCeJAWQ9/BUSxeyiP2sB9A53Lq
H8VkHGRsiv1eghh3z+Ba8KAkqGL4Zj5vJSWeB0syuhTVqlwlD/SW4J8t6O7QqsjZ9iW/uUlx3IhJ
x50BuIpWqXdBP4hCaeyJG5mZzycSXp5cdZPpR+vwwKiEI7YKDs3uo6l4GeaRudee15Zr0dn5n7iZ
maafVlBPhmNXo3RVHmhG9/OYVbZi0zdFBA6EmvnGS+R6ZJ3xKehoo9MT4/wArHLRu4A+GDoHI+7X
brds5Y2SiixyD3etssDE8AsUcMWt26jO4XYGqQkir4U2MWRH3PNBfuoHlDbZEO07lx8gv58cFFiJ
GZ12DXWOc15HwHXqqLDpBC9xonbqsNryZzblnC0Sl2LDnHhdSG0A7Ne+GOrcjf/r5mqCHVi955sx
oAFtkcO1GJh4MznSJJCTkYhIWEmB5C8FVJ6MQXpA5/45k9tMGCYZVuynarkfa0QU1hEjsYtGAYyM
YFuXi1N9k84nMUjjFk2ZFeiU201qE+oitbmPt0QN2wRMFwcQuGzRHEx73CdsqPss/j1wK2vYfFcT
EbZgphwfols69BE+H4R1p8VtH3jqPHZ43k4jdtwAUjzAUGNqUX0sl7q4xXolliyyiD2CyvNMy3t+
edZ5fGgD2/qWuDySom/o9SSI8uVS4gdBij2V8/HhXqzr6lKl+ZRohttwcE8lgye/nSQt8JLx4gW4
37T4Z8rz774Vb+XT6OHYcDT342Ig2gRaXjju1QUAWnkVTSCq2sskAF7kBipt+rdtTZ45mwb3m2mO
S5EbqknsnyeOhwFFYVEM00VWkge0WC7ZBa8mhihbFDVZF6/1/HkYbSgyeweVO0NnL6m+0qIaSfvg
QaMruqT575DPTBqti1hLazw02TR1JuY2EMm7MB8CSTIrYoTDR0+ykqLL1jReqIWajaaanSPApw8M
9kvV3aWv2lmM2xuJYxDUxFAsekTupmDffrGgblJL3hr03+hy/iEwgiX0yMawls84VZnbHnQWtbuo
Hin98v5MIsLyiZjh1h2K3w1/qStqXBskvqYDOeKrlFVMvhEBBg+R48ZISQxiZUEknSz/tVS5ITq1
E2jh/nAZz/I1sYeO+FbTkhLVTgX0x4ZvmUXON10DBNSfF/+fCvYitLBR2VotF/jywIPQI+r+oeUg
urMOckZSfjsSeCfi770P6EzrvEIak0J/dgszs3OYsUxlL3ZETBdAm2ITriCPV/i9QtNM69mkrKPh
N3HKJ/3lBEgQJwBq5rG7DSb+jCKOdwvM/ihdotQw744jeXfGUgxfMz11kjCBmsDb91LC97RGTlFi
310myQRUC/vIrRAkLDFnu5PpPxlVikX/4MZ+mAoiSyzlgcw1GVaU9C2Ky/YnH+VFhImEJ1sfwnMa
gViD6i8jYkb6eKteFFz6nJ/jspBb8M16qPhA4YsDLE5IpxSC9AuiJohdxqOiPbP3Z79ribiNcjsq
hOj4SgtG23rEXwJaWonXd1fl3/djWT48srG7EILxn1LJaGlM99WqEsPZZxgXNf3riGHON87B8s49
YW0T4DJveDjyWtnBbR6gmeOyFa9oXkASGCg3RIETu/PBIWCa35Ks8kfk+FRYCE5HHUC0aQ/bbsdo
irLYIhNrQzc632HEw4MlHinFDI8EGBzwnR/sx35ojMX7XkOnbTnUuTC7V92ZZBi3bf2gkghK5ozA
WPRKnfD9zLWYejmvBXUAdTBX9OquenCRXWru1/Oc2HFLbNx9o08d4xbx3xspSaqYYmUYoDPjp2s6
33be9t0UmGzGdYl4qpPoBjjzeA3qdddBSN6EL4d+iqGy0qlHhxId9LYSUDGKxn1fvz5T//MX/QSK
uZP9MybO105SecXN+nB4s+MpNBXLlUeAICCOt+IWAMBrK1rQbgb5Cx9rCIEr70oVehsAzALnYL4v
rMbQ1TqWOksCL33RpMJva6I6upfUjQmJ6u3JG0Zn9x9kknYcv83Rixl9VZmZ7DVLP7BaVNCfgVXU
5Eq4iPrwpMG/LHbYTF781SAq4uuzDZaHyx6tVUd96BBFO67ruMHk9mRvalaDyoP5WKB5WZHTPgL9
HSBTcf1wJHuiRxYoFHb4ft+qqMGO7E+od30hqq3Fhofa0uhOqjOjgHjR5RrkNOt7odRu8M2J2/cj
6QrM6IvLa+09hLp8qO2DsBr7Ceg2w6eu/dfjzEZXJ0+vG7MUtjG/FUklFHs032U3YoPCXYIKC/r6
HPWQomx1uqRIpBWTutRJaUMaeq2eXpT3iTIR3d9/PBvVEsgY/7nJxk26MOfooNBpS4bEJXGSzuCI
MUdX3AMnqgNFg9MR81E3/6ryWyqBS2MClSXSF+EpbiZR7VFe+fLoJy1cJ2tpbr9bD/PeJEfFxPYw
HVf9rNYpU7zt9cbW1pc60WlkoPXqzpH7KLNmk5xujJufV8mOLfe67M6Wvraydsb8ioYBA77cBDGQ
0Fw79e8j6KwAlkm5gYVA7ARYHHI5bUo+IL64wbU2P4RjnfQTMeAQqa25Jg4/nLkHs0mPdaBysfEE
88zRhZxNYimZxlYMo6M+3BC3WZOdvoKYvT/ViMaz9Uc5tPwfmqenGVZjPCCRo0nlnJ2WO//Y21Ok
FQLn5d2o2Xub8mtrscv4gGLXP6qMUlV1WSrrAk8GYlJ2jB6HdDwWXjmMAnly1yYf7WnBlqQZwpIq
LC1chNXg5BOHxuaKGs9VoFb+VHRdb95JbLqAQTxYvZ9kfY7doq1Rn8tVgTEUkcM93IHbqx4RDAkj
+Wjj0glvhthiQajlLCdDhPOwRV7bnxh4HaSH8PulYygIPAHG/0B2MrI4nOa4Ag8lVsZMQF+h2oP9
GIfbTVxmBuhT1h+SPvELfCdI8yhKM9KOPGsNAaEzNEMA3vwlpVPaRSW/8Ls4ajTkpWg7QhgMIZGp
sErdM3K4KCI7XkxC/aSdUpaepz9YDhHMVI9/EIys/UiNLHjg4cc9bN69NCEzw2F6V7TXYYhUPrD3
EPfoXEBawuc6qNPAef+ZiKuLuh7fE8XCvY6VKV3zUKBY+NMbeK42HApUsAEyYfBMaeDNPEAFvcGW
dmsyfgGJxMxvX47qE9X+uMamdPeZyx+CWOYo/qqrw4v0wJ7EZtwq3CpvWz1l+ON+1AhdSFwY1c5m
L70o4cdgXhjKErsvPNG9gxKr+43ZmgooWL0bRC5a8kB61XyX3Bg5Qi7aEN0cBmzqij3YnrgjZO5m
fnoHqfuYDU0fB0opBxX9csD01yd3QQ1rqc7bIvUQeGvV9mGuyzG2Hz9hux8vH4xVTLLcNF/4AMmM
pQiMcdMBremVrwZ8JdXg1/f1H7qm/uqU2AI8ySnD4b3t8SWV4aPfz0IsWVpyqNLpRWY9TH8xVHzC
ruxT0q69vVHYMuC8N5ed6q2Z0VGYMAYjjVakhq+u5i8LjGh4q+jrFGAe5EzUHSkb7/SFzJ5XqoM2
7Z0NCS8qmY/OMFt8uTn9T2FymnvxEeEJezpuVArbQy0G1S0tm5QloSR5CTFLjmVbk/n1v6y3isJI
SPxPqufFI7HoZ65uDkLfKu9VUHYq6XMM51Xs2knKAhRSYtAOVn8GxcF6EhdKf0OwW7ioaosGfJu5
8kaOO1YOjHKgtSKjJin5qt/ykDLSvqzP8oZcvIG5sIWRm7UY+IXgcqozpQvhPgU+oEY1odEVJH13
5XILPpChqCkFdT71RssxPTMESBk9ksU1QKZYacXvMP2NWUx80zvpfhKs2udHtH1lnaSs+M62fuaT
/jx0SKhT0FaLZ4/0axVG6Tj0uG0uHcjM1h0CxOhj9toSnhTA7F1YAl+7SKvc9bZkpW6we0jUZB2J
agzO/7JUDr0sQSTtqXFtL/UtLjD9aGhZoT2wOltBMLjSkurx/775fZS81rRiixamwdPeCCFMkfvt
6LcBMAu9dOL5cs/wAtkmCNOPXNygHJ9/5ktuDJqEuiwOzYcZKxW1q1j8RAf50NbXBspijqdE7ahA
OUDCvj453hntZ8J5SIMUoLuLNmVIE4GjC5+UOQHDzh9pE7PN0580MgJkVeJrM9+//oeA+NninnnV
7o/sR1uFMcrvpZicxiSJJ/Xff/bWAqAMNmAHl/Y+j4jTQovERCZqN1bbT/UAuPXBN4jwVivcL/Aw
fdNi+w0o9tolrSE7C9SFL/OAQPRKrcUjtwPkyYMVRyF/6Qb7PK1fR8zFgBRAVTuV6Zivg+aFaMWg
PZgit1FH7QbEQqLmHXWfrdpBPZSZXuBpU/b2J7Fziv1qcCcSBjLaGfxmiGNa8K0ezqOYJgb13Ijm
XrKHGKzOrbofJ4sMFEixKujHO1rN33gD/pibW5C0rzaXxfNEE6HUFN0Hv3/QGE0Pz13EfCgzZ72H
9N/RMDE9KS+XvRoFvBPj9A9AFqloShUpY0DP4KdNcXNTt6PKc0G6tp3IIajYUQEG3bSW/R/qQTqB
tuY/Rlin21bT0EGAoXgr2lP4McIluPTKiuuIbBd3KfmJzZIz9oCbw2WY7d65jrdKU1S2KtjHWueE
Z98obJsR8cu+mkUF0aRNLaVIg1+HYTntz98/SmH6PktsAzt2d1yA6PJqqeW2VyVPaMKUTs8EY+Ed
KSJkknMiNjvdYggskQqJItDcdDd6G8KgGsPUqli3a7wrBL34k9jKcPKllN5Gn0ClhbDSFjRW6UTp
LOBdWg7CMGvdIu3rnu5BYu3/isJLI0h1xfDFKKxCeQRINptFwhsi4etTeVvq2xyiqkYjbQ2I2mXN
jTWtQE6P833reDG6+/94nEtKxkrG69gx2rOlE1Yr/FBwSQcbYUJshvWOyrPEq3PzIm0VSEwzQcfa
W0rABXtrLmmW2236LvRx+su1KzqCSPj/3RKlXie0U5UOCcXhrho2fBlF5ktZpoDSXVeIJyUtbTpg
Ao/Qkw4zVhYrI7gJvtkDfnwl8Oiq8yKr+OTCK0ygWnutVS9qUSe308BH8WnXd7whIM0X7Qw0cSgp
F+jQf91uVcNGbG5/HPXvhC6tChHtdKcw+XW8l42VTQr31oNGsqIPG75sq0Ju8cExThv8xJPO2nb9
mMtWJgEvYGZdvN37wlvqW2XGFLRvtSK0trJvGxStD1nN6A7ymxkCYgG6V09uHn3H0XV5jU6OOnB+
VNxk8BkJIO7cAw8t9to5YZxkTZ/JcIFigBfQmiFfem5UOhBMNdRhvXzlivE6N+3//ITH/m3P1sSN
hDJaMSBjQM/O393a6w0AoXAFECn/7LtN+x69nqRB+BnXJKoILQrv/3eLJicDd8j7DRNjqciIQKFE
SElgLZLFwmTkcZ6skC2SCuHhfbrFcbUdsvrXbOoBQlri8fzGtDl5E0+r/xQb2SRFdWDY9TnPXGOK
wJ5G60J2XTdUvrj1iKu6BCK11sBFNF256/LoDKPIVKnI3dLKpyCbmktzgVtvnSc5/hv4HDIuVAfp
zhPuZDkbSeCoW5Czn/KNsxCBDvinI7E9e2qAeM2xqiQwZRRCBKcAb7/Vhnl/vPQtQhMxtRQ64D+w
3ttSRs/7uchTIjZLtuSuPYjjsRE2q3zQ2ixvI8cFGphVuQ0UQcT4xetSCGf/4z9WtnS3BKhDxYzE
oCxTZngRBKt48Z3MZaMccn1BZ2BeSm9OrX+eUeNjKbVnKWPzyD65P9vvEXArFqlHKqwmOYN8pNKb
PZtYMw35F452PTLnNqv1TAcG8sGMjrxsNxjxnQcWlk7RO9xuFaU+rrtY1w/mXx6rFGNzjrK7/Zdl
XBIogYcaCtnqDT7YNWUVD/CE0d+3iOjRnpbJ6UbNYtYc0pityVvXGA2TJOrXhWNP9zqE71wmIRvF
nDQYKAxPeO6ONSrPsRIHDRhtjoKsA9bA5A9xOKDdEFxeYHDszZp3svJHVoAXVZ1K8xZ7qNTOaWjv
Z0hhNWXhhq8KiCEuxw4UYRTmaR6xpCsINWRvMNaSIONW1BwuBICtEljkSqIx5YGB0FMhUlVGz3iw
t3s4SDhTuZ5lJ/gj0ppcb8opxy+a9QVE5N4mlWQpgOOwST8Q2qafO1nXuOZZRdTZFuK7aOJW/5I5
GQRpmV5FmRo0c21NDwSDiQazJmCWUgkXHnKKu0doiY7P5xrEbwgQp+uDoSsS6chXQ5Zurt47a7B3
2JGx5Zt8sJibzn4vhw0gwpurrS3Oz7wMt+eiCTTSyb3RtPhzCmVtOJpP6KdjYOz9uod8ECIV1aLa
B/ud32EaWceXxwjYST4Ggmg3R2yX2SlA4pbm3N36zXuaRsrXXagyWixROSYfy5kULgiZr2rhezOU
n+wfVXTWbVPxYdGyCjtRmyo6fbnh8VvggZ32HOw/TxRgKCZsexVPNGknCCIBzI5+XLeR0SYo37MT
YiOnZ4l3t57pC3AeJn7du28nAC8Gb2porZl2ElfepGmLyu4jqpQNHBTzKH8i7xUcuVD2XPPqar96
GsMv50MLAdOFKw3nX3ThCYxU+AFtSGNjbPx7vrf603QZNMjpgrpgPphx9jVBD3crsWWvdJjBTb+t
FDTcKkVKt2hAzIMfpvxv08h1QZ1hoYw3R5Sp7CWwAHd4iNwN2BwK1keKhM6ctIrwZVkIOa4hkiRt
OaEVfij0ws8SKH20jMoq6iceWCe9AEDwD+cQWcO1OynXOSYzhcnBcwSbtjZw6a44EtDm2JE3bxYR
5zPwcAS8zXdje9mR5fPgRbufUgqOsUPENTesRrL7tPquqVIxq9Qz7ViMd5Bxu/0hKoqFIGchiRgi
OE6dlNEPHhROkOUD++jt5YysnbYQ/iJg8Gpr2XCXZ8250P+FwVIVD1SPG5XnPK1uxmJIudHOeC+T
hPxdgnMb2YgKI/kPzsUQqR5i/M0BvZcsu82Y5p66OM4mlJt8uZjsQXUjDnGg9Lt/zgaLJID/4Pje
nZyG8q8/p7S/jT9zgU2wW21K2jft55pm/cJd8JoumdBVhZ31Lc9+F/lWrq24ypY7uRC3w7muAdkR
iAZPvrASPpBgdk5je5THr/+g7ZuN11JWMSu2YcylaK+hR8vLCOe+ZNxA9u6Wujo8evq0lqI9cDjy
8JQhZWJ8zRKvX6SZH0zpnqM5ezZGoqRqJhqR7pp/JhDBCYgI87czIK4TkasA0wcgKJG0RiENC2iY
4Yglwcm576gzwYCI0F8mj82mlXHEmDLvlgeaFuInfRo+k8vLtKNq8vjZFCFRpi1RClFtpkNHIqBO
fHpurw7Wh6Btm88kNLmeDFyjDkQHamewRHWRWEoOeYvBtILMhU41fXniGB8po5xNuMMA44uapulr
w0cs7ZB6Epgww2oQ32TieryiNszeVEB7y7OHiz0OIrn+xJIjlgD63Ba56R4lDKlrsx+BUPHDgs9T
YKZGKXKj1NLfwLjjoEKlvUx46wzAijzCOTGVbz5rjV8VOEPhW/6aD92tF7DT5uiWcutm5SXY5Y9f
KQOTzSd9mGpAEilAMWShdlfU9d6vLdA042jQx35Blk9r9fUGfTsNcfzfoAlWmbcnghzvfHBBN1tO
RSK1r84CO1+DfHl9+pug9HHKXZoQIQgrsxcKJsZQRzoKkfzI5HOLhYs1KucGCLtdF150a3yQ4goV
C8c8kpxxCsaGy02T9IjtJNjcajnH93nM/k8265DEWyaV1W4Nd45cFtcb3cqDJCWvR3C20y1XHKT3
L2ADEiWS5jeAovvn9f4SKyqtH2Uml2fbo0wTBQOvO76LUNMAtVU22z2yqzc8qzrw+SRzRZEeL7qB
RGfeuRGv8SN6oCRra9TjimGTJwLL/9VQFz5+HrLUG5b3FTS3YssZbVO3jNJq5+NR8Ce69iP83AnG
xQu5OdW/3ZJI2aDZK6uc61+HbByW1a1wkkfsYNbiBYWiro9FWPFK/2g6wAxi1KJfiKcfTDayJDyX
fdduCcA0JU3iBHmQph+WmDZaUbZYbdAjjFN0qnDU8N/yBk+IadBaKJJHnXDWtafysbUAR/XG9NR7
VHgGSqy24tedkYLkySVCLqH050JysIL9j32WSEsNXhDcHDluJixx3iKA5+j6lYpvN5S2/HOf4kjk
qPK1rO5Pp4IVq1TN/ZTt3WB1Rof/0hQVYRwL9tznglRy2txFfntofcj/otQ6qeWqZrx9GYfYW5WL
+baOwSoFUHgz6NexFWn5+AiuQnBnX1jDTxh44byWWS44E7HH7YJsErlXFzgzCwk4ExU0Bq2geHYk
o5iKKazEabOI3CiefSJj1tR59a/5Mgaw3I0S+ztDYuks3iRCj5kUCkFIr7LpyFziY1o2uJMl0Mob
akR6OfOs2jVlyUqYDxtc18hSpckvnuw+8pR3TNcTVZSqY/luKzC0AQBi64NjbqAQOLo0lr6PrV2E
mVSldVij7Z47ur2X+tmpiEltcDWiEkM5W+aB4u1j62sTES53e9PpwnUczezJDIhkn2QiJsu2NfCF
qDtn7Tj4kj72jKZ7YDlR/U5P9tN5NOdKAF8Iib/fSzEGCrvO/P52tNHT1PAyxu2qAIfqr3cgyrq6
OPWqM/pz0xn4o6Ig53+SQp+pe9VpEu5U1xsq56FYU2FJ//NPMSAeXDSStGgTF/X3JomsT42rCTsU
a4UE49qarVEDFVjDSZII1tpokM51285WHD74EramT2Ay+1mLp4l/D9m2qjPoYEfn+WGJR8VAgoEF
O1Xnho1dqqt0EEL5eKhA+ruhOzRrqO+Nim2q0j/uZpAeqsbMWBXjFzIWozhfiNKz3Nka/ZFSm9Kq
sEAN2a4T8rR97etkjilocoFoguc3oRiWrs/DeL+lsnxbix7IgXY2ojxcrg3uxn3kn9M10hX0x2JH
PJ1IwdquWtxteDo2lLkEWAk2qn6/QE/jVnSSGsMnfnXDJYaSGjYf4A690L950W7Q2X8reAZQsNLr
+lzUsJ8S9eGR0Etn1TL2HL/c1VM4+ah1Zf2wh9uTyl8DDld/7h078bfPxqJq30Ukv22TIaLpK+gx
mwmuqON8yxC/Ze4TeeqINRzV95DIw+drfCsLfJHig2oxb4PeNYq22Zx+OT35/KZwlUfHn51h+0I+
i74kB+ffgyExa74sBwz+ouYKRsp45n3JXyn+NtqlTPn9msWQSZrMeZHtkSLvCni9wxb18u+6HHzu
PCMyeeylg0/kBjU8RVcMqRgOMJ4K4I6nq/WXRdSN+kXNTFcBXHp20PlrwWUET7BZ6P+azp1S2YCc
dOcErmV6E1ee3MyMKZ0rwTGRFzKQA/ijbRZ/To3NieOx7Sh5of+U7cgacRI3f8C3fq+Iy6f7cP9n
2AG25gi2wYcNuSniWZVuVTb2yZPvQIJW6AUyEe11vjLwu0RmdBDM+anQ7ylD2KbDvmosYV9QY73/
9VCbabv5P+dqf5efGWddr3vmLONFltHQzukR+5JvTNVOT5TjitIr/BxvndMDu3NbvfQL7Ff8YJVx
RDHcjKZCIAaMkZXt2yOTuRgfhbJkLsx/uUZGy/tOkOAWp9mmkq0LUofinBiEmuR+OseZt5DF0TQO
vGhI0ayKZCzMS/vW12oNDqf4sRb9xy+8PQ+PMTo3ULk0RntSs/izKKXtJduF+QbB0vku9l9Lwho7
+VTLV06tjF9ok7b3b6Wkbahf1fdcrrECsBvvvpxBRd3WSayt8Fl7i5gf3M7Kdow1gZcpfjIaKyzJ
P/XLJeVUssqpyiTw4AXetfbbiBl/hFeTOL1m8aXeAGTN9a/Z5R0amymh2e+kW7v2rlSOE6yEF5BX
1MSQZflkrcl3pvvsgb8w/StEB2qk0JV2hDcbVjK3ABuPsHJ96McntBqcfWenV/NjrOQB/eE6NsmD
8YtiM+tMRFy6/MeVlRW3Fpk8N2m+t84IHh6fSyzNijKh/vHn6yNJyH+YmvoVEuFDN662iZVYznQ3
SlT/KAPMhGn/BBmP4HDrp4jGk94RX9H8slU7EM73KFTI+8nVP8SbLVu5IiMnVQfGElAgU+wHQJy2
AncL1BbHtnvNPGzs9laQFtXYnUIx/4fuGbNjykEbGoocHAyeOKawjwuuOm7jk/Lvjdn4gHMbZzdr
y8JjsBmH7c0VeZ2PuVhGk6SGXQeLZXFbOuDvKs9RNt96PECTq0y6oAoa6rMwiL3D5ruaqX7wT8Na
9LBdMZzXP2ScFMvpddEZjBRC2sZ3ZshcSjHv25M0KSRPJGw9myrUbdpChibxDVfu1LaO8ab/dabG
QpL7DRnDIx1UQvQMZ4akqCoPFdPk4dOvFMhVcN7UdO7lEbjDRV5oJZ1hwb2uveTMOrvg/XpGhX6B
D6aooJ+FVLOJQ9/ULb0mAAacRAl2DwyOLE7F/MdGffRmDxS87NQ748q/D8sBOGFyE6rsTBuvlNAt
10GLwQqaIqGR9MDGM2ej5UAoT+3rjiK7xfN/jhP8FNPZhhtrUFnMvSASO66UO27n1jCtK6l9k+qL
T2TSwvS51fViKkrEF4zyZUjGynwfOVyKsell4T1LDELHih8Viy/Gzn/v8wDecgRxN1sAnmvkrtq+
sEo/XBWWFnIyDjLq0opzd3I5H89WkkcJXpi4vgncmrEYtpypPgI7s/+93z72WFLaXvu9xaZ06F+3
ctkq5N+yREp8gOZfDJvaknEqC3Pnsk8c2J44A+Yy2XK8gwaWPiRMgzbJRc0kKO6zkhJmuTDZxhfd
ZisxEeU2byXmRgr6FZ5lHkJo973GtwEHL8rpZO4DvYSI/7GIkULtM4LYU40IGDQbrM34PPazx98A
yWysXPuzMmveQdjkPgaTXple0sr29skB4IIEZBvfBwr2px1Q6FIm9hnQyjelY3Yg9i87cFz8oVLi
XEdGVkhlIagWNxKafxGD49/Efz5EdaC9Z8nMFG5FXBx70XGHhAv8IxoaHjqc7qLn+JTYcvXntKkF
3hC6JMoEe2sKAPbu2Vv1CBMBErNzqWPb2lYf03FbI1UfeUFyuMzOFImSPBmOaOAAWLOxlPUbTeub
8gpMAaBDPlRLWXgOTNymF45xFDKDUXOkEWOuDxvP4N4h2oybjyIN7OqUdneTnsBuBXZ6MePwzhjJ
eZBfet3xDjqZS56OSspIAaxvaYNGgSXYUkzT4Mph5eJZn4VlReYWWEtOszd6Qph9ifOj8r1Ts0RI
EiIHwaXYCLQYIfJr7mbsJZlovcjoLDvt/Sx3CC3nrcAjRq4U8kyhq1/lO3yVsiwmS8SMb1hkgRtc
W192FOPeFYo0sQxp1fNrYk2EopA8wy3OuR0O5qtLJ/wpPXV6oeSYHGWZYNlZKQhmqAo/nXZRsjwf
wr/u/mICn7nZ/Sy4O3GB5Kbjmpa9CWS0cTKN+jeg5Ivlnh8FDmuyfrOLJxbSvtcnjVp/QEahwaNe
/Kifq10xVhGJR737xh6+Pq65xwtdykVqzLrfKCv72nAxdVYTcBmtFuGCRUHZCml31yQF4yn7L5cK
qN/9fBuPd7Xr3lMhu7QW0QqlbZaAzFFGR07LK0mp6an2KzmwHkVTPTBzOixkR6vYn8MuhlMUsUmI
NYK5L2wBcIz+C6D3NA5nlNt6sRuqJn/7AfFZ6tCDOhoHlftNtGzxEFcWpVf1RE2MThL4p58rQxkB
n3KgvocP3510/SU7WU0lRqQPmgVRMlVFgrCBKjrzAIpPLC4fUQi+86DDl+xLd8hI/YW9x59rywFM
R2KCFLV7jWaB3KLHNqm5TWO+NUGJc/37H5W2JYF0ARFOQTaGzTE62HeqpldBDmlloDO943+VnjBV
PUtMNv3rluLQvQrPXrKq6xMmmH46ejsYBMyxrVwWH+GT51YoIMmXmJLu8JRljeZ+OxBvh61Ojctq
usFTQesSLPizpTQ0aNDIuyohzrpYYj32EHIgtbkU5EGWWyAFKfz5jOlamOrDxTXPAJGFaLMby0xX
0mb6Nq56/B/H9X/YDyZDEUbCMZ3U7o6RkUN8Q/v7ifxVBb7Htdr733zL5ElUoafirQ2o3lYJ9z0Y
sz+D0uMa3YGaBbdIrN8Kl33QGFxGvR7AmG2lhyE3VQAZ5pMfuRLnPTA/9MfFYQu97X4HPIDSxMvs
fCS1fkmQCa6siBcyCTlUdR856W3GGdDOUMKp51GlcRCCBUo2rRP1VKGWg9Ae0Rwo3lROpNp4m8Fj
5mqTXt8rvdTBDKCeED04neqdaEYnFAECfceDgmjCoev2MrA5W8vEUSgIKRohiqTC76bC0tIEKqGN
JC+A7E9O1jWE/qr8Wdu5Z0KQbnkqVhEOJFcpB3bbOgR3Cv80dIgz7hics7ctRoMU00l0fLS45dCp
FXTgX3uQBQ2kI5tNZW8VcGBm9BwdqZjABj96+JGoItTwWDs5rwhcK0yFD3v+25/ftxtd2ixJCI6L
qtcrBBe3tu9473maAjLN1lQRUFcunYucwcFCn+inyQsQ8KxvuAfjKqO6XlZfQEmklwjHzGnEKiEE
jF4J+md2tngJ3M/ooEIS0EgLNTuyPfwIq0MDKz4CeehjrYacAjzUidTJsq7uP8Rh14fjj5Ti9r0e
95KxPYxfkDGTztbmo4hSax5K/k71TEQxDNNL9FpS7HltzZytnDi6/1bRJnrdMRYmyRWRP2YMrHxZ
0WiBfIUoDkkWBhQt8rwXu38rHS8ctgyyrAQ0/53hU8llGnpUUqNBV6grkyCVKTCcls+WPjc0V/sg
OO+0DAiqLyNNmqXPBlJ6NjtiiQTra2jDuo5xxcpUG1zZ1nmOuQchc5tNvMEkzGETP2cBfz33QaBX
3lEYnk7FnvpQZBa7cs2JLJ2pxzPOsEpUjOwn732vaf8dBilE1ASLklQbkU6JQ09bndd5scjvXG2l
NuQjj6xrtOXg+/sngsYiEBmyvLYyzPQr6yV/ahF/3ptDPmabpLuMZamiv9uweIMaze/U3qqB9BTy
NZjVfUevJrMeaxk2s2S3oRZvNMdgmmpJgAGhtp9XjFVfmin04Abe30Ijp39dL+KsnQkAliEhYb2c
wu3/SCkS+N1u9aC0Bu/pZp+R82TkthagsiJK90zh9rK3+jlEyg1L/rCAlR2fwG/wEVS+p1KG1/u1
1y63OyKzf9R+YbbudIXeO8jdPCKvuaPxrCml5UcoE8SoDsrVHvUfPzxOTu1GZVtv8fz8MphSLwwr
xLGzfl3u+i+fYJF8B1i1rvot/uy6ZEbUO+Skr6X+TfDsFoQlWtw+KC1l45WnFfa99TB9FfwStAij
uISlgdlC1j+mekVJxni+CjjlhJGlJBg9DzdZUypQrAEoOIWDSxQh1FfPl39+9waT13988F8iQgV3
PHN7PXKMw6j7JXNcL30GgEApcrf4DVuwPu/iXUaQjV0XCJNY+RHvE+fbgyOvlvbsJfMx0IgEdCpJ
sKIi440JGZ646x15T/YRahyNwsiWbjudJK/31ebBAcgE4hHlyrFwIp/c25l2+y7+WR7iDGoNKd+V
ZXrIzcl5YldFlgsO09Mi8gIjpEOHr1WcbSD04scl3EIXGm2i38SGxew6DeIvyY61qpO5SCkqW/Bf
OCbIfOkb5Kan/T5r+ViGzV5D7ohEkBqluWd04NRjPVnf4av0MxNFciFt7IguHh3lfkUqrwZ38ven
trag8+4pvER+HOb+0k00jKlwwKfcWnSaEubCymfhYvC0ZjDLZ2/C0JN5RgtnAn2llBuVdwgBS+9Y
vXyYEQCMCPQAHgfoQ8uDrS/GdXSmkna/46o385li4sd6qd2DESRbyU1F7FjxVAHjpbw6wVAqJNzR
RuACLWLYN5RvX0/5HpNNHQTVIkH3izMAhOsZwTAwACSnnVFUl+keTKZsiyeCk/NbeiJygkcZU1VP
4XMGdTpXFPsmnfNQZ2JX2rx2i+VMvDJx33bgJSDSP9xq6GCKzZSUAM1bnODqirUhQ/WxrA+bcQ6N
b48aImwwucLi3q1ab/22mS8AGoOB+sux+KwfRmZuOqirT0oHoLyZQ6cNlw9X94Az3RfV6VxmtY5L
uA67PZExt37OU7+6h/i/WVJl5fNerTSjEH56MPfdTrCmJo5/iQ/RfWV4ksXQLv69rBXbXDZ6MnZE
+67gMv3O19xeW40DAn8g0pXABg/+geHgwjHX5X7URznSNQO1M4kSPpSnAOE5D4dbzSjnL+G6ahER
uhBjmmv8tRrDKJVROjPL+LxSVyo0OoIFZoLC430YQsPM9UG2OURLUeI0a7ESTbF1HHH55W9Jkw25
EEpMKwQZSu11WLYFTcbhqTIh2rljEGiAdZcVVZi/xeMEduqR/pfggHIMnqMCtIBU27Q7W1Z3QfSB
B8LP8Q4EboBFqjwLVO6u3mUvpUXdJhfQdNkLSP14FxbJx/D67Uzz1kMHukL/ULhK4Gg+kV0RCDW7
E6i3eWEkuS9Y6xjw4zfFbobDQo5eFY4+O4wRVv54bjVRWahGL7606ihlf9/Dihe+MFAGKiw6feaH
AI/o9N1Ix3H91wOks8+JZSnlmCv8eQ9kWrRg8Bc9G6Uv2q6t9MJ7h/4ZnFiuiHPyFpJ5ym6d8oe9
WHN/It+r3uxHpwk3HhPvWJHQYyq5vuB9wSGqAbZ0b6I15BfEX9DVi3rBjEC3FaKjCgyF++MorgTv
+wozeVbj52qqoEMD8BiFjhkdv+g00PXiGiB+nk16GQRvXy+e2x19y2HwTA49bpWiePASwsR19JuX
K99t9EIwb6oRHOQVSUo8avUO78skhuSJnuyVtj6ULbMx/Pn+hd9mY/U2DR42p7CLwIvS0hiCYQ2+
EDIlGOunMIMWfCWyyjqUEolcAtNpF64UON+C+JEoYQN+1hMu+plybUJNPZCB/cM4RXMMOvGpBFma
WaPs3rFboMtXBodv6kN8V85U2OcnJedf3excZIXuX6wI8yPI6iAwXMEuqnEishPyM70bquX2P1UQ
b6JRLtCjoR0+EIp9WdzJ0f9fekUjKl3/5QhnjVfv2yBaRBoYvKR3uI3/lqi3gTRyhCU4qeYWfGNJ
tQEAyDe7+vZv3rtaC0jUU8r7ydBfboN252CCUxebqS6b11SowuSw0uUCfxOx3Bv9sSYfbxX2FkUW
Od4D0+rTOM+2rdGGgz1CrrPHkPoKHP6xZyStRkXIFweLfKWVMpVJpB/h1ld3qQniO+Jqsaa/vXnk
wTVhNjdQsIZfwee/65f9ZtQ8RsTsWV7HZc7Rx6eYUFg0BYiyh+apqih0U6kMyc0FiV1xjaBccOYe
RpsHc5n3W1N7c1Nt+Is8DIlMRAA5qS0HlOv0L9VWgv397rWEu4b4Ex2zCRox1yw/NJQH3G9iQlaJ
VtgAw3VibpSK9dT+G4imo0TEYWDc+WBcVJhcjyS9HJ3znNGVQ+eHxV9lFJD4mmOdDI3UOLF0bPUI
G9WimtJnn/gGh4q/6uIOa4hoE75Vbz8rsP9/lG9P410L0qaFLDk62QT+jpmRoLh0/TrD4TArIy7y
RYvV4DPcxxiudhYzfRHm7hCtp+rP6aOBhfxCrPcbUykOV4aq+d/jcsXiieF9jb/8cJyOWWKCwaZI
iBzkYUXGf6AtUPXg+qi5Wa5CQUW/wGd1k4ImaotLiixiNiZZZIO3W9J74aXk0w808cyAZ2bki23r
VxaLno1VYAc8jTZyvCodlGF/m+9SytBE/RpNaSHWRU/8BlrgdOvWLd7GK9/fi5sAmobNncRs8HRN
HBXBjr8mQXi4awDNE31x9pKP4l5CQDRPB1hj5z1MKi3O0w1aEtvlnewkVHndwTyJMV9ycpl4GoEf
dehaB1ASS3ummpoVZAyul5Pzhupo1nfMsCUMAf5UAl+7Xpv0BnEtkJgZUAHWR/9nrRk8Qhik/Vj2
S6nflpCZcDRgRAjWUhn8ruoOv86NRd/X1CqjpT6cTKop2t6ls4h27le0yW0MT+YNFwovVP3FrznY
sOLl46g9VCUqLtXfBaewc2WRBjNfJa6+u743fxJbrRG+OiLOga2GHW/NbW9pUZ/j14S/5Zdc/s79
jyCnAJfqrIppoIkwYfpVfLl0iTwQJJGrUlnU+8mRPH01p3MoK2GC4nxSfzzxxgCupVd0w7J/5Ia/
aRFK5mZYINgFL3zTTF7MJMjGrCAgFt/W0AfK7avY8S6erKqdpnJzp1zS/RJnunzB0h/nlYxwIfyt
EG8o1rR5+ZaJjpmO/xyIEnqbqGzarc7M0Xp7cy8a7ueWgaiCkK/Gl3RDzvsQ+bsuW1nVr758Z0xV
Y6VfCJ7eheV2rvCu26WAhONIALKBH5TgEI/9f22yv+Vj+vuSiOnY3mIIkJsNPMqyd5BSOWjA6Q5M
oTs4RGrqJQlm6Knb64n9VyL1FDiS1eHMjm0DK72EPpg2lZIufZF89UER6XOVl4bmQE/KRsI9qN2B
ZkhsT2GTbfR+IMR1t54FMJ2mVWawzODFnIQZ+MtHRTKBpWVmh5Ls6Tb91miTqdY/P1HCE0qsKZxo
mpt+bMptxhK9LpnFD43A+VrWI7elfmj5uFiqJlOU4nLRdD8CEu6taBs9zUAADjuCXVAX/jVxxepC
wFNiDnmb9GF3cQ/a+Hz1CqJxsMjtdOuNRyHtZP+59aWb1yIbvE8BshbpOn74VopCtQiiJO8n/mK4
zpuCMGEJZDuRM8zS6gX0meQqcnoe2y62MZVxT+t3lPLh9gkAcKcE8HMD15W2GxqppRwiIO2tVqSd
ek7DuQQDgyDowBNup4nxlwMOEw6LDwJ/fKvlpQT50sXwOtAlRwcEAErMO/co24UOPo/0Q27huErD
JhqkZYV+1S8rWhwdgZFzZC0zx9Wl3v76cW+jRNR1f0GysRJgQTxmhGXQQoRt1awQCdricCQIGjdn
5j7lSH0AfhxN4gdU8POEG9VHAVh7+8u2ne8XAS6WT89Xfc9EC4Gnjy/Uob+b5i7111qK81r7b/63
HrAWcrg420TBIsnsQIE4cutmcWbzbTz/o6xSSiryzV21ASDQzwxW+iPTV1qNDm8qrAQZbQ6cHTzX
vAqbk+43FDO8E8j3JPuWLUIa2tjSwHrUeR0CTTOfUj1wpRl5ZZhyTvmP+2rib5J1u+Yct4RmqsOW
P3xfLo6ffVw8XF0LiW/gx3PUvMYarB9aOeXomXqUnhWxmJFByUKXzHyD2QyxEHsfXS3+MA0XCZUW
XjrIJEd8Z0KNpPEEdjVhaayXe+Ghvt9+3M40snrcQaYme1yZn8zL01V7ThhpjxLlVfeOYMwuqcut
Vul/9T9hK7Vg0LO2Ekz9YweNArFpKLJ5gnnZJorWI9Olq1xCywqCUH3NRcMOV+GBNSLrafrxO2HV
mTgBbQiQdLXfwBldwiAVsz7Fn1tF1CJiDlPh82+SHI0xTLAy01wNUklWDXolx0UOxg4APb5d3XcR
nXjiKCOcDrg4EFGDxoessBhYaasyodgDN3eViZTs4Mh0PINP8on3PEE2auFS+/iH5LbQ/1MAC98C
wiPDdvpp7zYijQWcM/ttFoanX5HxphoXL+V83/mj0RSc3BbHe7hGs2MrOynQ+/GoZyuMTfVrHZv+
Y50ugkcpmR6fMvq4aIZVI4Zciz/JFtr5vE1Pa+aUn++5EPGkSK6PQa9ZijpGZrMRY4M3KUWB9DuR
MXfFGsgE1jhS+INLcXc+mlK2t/xDSRJ/NbF3RLkfqFHtxgV9575MfOa8m4cW4/uxT3WqPifrWnXd
x0ouAwU9t/t8tCeDzAyEUDRk6lTcF4jJDCQU1FNH3V7FefLKsPiOl83XZVphd7SUhZ52M8VMzXCW
2ttsRXUrqAwLa50kgv5kTJS6ok80/INIvpmJLGQqwKqnqi/4GvhAXsoI5IRm+kBLzocPfMVOtTGW
GqDsr2YCYKJTOqO7ApC9beZqli9KJv32ihdxNJNcb8N6PxIacP2BIujzgrzpjrzdF8DK71b0ntZc
grGY4VnR3mU5+SFyd2wR1xWKDpD1GetahapfOlzAbZRgtEBHWWLsPPk75ubO1dm7r3aLaj42X+8s
WUp3pxftY02VG/VLjyOp1wS65AhEONBjiXjEnSGq0LZemQo1IBsFZx4YagcWrSOomKUAnd4O7/mi
UP90+byTBscXuEMS0ZeDE/9Jqa6mEqWtRh84KCa37BMMY0vbWEFbLo6xud2kvhlL+8zct3CktC+h
3irPnGOlOK1EAqOe1edgqyJ+Pd9dCc4UtKac0nrOYnbtheDS2jxMkd4g/14dwzRyK/r/WXiqkZHE
bzGjRCu6gz6/Pc7ryGNHfqW32Mc7ccuggUsDGiTwMuNXOzjsAS0ReFoP0vSUtMiuJtkhlrvXAMRG
P58Cyglt6I87xuFYLzSc0Q7T6hbr2n9ddE0wFQ0dtKUP8yeRT3OyVTSwVdM67BKAqeLj3Kd1CZCA
wAO4TAkBBUx40q9m0OusQM+DTXf1GXdH+QLc/VkyCrYtc/Uj354H9L0GD6nbW12X191xUGHjl+uG
Vr8wD2Qn5jb28cA9GLUGl8rX7ZMcnEh/gaghznkGF8isZKHdkEMKtg75rndtCkVVpxUa6Mvxqnkf
i4idf+B23a6AWv3lwg5FHfKOXA9YlOl8QTFRCk6xu5GmFwR79fJJg2kGJv5lBQg0TS4VsOuuiJjS
oUd+19/QgX3Cq629FIB/LokVr5u5Q5KmQbasrFt7MR4nsdaDimMq8FS72/YwhC9+bx+p1ziLR744
OtaqG0HeI3dQ3ky1hVKasYbCKTa/JxTG1/myxCnaPJ71jMwG0znqkj300MxQtwC3ls7AzIBMLalB
JIdDntuc3zf1GpOKP89EAAYULlKMrd1djsAbPfILJ0cWvInnrVHksRb2sGGVN8rE+mNWDxwIpOlJ
1tRJb1c8uKEl4yHauPjQI9WlYNqjpUA3SxgTBq3sx0xIdYDiM4ReAp530DNlmyo0ro/0Q8Luj6kw
62jnT6EHnMkOKMGBL81ZwySmLV6c9uXVKKhfIPBR2+B3VW9aEht3RXje9JLJL2rS/2QyLFqSdY+H
TfyFXue93I3rH+++sbC5Q14k587vBOQBz8t8HX19GGdd3fbGUz4vBtaBqH50BUaurwaKUxnQpRNw
Jv+Mf9H0qP7/SQqH0VLm5qz9XpDlxm7H1EghmFD18T1aRtujUDioyxl0EJzjCQ8xZ86Vg2WFXAMS
/62WkNdcFotIw5ngcFZrFH3D/wT5jMyrSsW/k2p+7xa4Akh8spl6IXmgbdXTryIoskE3tKZHISB1
naS4t+HyyiXkkwRavkYuTmNfvNKlGgTSWsCXlmUT5RsO1C6TQcYZ456skLt0esTt/6b2hrgj/cOH
Jpu1bCLXCMV1tJzkLeWVh/FEN+Ff8pYp8Bp6fzczgPs3gtjCBumYF3X2/rJoP6qPptt/GrOPk2Vy
D2xMnKiwQYfAXyc2AK1HfrzY2Gj/gG9a1BQsEGGSfkvPZRV/nL6KvWIrCAwxRRZC6n8Z2mFcKVWT
bIrXLeYas6nVfiqqHr/GzUqh1PrIXi5URJ2bFMZPR6ZjZcOnp59Jw3hoNyv9EowykXOmdvlpD2/Y
8i+oYa+tfP6Mj5dxcqWmEvg93b1eszxkgmNjjxjWEmiR5RA8FMdERrq7d97BodHS6uqqo9EebjdK
+7aSXORxp8Kct3xFwj9DrWltQFfFknq3NlnX0gdXwyZU6DWRps3LY5XbUDDO+H3EOFFt1G3/amhF
eL/nt5Rhtpfm+wp/wAhcaDnybyUuc8f2UQnE/v2g/PlYMhDiKMTUsGZlmg/LObynl9Xu0yU4JLHs
BJncXFRvXPGMJf+FyTSKlwNLADtly8WaTrkT2uc1+IitY5/zPYIKUcr2WgxOsDn83T9F8MLts1+O
j55XLJ0D5jh39+0RulOcU/CfgYf00KoX5rzxecn1xVOlhmwUeILA2SZfIGt3Xvao9k8ITqcdKK6c
pQqxSYoxjPZFtlkQ9iPnGcpbZo+stoEqG6eNJzTYYyv0pz99FGn62YKcoG4GKxwSF+HksaOgLTva
fWBEcezvOspsVqYcIvYCMg+z7ghyeBSDNOOeMjbn4H8/XBjrcb01U0qsa2/JqTTcj5U8aZH0OTgV
Pd7Z8jsG04MHnO/WOuc+l5sTZSOkO+QDy2FUS7sSi1zT1Zu19ot23BuMTR6snhcrOYcj32DyWfWi
IoPFpnzxI3fAMF2E8G0MXOpLN9uRMR7Y9meKDdBJApWt5uW7GhrOIqtSX6GJpzjAZGOSNcEg/bH2
s8YUViLbntoz890wMbAokCIIIvt5MIRGnmsAGoqQvdVWRevMErp5wBtUifHbAB1/LZajQseTrHe7
LAc5tjZSmv4VwPdKFIahhGIH8s4rbX98VFNxMpViGha82zyE32WSCYLxgUw4IJ8NZJiJqorsrxbQ
whB3ubSZ3xtT9qIFet/dzfpNJYdHy9v/yUi17xjiSgcMjCZYpjmVbA36MOgdw5Yeh+n3u76pfkPI
8dSSpAPAslqdEEkWelMo3CyD1DOJLfSAAh9fyhdz36Yc3MN/TdRvp8OqACIzPSnYO+UQ4qHsCjKK
2rilrvwLXHDTfzUJ8pOL4dbVAZktv2mryVXdz6UfqI1xTv9vJBsX/iyIHW091ImunC9Sucq6D72B
X8SfsFjdpWFjkOtiGR/9a0mDiz1L0Rg4QZk2IJ981K48FKyL0hZHmTJ/SUqT9LGna5tROybdz778
ltyHrHiVoPb7FvUfpbFClm1idtHstoTzGuyRLmV/BjxHNMdVEHbwdzJy9TGwP/LH0d780+s4k7p3
qH5ecOTAYCSP8z86I67sQRrDuOSoEMPK1tGcXpsZ4Z0NcwZm/zVjduOEy8MfWioCJE0VydECx5f+
GYRIHC5a4FM3Zd2MZxofBXaN4HAAPivKJdZBBJKsJLKLuSPR+q+kMELTUSZAqitwNau3eTwXrZvS
uZ2sciTiMrYnj+y5NZfI7Bku/tFtVJPbHHDRjJTFPMURmNhxFxAMscOPi8TrTjRjY+93RxWQ91of
PUXJaBLRS8KjuEVf19SOaFL5IIIXTFTpBGcRUzOib9gK+wJw0miJue4kcGn7AmXOk43gMLiFHN5r
XPfEASrP13ZD4Uc9aN9BnYMcmzr8iRT5oe6/ViEc7E0SvW57GUuvSxRL2lqJZ5mbwmpffweWeFlq
eykG6cL4vw5NET83Hedow7qio7S3yiZr+DUKD4dVLUfekMN+gF4nnFGUoVYgnKx3zrWrJ7PJeHMy
IH/bJCwgVId7mfmvw95c0Qv/RI7saKJMSZ/VkL9qDklzWjI6oq3EuBfRzWa2YALxg8c2I314qQgQ
FQOvcq7dz3akPrRoD0qknNAZTNhEFkU56l84D5xdTuEu1k4d0W/bFRc1XSR5prneAsPnGD955BRe
uaT5kHWccxTjrD+UG911MiXpL0iBSwem4rVD6UdpeJ6zx2Jkyweax/qFI1G9Ov9y/NHIKS2zbtiL
ggp2a/PDRb1xGy7iashN7JzIc+9E0fQQt/MkfVTyz1K80N3p6MkNSaaAEhyGI/acDVkoEKSpbWwX
DKd/CB8/gggcUesU1omTLqReZcaJ0eDLmhhamCIunrbrzqPuU9dnfcHS+57fhfbHVw6o3ViPAsTC
7mwMdFg52dMIKGYAR66gZijXZq8jnCYD4K9+koc5C9MIaaqpanUOr5hKCWoxiKlRtceOUfqoI+Rb
PIri6Yn1Xq53kvMuUuuQ0WNB7D3cbcm5qW3wovOJkeWafP70zz10SQ8B8hGlW4cDpj4/+nWixoIm
JNAAKF8kwVecG6tKboZqfD7heAKChWFUMKmTsPgijkfJWw0ryVgy0CJJ0D+tTUXyTk153gOYLji+
8G55MTp4/PvCKriNIwpc6vhjisgP1S3PMsoJ0A0lQYnDF4xjngBjsES8Ty7ctCS72C6OAJY8cYGi
Tnn9yHHm8fFNC3u/jXmMQdV6TawCCkGN2v2Et8zd93nv0Ib5jJHGs7PqHMp/gQNS1GRHZLyjaFfb
PUQ/jRRqLirecTNzg/2bJa15fdbDXb8zIWX0O4LhDU7+xb8bwr45tlVZU3zrN8FPWP6B33tj6SOE
yi1SlOV0UjIfkvud8OYA2ZpammwiAz/bj3n6hidzLNwrqBTnpJ2gqAYZSvPF4xRAVhG4NUKIG6nN
6lVPRVjQQniACX8Mzg4MIVo0HpOcaLGFgtWHQgl316hj3M3TrRdAIdw4mVm1nA2S+JcunAMxqim2
VyGHhSkgtN1vxvV4awxuxf6I+cusBw0VTVgoC577LnSpIhMr4pUBqHmkqNdZ60o77It3C/WfM1n1
BO2Nv8JYsOXkCMTixuP1d+XRoEeIdgrF/C0jZ8h3B5YTL63ks7wh4R1Zzx3E1cMWUQeA8NMsMnc6
c4asTy0u75zrtrzmALul0R3MdprKFLIN8e0+4fgiavjvofPRelzN6epsU+D3VmJn74sXxnxt/y8D
oRl6SEsES3RroOTJtqnwOfow6XTLhJZY0+KR8UbVtqaVEATUDcOEgFIUI7j2Q/2TXqbUgrnRXZ7N
yXhPE2a+5FCZt4aBOfKPa++uYGtmlEpyTglbeHleMChjV7OYB4uOdxYl2IB0uFw2UvPX5N7FUw6t
MnUe/RFf3qxoSv28i39OSzNs3914oLsWTIvNSvVIsCJ4547OTp8DN6saZiAqJ2Fyd8x+pZumGWp6
4VFI4vjzP7J851QMUTRxlUl5UlGlkG3NREdrEJf6rPMflqgjThjdOv6hXbhivUEo1mt6tuPSVeoA
rYNHE083zhfCXLSnUY/p/CxkcgWfKjs7T8lRR632h3FV+LwRH7w/tzcNunnMrXxtAfR3Fg18De9D
K3dS17MQkodLBZr/yeXjf1to+vli6BRBlkDEu2SMpcIQOdPetfZaHtGVTndsU3CDyXMSdWV2PF3e
rz/48Ss2R9Dy7XHXf1vsaF3JkI7gel4IaaVk3noLPuMYpYh7+jIdEnen6D2hqV/4aPtZhWOhsTHi
NsuT62iPse9CMf5hpUrhPM8MO6AnDQaB/VCgPYaXMSxj3UIy/t3Np0kI1KqbgiuAFkc98Pkp9Msn
56jIYcKy09nSy0wa8nA4B3HcTFP4y26M5FFfXyQFl1UAsUMrhytnkQiqoJCnpDQgEfDciAS2JibH
3fOhTP+xOQOkgPD+K6DgN+lI8mHtF8tIVfsfb9IBFhgjlhGPtzAiKyH4KF6pUDRBE9BPav4gOnwv
jHmjXo4+Xma7FK8BaUWGoqdsZIkUxFGWJdighy6fcP+5F2y7Gpwswrz2K9q+YMRNK3ZPpl+6xm1Q
6YRkAR9u/k2V9uGJvwcxn8/XLIos/sOu2xIAl8n8sp1lSmjofy+eYVaqli0C3FOzcOZzwsl7N4Dl
RxHowB9wbgC7oGKxYmatYZBdf97LuCOs/xZxeAjC0zSXDojoZIJvnDQFQduRHFueD757ih5pgiWK
aDB6GqbEQQZfYybRRfVWmWIKiaNy/TN9UE7SP6ShzQ6MZlGZAUyeobqmxKuqqdHEHrXuUDooCpGE
T/S2g7SQM/4/ze4n9L0PTqr3O/shCsgKJiJSgP9fZm5ujWSFRrMewc4q9sa13xAEup245q+tvE7i
6xbovrWwWu1w7dOkpoPoBxS5wJn0DusgPVPeYbadNTeuQuBIVKuAc3VUZQmKLLf6kDJuaeFqONQS
6uT3KXMmi43Ex0bRiYvewUGt1cmd6qdHlfQEKpi4skp7fJTDAsXblwAPmCmAb9rQjv1Y3xbDjGtQ
Wi73c7fi066ftug6ehx2FbIwk9n7a6cA9UXEERYsbWP7btpyDcu6uQbywqNbakXoY1MrWMC6bRB6
OeGv1rTtCB2nWDrkFbuD+mZM8IQlSwPFvJ5S/Nx8kwhBzwWDlHjKJwOlXXZwRg22N2UsgRsNx59K
RIscquZjzuJRDe4P6uIjVyYC+m4h+F+GVAT4McDI08HP3TzQ5caE7cXpEefRj94d0Ao9t4J+ZTYB
SDt00ukRcT92B6k5z9jaUbFA0m8l1JfwvekELXJsHKVtXuhO/Gp7D/ykgpgiwYBfKqXj7rwDB9CR
t2Wvq0CtYzQFi4m2qgFPIyJ3Falzk06y1bHVEi1TxUJm7jGnycLKDXOvRA1Zd/tiIJgd4yL1wcan
5MRl8M7DeKYc6nMPSGMN61Hj4J4Nb9wegF1k12mIIYrb+jOo5VcFjG5Zs8N+UrHaTF9l1X/QnGkn
FQoDekK2x+bPA9xUtho7RBNJWB4pF2JvjGLcmiHeTO/xK849L5u9QCRRsfJHeGgs0u/P8uXZSopG
dTBIVj+S+/Fde245chq4zKr+zlTPvzjpsZluglosDZMnFwHGnBoYmMYt1viNQHE8BqcL0WwPqrfv
HSD1licNLAFTT0rviIAcHQm8fCWFvoXap3K0KiAa1z5X/3TzdNFGxymL8GXZH1P4taM+A9k+hFXR
IheZIDXtNu6+VMWMb6ff1pFXd5AkbtijOKJsLmqyPWeUjvSXuzyOout6MLiUIXa41DtBI9OmyXNI
mbpX8ulQM78K0pLiL/40EpUF3M1ViO/eg+OJ4WpibWG44yVyrq9vZ2pOvljIuzjHq4c3gzYPisGM
rMOM6F+CHk7hlJbks6gbDnF83+trGlRMiD9U9pPo5uY6egGnNz6VH4cfkf9+rFKRVpYJlPOLJX9b
k+XemdYo9gFx4KJ8yWZlcns7UPr39nsRL8iUHH0lZpqwHOIwY8Yu4TiDBF7pRhff/Yo5FiIfpwLx
ZX+/g+PDNpl69pytBZmCCGTVMY57ESN17QIKyStSQj/f3o+nRQ+1I7dLy+jtrgJlt73Kupui8z/3
ZDH1S9SVrbnZjBbO6LF1CfA0ZBddF3+3QPU5vxHoneFW9KGNKHjOXHgoItXSQsfzd1tISDyw+Lsf
60v9TerLJEmnzGV5j3hQK3H1YrADb3lDe0sFI61QNCUjKo6ETZZF7+iTy3fb6nIWIpXWrdXVI80S
Q2d6oXaxnFxiydPr2HJvQjiRg77Mf01xEo1aJvuUEIeSxkmT+pBv/VKM7sc14bikCQJPiHFt8KBq
ecxJRcB8M6XCmxIaRldc0KaBDdbRtx53E/jwgSJ86G/pDsBFDXWn0Uk5JpCGwDafam48RwMVUSFn
aYnwm9lqatgaU7LNZU8sog1ov+au8DEIqBYOyc/zjcf5iL+cffw6qLEcXljq8C31dGefwDG1Phmr
oG2YAYWuLBwR3xnWyYJupoSn5G/VG+UKFiItewIyO9eWXBj1tsCdK/neGruNGpHZ2v3j81peA4Pz
I8UGUZu/zkRpUCHZ1MgEzRyYH5IT4CoMOameMmBV4Fxnqi3YmXr3yUnNxLHRK3iLms45yuX0Pyjc
Coww+KX0gApwMUd6uNI0JiHD9PkxJI75HZEiDbvditDHCmpJ8Fb3/vp61uvqUfKM/hlWeSuadUU3
MTmkq1gsveub0iYQ0dciCty22kMT+3lV+FQ2GlIgzZnoUYWdbzqnWWjH+4PikeMunozuJ6CGzCos
PV2Z1KneV3ylQTjiMUNRunpAAW7gWglYHzxdh2hXxhnfLpistPrDtg+L5uhieqClTMA4VggvQKle
oZfKWv52PfmB4WxRImp76WTbxBJm6unNytj9zMQZlH/WqKSSvTER8oI20NdjxHkvfEW/7FoO/z+t
Px/+ZU8bls9BcbREkgtnqDP4CsMRfWIMql+N1nDswlXuUg0kOgBU8ZeZTJ+jGjm2w5s3cNr0Lhtn
uLjg5TDb2UvdI1UCCAtT/pmG7RoRAy1zIRWdJcBFe3xAajIt7W0MvyIyuIyxztXCuEjN7FnYUXR0
hbSnyW3l+1C6OvovgJLBqfk4PcsRtSD4GLquK6ms/L+/h5ePW/6VNzLgykDDZG79bzLq8lck6kVm
avnuE8IsT/hdIGhkWQ12KRMc2Fb4EsqDuODoZlzt1pg409OROTDrdCnxQwmtO5ih4C9p+uI2FJBN
17Yw5tPsEBY8rltags3lJZ2YIqhFvFi/EQZH96mE8W0F94W9s7C4i4IcBnr6ihD1CLg53n39r7R8
uELmZ2JZBM13J0ArQN794olZedmvzIUNNxkkMzHojUYD/pIFT45cXt7lKwdd84Bd4P+jesR/O6Pj
f7dA2mx4iCB1UyYSPDviQDX1Jtgqm76UGbBKE8uQSa42e49XDdX5pSWaAgBxjbC1XPQv1WihG4t9
HHILHEWlRQgxhh/ycW7AB6dJAoZygCF3K0WOFX05dXPjqvWVRkSQOTEkBiFwu9Wd7EJVMhCnlJLw
DKB+vznJHzNfxSnU9hwxTFGsEW+CNQYaoqo9lQaJH/AuDLtt2+sq62OFaVR3NqHyD9zEroo13+w2
mg80OUCaR/l3/13RFYrBc/CGwd8a+Pv7SW3L9ZLiN0og1jLVSLl1E+soNqqW4A4xRjyZ3KAFWgrF
YKnJuhcOh5ioge7Cy1szWU+ynqPKwZgIh5w684Jtwxx9ji4JLdUreQ0nI9/+a3InR3SjjoZYY3Ot
cEWXytqUu8/9lCKCz1eZrQn8Q66Utzd4KwnjyHnIB/mN26je+isq6W5vfQatb8ZfZQ1zeAz6Ke6v
SiHVwsC99JAxP9Anfczh3rJyacxnQwWJsE9QLaScCR9U0xjaz/e8Fh11laULm2thiVA1LAXeBkZQ
GdSO0WDUlpU9N4A1s7LYxEQ8hbUk7kdIdsXm1QfVi9NgXV9kLXRMhIIKJTFER+OfGeEya/neZh9S
gu3wWQrH9d8WI2cz3lnDbXI5wIgnhAI7dZuAv6TrMbKXlYSBvVDzbPbVJ+kpa+FXef6mNmONmXm3
DR77o/KrjiXGUe8NukqMZ91sqHfBFq+Vacys6GU9GHXJRU/MnjTs7GIOeB8lyuurzPi/2iJ2Qs3x
voAz6AKenYgSXhb5QdvDNle+RcMZeznx1fxInAfyb7FwGLduCL3Jium6j0QChQ21zB7a1j2A5XgA
MmbX3f7gDrioUtoXTCGj5+5mRTN5kwYHVqVsp5TbVXwaJL6crC6ZzIoTUjLjRdfQatGFx90Fvv4i
JfV9m+0q7lm8s4FhshqIrAU2tqK0m1V8Bk7ezUxmRiynWIzfLwM83oVM39i79YcnWQSl4igDTDMI
Q+++Jen5Xi9rhFDlUtLLapvWHhHhsQ1RIe7Y5kQUp8MUoPPpWeTxcuWq5YDyA8/BmAZRWRlsLF4W
uUjjkTDwDwdOV47v4hQhz8Gh+ic61uhEeUJ4yLfCNU1q20tAX40KoMACA+ZQHREdj+7LwlsCse9r
Jni43anRkC2QdYsCZrg6DCt1Q1FwWf9i0fuGVsbSK5wwU42gJu5+MgYbhWSVMUfp2diJyi6ya0GN
61ag0i+zNwd639nESgvIMNLGH2WT5SnCfUzDsDT5WFKp0c1rkVUM9x6RHNFyW/flpWrwWjxRBWew
GVItrB7bxydItX/kkaz64qE4rg0mkBApM3V+ort5W27RZbZQaY/WhOGKxQwXkMbRabRpCQwkQ1qq
X2Le0tYGgVdYVkJ/Qp8M2GlBOg+zPmNBo19aUg0TuDIml6MAzot6+EDJd6q+v9BduK3i8sWdANis
K6it9dToUvfMCkZtjWj6IQp868KpTGXDcUPFXvOKmgu2WXmpa99G3i8MD3vC3hKauZM8/SIlJwRR
Y3o+PtDEbSJQbY2KKSUWFj4N1zflc68I+J3ACDLundNVi8EzPBoePENdvW2oRZ0gVNJVeJEqO9h3
Q1dHrDKcyMRRQjG3tHeDy7K1PXhH+N6saBfpdWlJjqB4DrQUmSUbLezmgxqChcwx4BGOifW6WgBG
A2rE6/fJzP8q0oL+z6+JUzcs84KmawqHEk8m2Az4AES7TOKxBgJtJLakx/40n74bN35+Wdf0kNp5
NPr9P3h9GzEYLnrVA1F/6gZ3Oavnb4MLVCm55hH3IZMic+LCbcV7m1TyRp6O5lWZS+a3nFYc49WJ
h4ELDLgIkaqBgExKUuPjlrneRTrUjhhL6OVK5aCR4rKq4y2+GUEviQjEzsRIcCFxJYe6GwToJkab
yUOnulXC0LILklUMjaPWpEkBUmaTWkpZ6DOM5GVLQrlsPr/qTXh9DUv5JiybRARfpVYzwqQh84AS
PQ5XZ2Of3Gbm9w+sNOYPCcS1BJ2/PMHYICXs4jx5uzrlBzY0dv4ALTxYLUIw7g0j/GlibNpS1MsU
Wjxb/f5P+Citf3ukHSfbyLk07jygn0V7F74FQIYbX9/Ua9sQ0l5QnwMsZ5rZBY0YaqXYn3UaBB/o
d1XtkBSA+E2DYxq7yK4++XISo+UsAfGLPqOjHLlQPo0GWBNtxIDfbMetlEthy6ysT9qeZGt7rVS6
XFwskNWZDHqe2VgBZXvqIz6pbTqUgCLPJXtj3NVLQ5n45tSMrRYKoCZBaRkUJkLlyvGAxny4Z5SO
fv+gPEWC03aQkZ6jiuvzw+mzsD6u2zWi2ssfA6VA0+vNdmgevhi2BMc3MiNBF+ega4fT3Pwtp4xC
56YQ3GxHVwXD9ajLwoPBaWXBy3aZCPHGHRZvGHOzRdgKp9BCLL1ILZ5O3pjlnzilodlN7xnx+zCw
ldiFdeNf0FvRVultcxT5IXKpS8+o7CwBaKs6DuCrL4V/V8txCNzE0gfmFJoh96V5nT7AoVtrfN8G
8Y4LN7bGMOgIp1JwZ35KkYCc69ez7iMhmlVDnNMrJ4yQbH690rprSmM3NJfGfvNvSVNTxeHhnUUg
cMPVi3Sx4BS02lEp0wVzMlRJgEsIctDNhd//hDVso46aMkRiL459LtaB36Fe9WqsIblPezluqAEu
fWR+hQFabsIe0N75x4fnorDZKivtYIMBYVN/YNQDa/gwrz1/fDZOe1rs1p1KTa5UXbBm2cJ/+1W6
segYYcCKtEpWoLRkQTz3ijBa93Oh/W6aXRrOXzXDv9K+4yB5s8Vz779NFKifOEuxQp+upSALDorz
VEnBOizAlllcxBLrtTOqkZH6sJCihbp8VTPN4WBH1BOytiexjeG7SnSv+c1QmPaQFwOOLbKk6bm8
49L+V6GDX5oLKK6tckfG/0qVTZsLIxQ/8TpvcKPU5fuuz9Cy6BL3Bsl+o1ex+s7m7YXvLjtmfiYE
56qJqiIGP6IvT/6rICZpbFtzHfD1gtxWKz/T0CEgC/G85/aVpJvkJz7kirwRq1g8RbJYyx3IMJez
8Mo1Qy7SdJ668BfQVB2GlMfB9dye8YjRcb0a0uysyd43/06Ca/iLWtsCDm/QNojLfCf1ENdlxvnU
sve/EMTGi2drPprPlYZ09xqiCPXvJ+wL12pSb3dagfncGIdBraevU6dM/oiBCRa8jfZlz67mOm9n
g6cz6k23QkKd3sAX/6zuGb+SD6N+mdCpy6fNnJK0480NzA4L4G/tFelT9hfzigZjD/Ye+eRaUCJP
aBJjsMHLTceSHmfD8AA7BUdhsXRkAdRHpCL0tfjNqVlEHcb4pCwION1Ly0ZiA9MvgjRPULArSEvE
rl0jc54PE/9xQSp6ImVU5DDsGJUXarcyYM5WiKLviuuyIooKziFWDtj8NejvNczbWO0yefVEnrAW
JSXRqCv2IZLDwUmtUbW9zrhODqZTrRfrPy/bqLv2Lp8bqmFnGvzJYs9WH43Tmdo+Pcec9MIEd3KE
/Iy9OyKwjaZ+g/wIaea6DiO1PhZHTT9+uV2BkTlnwKgLpEr0ZZ5ANdOc7N4ESX62Pkc2or9Z62dh
HZyNm+OE/Sj9mGvtA5faw1DkblEnwmOQukhiRzKGLcFaFXcMSaMq0dGFQXXtQcpNjKQMVOBPKxPN
EGjzCoyb9azT3MJPrOqgzVGa7hsNgNfAXPiNrTEPoBLhX+HieRBMXVrv4fI8Ybqzv/1WahauJswj
86mM1fYWFQlQzkFuo0ULb/a16kIg8FC+f4uOuEC6DJ04yeyvl9ZStLrJNVto8ofVser+K3CNJ3X/
iODdsD5z7Ix6N8PG1/4FXecuU72OXeQUI/VIjLD2Xi4bdmtcxdt0kIUgkCOBF5rZ7ZPMLUUe3/Rn
RtDBx60H/s3da/N/MMv2XWAtxEmihmszu71PzMUVyYAfHtKD0dgQeBo381pcgsZCNYYKCKnEb10p
b9NMqtCUXgJXvN2/kKOasXwdphsPnK+q/bPXF9u93iRbOmzq5XX0favwfQiW61yXU/7SRnG+LAfv
TYAhvo6tN70wIw9Jp5aGy50kbw1qqOK8DoGIglDpEeig75I/JDTxiEU+v+vl1ySIqK1qfNQ/gxae
KC7C/W1HnBixhl+1WzFgAgWcKPRDy0cNJI/z1k+WZ9ynVtnjfBvFG9hXi7zQstv239CqgZFtdWXp
veedddfVw/toBZYmHA7ZLNRDB5ZAqeKDqdAfcIxUiujx2+GSS3U87ozX1Nv8MjvYFd1u2nEffXan
F4A5fhDe0i9fqbVhZRlwIM9eaRRtnRCbzDMDabVxbMGTWRBNFL3mA2jiyXQeg4pzhuvWWiDVsrc0
E29CMKEn99x0Cp1lw5xgNKmPQ5L3nsDChoM1+AJCZj6FlfG2ggvLXQqngFZzv2goLeKEP7xPZv8a
0i+WvX90Q2pi9wepQ1a2H5WUcIlE+P57rRjx5usGU97nZz8Gqn5ikabxKW7tChWAt4egCqFj2ufH
qBTP8UFzQQAau9awTkK2K6Jy3dGFx/kPUnODK08Ssf/BnNnOGwR3zrdZGeXDqh4Z6cSlQNkbG1Ly
f59AaFevIsYc02JRRc7XJNCeGlBrwDGF1f2q0NNrQI3x679mMEjsibQp6Uv0YPEfkHrV2koD5LcX
hAcXpTMUXmyLsIGCapA+kvLn+UyYMsBwcDk6iLCG88Mz/38FGvEzVues15lP3g5cjzFPz9scqPlz
XPDzx2pS7epfEO2VyzCJFv0an/8Dk8sWEQyfhg5w/E5OE43/ISFL2pa/CahWEQiPct217yvipy9Q
UU6aRQWa1ITi8ZSzIIf7QOSm7JO7W2bmmUyaiZ9D5upeQwpFqvudvNIE3yeZzSA6HDwrzBjLS7cQ
fP2YxLhDJC48JBtSp734a7ncUrforNcBGC7/NrtTiu6XL1YYeiv7gfrQk751G7c8FUa1IHVLsWrk
P6Cvn8/T64coTq4jYh5lh7YNehh5GpBJhdvEvAcMLyiUnMxKYVB8EynvyXb4cWj0pmnDiJe3WmNN
f236XGPSYYQN7rD4FPOblT7qU6H40g6UWctBNXESuEsdRN5CIWoDey+x7gBE7jdTKr98lDgEsvCC
TI8APmxdVkK1kN23GEvY1DGur3iT1uhAEcVkz+/WZA6+QJJ0HBFLcSNxr6ADF+N2tuxbpS2OQwJ2
JGmGc/1OHW66S07PqP6HvKf64SQo/VXaPSHyWXDRAaIgpZuLf71ZgGH/zc9rr+S5R1R7RT6K3AH9
jXcTIwih/lqgPBK5otJruHAG2fow0EaPi2rW4cpzyrfQireKPVUCA7GeCHz1s13Sm9cluqV3Gs7z
6fff8rQr78f4AUU/PI+DsR+jjI79bDCGKNe9v2oqDPjeh/HyCTC6fIzEz9esrQIIWMddIKwrOBtr
770Rs+jQuhnm9X7x+EV/+fW+CbLJN6/5x+O08GRc9YcFGQlo7+FF+dtOKkaXuhQug2WELi2DIUNs
Yoiq8iShjA6x/ve3mGCNNdv4HfHo1fTw7pBuResFr2sm2UrohBZM0tNp4Ft/7SR6v8iQB07c8xSn
IJd+GxlzgpiA4vip0WDke2PonJz5+Us/Vr1AG+zVmVrxJCkd7gY0SlRrBCp+hmu2iZV7ygzmRGhN
dt6wp818i8quBSADCNv2IOlInuMZL+K5NLqjd32Njlv2tl87h/4FpdmtnOQ/a6Gs7mJ92E9Wh4xZ
hTpCesbFPaiRpdimpluPNrVxUJx0Vszlqg7hUUH3ZDOMS66wyY57WLqjQZnwphmiOUYdZGNYClmv
RdvnFGDwjobpjxDkiHnTA+NCqqT6d7vBMSkOgPtK/qHUzZdwZ+3aG92Ee1EsbRdteCss6x2MrhYW
/i+lfz8WeRW9eoKVxnC60j0uc7mKaqpQnPNvfe3PvPCJDIcelfZpVeK+vxJ+Z2pIIPxe70uJ28sk
EJE3dWnLMi1ptV1fJNozcSN89eHWfv+ywBD3KBs1SrgvlmVYZtroWhdUMI7THXjcLAbE4qMu6B2h
TbOUk3WCP03pslZPzcWnUxtr+iilXh07g158mYOIU0ugdbYIsG2R6q9bvfyd0+hH8QG8uGtsbjV6
9KN5yZA4vEf8ovBEXLOWlwrOIEQkelKZteOQkRtL9M7rO6RUSTnLbpPF+ybhrlmyAfcYFjG46+xc
JMZBtKoTXJ+odmSb26yJ1S5MdbI4mixiPiaTih7InmzJnFvNispZazemdCD25gwhbMliCHeWl3EO
/5rtR6cWiqh68iChKxY0YyGIOiYb07+FKtHIma0fZDgjakPMyK5bffyul8COvqv8rbzwWBd9odnp
uhggRxoC458CtemX1V2+w8cmmAQAojzh8Ahrz5yxJkUJnmManNLGPwqIGQQ8Budp890uyxSYRwfO
i5MpVBSTvj1MzlrWu/gkV3VW2tPPOHiozKtaD8bYB/HEkRvAYH1DiiUX/17hf+gK69pusUBjLTjx
TbOo5SRXLstlE9bijLFmVqV7D3KyUaw6OUcCUMBfgUmtJ2e1w5MaI9nA6TRsJym/u/u39C+Q09WE
vTq8UAB98aPzyt177t/SYW+8zdCMBVprvdhn6hE/k/PlQAjf7eMfAevYjhFZwodVjCKqdZi0DX2B
t7E7CNjaEGwTnAU63/TTUyIGObN7ohuU+YlHO+HBidCw4JFAApUT/8SEXcjxE+UXslEOffwVGyXM
9vJkK08zLwTcgMDpZ14SfE7JXu/a2YnPai7gHGEvmaP858pDvSycKOsN7epKerIYHe9WSdydIbsR
bmN9Lcei66ZrY75IOyNc7T6/wSP9MT1SAe1iYgk78Kzc372+8inDzVJftqMxvY0T7R2KQRhncChy
VPyy9o1Wjx/YxpoI0Pl6KpYiEDJd9nXkP0QZXVNgDtu5Kx6CX1qecJ19Dx+UixkRe1K3m0mTFB3U
pFAQtEvDq+LdJctPjeStWzDx7hNtf00hbnoFdwTC/5nIjjVKxh6H+L63Qj1rmfvfQ1I+/aMRz0ld
Xe94g57VkF4cX0hF3UqVn3vYPJBLIR+xTFuxcXcuLzhghnExWLpkSN2HURMovIItIUt/TVubA5gJ
QQ9kBHTyJz+hbpaRQgEy6ZzfrFECOV40IbjzcAeJNb1cFDvwNnuNdQsdkEN4cZPw3xAyvalunz7J
whQ/ydSReQnh1JZGrAfTdOIFNSN+Iz/HUEPLoRlYKIsplIJHG8fXb5k62saKfRS42C6Sd1tUpTeA
PiZ6UQB2m6YANzpXxERJERZvY6jm4MecIJfsHY4S6T/XI5sXC0T3kdp1d9jsgIfHhYdTuKCcRvJK
RnmKiIIn4Kr9WF1F0iQdzTTUmme8PAstZstA+hBy3kTW9uvj6M8k3pazm7e+2T/nF7G53WCsILFW
Gp95C4WjHeBHy7r8QcNA+Tmmn+UCWmSvMg435IQqEhAZSMojNQbZdi1RhRWCnJdTdai3WovMcDFm
dsCDHuNmWjq+48nWkoY7toIwq7iDl7+dWKmqkm4B31WmthaL9ebus/nmj6dvIma4aMXUeTOF/TyK
OXeOG4AEg8VlAD1JYfkgmm6dGwlxxqrhZtrxq0UmG4t425eBFOwQu1f4jY54cbpn6BE4rdeYHX+o
ftY6NMyGpzjMIsU6lbdg2bU6jvIfswq7fF4q+oGikm09fSu+U3qLeAY/oF5aLSQkrlUhUgp9zKHU
m0odVIYbu+cMt9mxO4W6KI4NVvnHfvkA0v1BLpVl7n/kyIYaewYTllt3gOEZBYdIhpOyamdwypQS
42E9+6vVzsZsbJo5x3o2hLkR6yQ4gTdBkdx0ZcTFd6Hx0X2zH+NQmHDptyGZYgSaxa6mVoMQLbmy
EW16pRQIQHtOSNSLOdNWXzU5f45n9M1mP38FjNObqqtcbjXWzheXyeOg7rbVvr6Ify03L96PYeTA
A/KcGWsTLqKC9TLiNIDnLfA455N7av17SK+N9tiXa8XbuDcqOJyz8c7ZFK4B83Z0gi0jvjC8Gzvl
qe4845ZdySQAgQLqhXIHItFg1djaNoXmjoojmVb2R2EINAzkL7pAZVx6bZIp9AWvcl7rk5YznxTb
FcsmeweMcUiuxCrLFacbcmPEyyw1r0nPCg+68RAMWS43VSlSf67FIXn01nbGNdkWobY2NfnzhDQV
/IBHA7ZTh8K4FNYxOm3yLpKVnkz7wEBKCtDAJP74oPkLUz7UbzGEvvvKUhmtLEjg60jO1CVbLOrl
wQ/BAg+IgglFCAwFrbP29h1pitgApqe9tI6uojbbwc8YLl+IyPdv/KRwWxcYSMgjd7cgtxosrW5z
rPOzVqV9Dv5J6hGiuhYM84gs+mbjo4+4zJnEj9FmUzTJZgHvEP/WlUqAGkStNeNV4oOvfUP7LrPv
2DmYM3hq/EPlgGxLuCj+JbatnOiefjCionr3oC6i/o+ydaXllsoz3GYlm9SXf7TP9SHNGQAgM21W
TEe53Z1kxrBnLETaKjESRpFcFclSlnchPsL5tnNDdhkPWyEZfkux/EoiKvyw1NRFwW37zGkSkLhi
RITp4O1siU6dak8z1x2vjNt8AhQFpigQKeg714weYKSCuSuXaOg+/cT2oeJxbpgIZzJvY+omjvXy
V3+dW0g5Jz/CgAZwnBOX/nYf6oH5SWXTsa3mTzyoyfLKXwzO7TphIvzW0wSz2BJ8Q2/jCGrnL5VH
elGqtnc8X9JALxk3QagT+myTDXDcGx9Kwn+an2GRLs73azV3WhlJultkd1J8e8M0Li5mZVX+Iwzw
2SUetGQtDg+uZJq0RWUBmrYeUzzfauwRiCOgyPaRH2TuqQI47Vo8WXLMavtF4P6aK4wf3jWcH1Tu
uWNeu0qzJ0i/dft2JFwQBPanPRVbAvFk/qspRZ3K9Djx84Rc6WMtiyi5oopV8SfCQWeXfo+muuM/
MJ4V+ukZoMLyhzuCvkwoje+dHtcyd0KULLE3+FGFRkwaoI9X+cZN7ob8RVNvcQrWeTO4yV4612bY
2dRMNPtbzpLSzbLqO2ZG8yiQbVT3Dx4Izz0puvUVGGCtVi9cX4HWyiQC6lUNE7j62mGnlpDzkFJO
qneBNKOmJaXVvKregFpK4w73QMvb8WnKnefD/YhonIQCVHKaFTlRuT0yUJnI1a3L1Jqee0E5Pikg
x0JG10T7Lvk5zGRnGIB0mJMH11IgEnphMFt+K4S9Gh/PmqXQPpbKX/JPgcw3GCTuZ6OhhgvcQmw+
eIDbg0zW0w5jw/X3EYuh4mpcHM0knGPMUV88wrZno2NCWi48dJAPZhJP8WHjXHlvoS8EOd8fhJWS
XLLpAPfK+aZRlMmISq8pauJG7sFgr+SsbsqPIS+AhALlUsNu2H4qEtKLPbKweYB7LY8c3flGpJoy
LzIv0a5mJ2/w3+DLSi24y0f+b0x3RHD4KpahnSTsnpCkkU+FUlJ5GJczVr1KnxUWg2VeL/Y/p0U6
jbwSI/ZV7wE3N6DbGr2Ljjtcd+8pyHH+N6CAjVidPDApdMYLmj+1pHVykLahmNmIyi0gn7NOoBeF
gOMQQJQ/KU0zF5eWLJMPqijDUKAYt8y6kzZcBGnjzuGW5jSZGQJ0/68NbMoxbMsHsfM2qghRMWMy
/juG9nPrqrhcMV/Ps9XFrJzuJuUW7lB2tVFFVUmoq8cqhtf5i8/wAHuraE5OyXE2IqdwkNozshYm
ygSAumYh+TUuaPg3EtQ6y/G0oLf6439o+/PuCvj073FRk1kklJiwjxqiXpLV1CUfLVDJUh7RPVq7
6I9EKms7F5zucx7p/aKRQKYcIDXBdAe3EADgr67n6fmthsTpRs2dai6kxXtXUcwWxUxp2657dGH4
A8hkHl5kJIaohM7cNczMSaNbtAwwD0HpRdfDL5xvBiI+7JMQySp6uQ8Fk1V6k4rOos6MLkkNAB0Y
j7fMXtpnkJmgLHNWT17+Z5L5C44hoW+TN7FVR2iAHKEDA91tW9CCZ6p8vYRLjVWoXzPgtDGPQPZJ
vummEX9xm5DZEp60v3kWwSoxfr6wCcyxRIgAeYJ09gF4V1g9B3TsGnqW4h7u8UVv08fZpZbqzyxZ
VieMnDil7Nt/yTf2D0l0igoyQpfG2+8NpXThQmbr5xGZVgtWSYVbEhYZK47SxprSvz86zIWmkY7h
OiSKunvCPMDBFv1ZDA7POG0qmf/0yqPp+CrpsFCHPKZH/aDc2PQ3WCO28K7TH8pym+AXR8DP60dE
tvdr6h4rAIk9K5OGZJomNs+NyhIJndHqfwyGu0SHu60jUNb65OgCdzsr7Lbej41YfYLg603r67Ck
MzIHMAv/W6Q5rTmW0bFqpgaXpxSf47fP5Rqmx4APr0c5YiBEBzgCYS0cRwODxre+/0EnmhpFwKA/
8CWg8bpyGsMc79eh6YEF8AnORV7fRIeL3RYYw5ZjACQo25fOXIsi4n2vGKjlt6H4uq2vM5Prcotj
5X7e5rA0rbi50HbxbVO+SE/KrwfPGVp1dy29m4yQdg1hqXNmHXzWqHvwz+elcXa/0j5xGk8GmUKa
6aTJIeV1lfDiy7oI+GCSXn/fol3PiVvH2VnSeJ7IlV7GCAF9qssWPSJ006DLgvYoFqUk98WpqETI
Fh8KPpcxCMjZEyPL5/hYc47X9Hw8uGCHssj2H5IzqaQoU2+n3I+8NE9fsgWvFx+ts0IPyHcVZStU
sy+yL/jKWMl93FTMh4hhqsJY/zCt9i47Pn3S0vAzD4fIJUpYoUudWKGExWne5R8nxnBbiiBICpIn
Yt4bqcS8uKzaxrvquWkCg7k9vOUEtiKN7JAncZ4o5IGyjYm+QQ4exHcXLoKgmasODPuCRQ1N4tDC
e8FujtzXa/mmbvcB1DUQRnFwYvaHMF6Qbn5yu9qa2wae+KqWE7RW6+vJn2SMvBWv8l7/yMpH52Gc
4fwrw/pjoNS2HUZr4GbOVCw44IkUvafO8zUUQpupDerSwD3+T3hgUfgYbUdzoyA1JgicJcPytzny
x84GdbORV4dOGKS5DXeQNw0MoM/DyWGvlklMACgV1yeF+3PnmQyrig1GlBLh5fBEwu3rouDRcSDx
BQnrU90MFuqIJBC95hxeXmuA2LRChrP3GZxoAx1s3Jen+OjNIR1B/uYGQ00ZUaoteVzlVxWIsQRK
bCOLDydmrJHBczZepQ6qv5fMUEDO7vHxcnwaqfRtgACHSmo4iUPKT+1ugUEKEiwqm3P3kNjZnqPl
5Ms5lvblKsm4rSzS5dGYzPoZKTX4SRhPILDDyVVfBEOLasjkA0G0yD4tkns/FuuH9MnmFcDQCgzq
EBSx7jkot4kpSyAquA+QZDa3aduzzc6o42TQmokxArS8IpJ8DxS6TmFwDmwInn/7Urz4iAEbN+Vy
zCOPfD3MVWSUhaT1xK+zi6ZMZWuKneSfQ5eqWHldCuJMtg8tWyqnGXlcxacQTDbbfJMGuZWuqMtK
KjK2yEL7oo3Vs3tvmrQxDYttlshjyo0KBlBdikJKky9ylpX0huUnMB9OtD40+88YzHzqWbjixw7A
4IF8FQlodERjVezVPsf0ovWmHJapGEiPHA9O9yc6YPwmBh1YRthtiH++94SZR8bxzfS3r9dhiZi4
mVH6UtnZ7CqRFnj87Zd3im4iXh7N1W5z/ljo9KTS0eviOdDtWk/1BTQLOvUQ/xUcwn8igDeOIh24
rPb69FfB+fTLt43K+RzPwzsveRi0lXtfeT68aqJB9K5oB+U1Bu3RCBeI2BrLYbNLh9X9Mq0fiYF/
TWzh0Is1te0apuI25WUh/Ntv9By/6Kgyeh/Sn0X/7ycuOO3GfjvmQ4iZN6IDbjbhQsqRmkh4Egd2
+BuHeJoJWSs2hJpqVjGJNM/VMs+uLQv7mdvJ0VTsj7NHbXRMo4EIPi62X+0bLga2ow2PM4A3LiYY
AwJT1HgvrZIaPyR6zfZ9+rQr3H7bGT5BjlGciY6ZUf/Q2Za7YU/mEKy2U4Z7RoNo82iSBwgxC12v
7Vi9ALTnxCuskR8NAzmug+7qUXn+9xFjLVtE/4ffIBZ33shZWYpP+LEj5VnHmNgA33w5pKePopx8
fvYiAe8VCE51K+wuj5Cc0gf6A7BMadzc9aWHy32xDA3ptfqmfSkaYxHWLBwn9n+5iejNX1BYFdkl
PnP0tpjWGwHOtl4RNWoxA0Wnl1PhY6PSpewn9f7dVavV6EgI3uOJpZakRuQkARyyYzp6DA3XtVjj
qOSonU4y93wdLP+q2w9AMElCT/sza1OIG0oiCqV8ZWQTT1fqCNG6ELr2UVAsZIMtCueEBOXgg1ey
jT9YMou6I5y/p0BGTcVmkRp13pltiFCXKPI6ZaO4YGj7KUJMggAhC4b4qWEQVQbBgPut7sfmHrAZ
9VbzO8wvOHdmNxGAhEs6cgSy2T5XtLha4/ZEUEKFGgRBkfbTCc/Pk1cgt3rdWXCC+dLsxXaRyGjz
7wIflfttOsAS8UKfWSwvash8whpcmPOkud6AtupFhIx8858uhNN5Ik76qx+ZkXrMLDvpQ4o5yclC
hha3kwx2uMz2kLYVDmFVDUwzcZVFoU5sHzYN8RVGvQNLuXT5zVi1ck4aYsC+WR8LljPhZ5ouiApC
1RRgjX2b0G3+yJLkbESBop6M+6I8uR/6WW0b4vWhkAy9b7d7a0YW9rXKs5ZOntK4X8Y+EcIvFlMD
u8G3hdUlYigBcLAeOjLCSm4gh1SZnUmCjxTNe1cqjphHQBr9E8hZIaW73mHkxYIU7beNmimJicHK
vTr+38LZoIb5jXPq3CkqCGcquIwupLQrR8NbuWfVrkrwQQrxPuEUe1k6SvIJKd7wZAmYXmvrW2vJ
R7QcC7/3cY0ufUyfKOcU/TIaL+IADvwdsDNbNt2gS1uHPYZ4rmAJeAKs7qYK+qJWlsit3wLsINlu
lo9zVVfJh8sJ+smYyU9vbx9v/ljq039nOohyIRFYRrOGsGuWgc1VNom62Q85XbayCflccIymDQyj
4MNljt+hPcxTW8/SgNdwIVCEgaB4dwLdu7tLTIrGfD5wsEINRigS3EcKOYcUuzAzZ6+vvxk69TvH
dJhsRARXsA0jWziI05PmsphtCnMoDXlbXG3OTMkrlgmyYSvxk35j09miqrD/nuY9BI9WgKGY/mIh
lR+YOA86BfyJXqIGFgi6bBCl6r082L/357MwBVHJS3OXkN2ZBn/ZzhKmB3IDoWJWm/u966Qu3j6x
45pGOJucL61dod84xY85rySZ4Fm2RivdGcN4e3+0aiiPrffLoBB93KYPYnu8VriStujgC+RJT1Y1
A6yqjYiILj9xJsi9xHt/NzoxB3D7K1eN/pzQsBKkVJM2D5XWmR2y9B75w+fQqgr1KX8RAgnFxPeL
Vl4fgLnLcWW6N+Q5rOCvMCikic0A3brefc7yd9ppH0V16Zl9RveoJ6jmZohwk4rM2gu9oD9Y2jcz
6NCTVua9wagccv7LZPCayWNZ+GvM3bwPny0rCghytLx7GoZUu7QFMRICNe8D7EKCKWjU6dbfd0sr
0i0UgT3RSJHrO7X4rPfydL26WLqZArM5xx4Vdo5LJfiJrx2wQX1KZzKwyDVE3a/GHAiqfDAcbb9D
XABUtLlF5cdL6o/NlFu03B0euH6fyw8SjX0qIopPHWzzySN3C0oulBvAVoqZoaYbsry302IqlhWC
Tm/O30exUQrgLOVlbsp9P6Xj/n6UiVhkttzMS7dLGaXDHLRDUzQasWhMFFh2PjdQajwf2YQRnfIa
RH9pNmMUq7nVf6TjvJzdPAzXUFs/SJ12P8stDtf+fxjw+a3FN11DDOwCfd0tIObwrZNRiDY909lf
4E5ybrDdFlxsdGfjRZozUzBJZEm9ski1M/9T1bqdB7xSh4bImn4mruGtpTCQVul1ELD7cN+VcCeV
46sxklTtPv9Sr6qXlaAhow5iT8yW4Lf9sdDM3Bf1J3KY6tF2AYRNDLvC+HTD2ad3EeFeMjg1EaM+
reqyJ7wqcojQJ6A+NWMaFRxyECPF/8CnhFe1rUoSxIXrWMX2qTTnUkjQyPVE+kTjdQFKsHcNH02U
oj4Lr/pXoEmLpKdU3Wnclu57EnYVNI0bLjtzRdCe+K5EM1FU7IRGrUNyWljvRvVQTAjpbdG3PeI5
i8y1WfzB+Na5QEx6NugTKolIvFB5V3+G8ADLjqcM8ErIegAdtPrWKphXwg3fW+wYYGUAVytX6x9Q
EWBfBFyoez98TfjZnAZ1dBG3ye/GvFCd30dY6TuWToIb918tizjBn/Zrq9jIy+VmzfMRFSzgrcLg
1PWxBOenleuLTiybilDV0WchCc5azZc22M0aTfFhZ86E+MZ6fZAHyxWRQ8B11oP5SR26qFX1Hbxk
Xi4YcTEOXg2kfoQxN8P2sN6SN/qzm9vvXWcUdCf4rieOhfb2XSZRTYZWcA9+raEIT92F46Oj/rNG
GwwFItKN2kcVa4zoUkoyxT2P96e01oUq5iYbFhGJXovFHKOpXpB/UjlEJUUj5AQ3e8PRiNXxzCyJ
p3csRHZgiT2BoaaqQEWEPq0Ys/OlIhI/8gf6XpHNvZsDE/ew+vH4YXTzz4t73dyrW2XJy7MkaS9G
PLS2AAw/IL5FhNVm3X0fNBatqMonhDCkM+kBeSCiH4JQqsXNGnMYQP3Ehd4hZ4fso+CuOLCoXaue
DIJpvxDn5NdrPlVvcZNqyJ9Nky6rRPtXcJEcmbmyxlhiY6hYgrH4P1vD7rtnyTOPbN2M+XTGFJ2O
RILrBWaArbHOLSEQ3XsmCC3aEMGqGLnU5t4iAJWLokVzfRYxGXGVksyaUSBaTuClG3+L+zZ62VA0
vMO3Z055B47k9AuI54KU6V9rgctTzv+t5HKQG0FF/cOKtAQIkq04VucN5ZYOubCbDsZ6R2kdISNZ
/jSNC3bt4kxMlsiwo8scyrBdqmaMWWGYNJIdvGYaZXDIDMkPuG5ZhEZnWV++9yUPLe8HTaBD+fkW
SZdtzOolej15OlrMF3fokaopAs52YsaUDdhngoK1qRop2Oo9T3m0tUOIh2VsYP95Lki/iA4IiJa9
RhQTtaUDJFDikRuSi8anD2jyCw2MNTVpv13dAVaZocQqkTNOYesjml98sN43B9TyJuk1Tm1x6w+F
6DHNEuJnQsEpZrjjWu94CCB00FDPG7ng1nDuZADSAYXxj/ECUmavLJrylCiuhAw8OyPtFQhen3Pc
pBnm8mFE5faCC9nnCOabTG7u/714n729Q1Rc724bhHNe15uRlaD4q5bxgtgXtTlnPFesGqOsA4BO
+FSiY8EsConQH3caZpqerrRLC4ovNImaTw/HL1pAAeUzf4GlK6rM4NQoSRcneENymfwDNsldun5X
WJP2sEizP7Z++W29GvpYeHpyGwYXuRqA9OYW9rtgN3CRr5ykYKzinETZFqhjsSg+MJF0EW4A407j
5QT1Hr8BwoQOKUVuPEI04WdSffeJOyGF4Fm+9MpDEiLro5cYiZwxna3PI9Wj6rxlJgQ9D9qGofdx
Ru1bGVabDkiS9Z4NrPXZj3Gr7grzeBDiVytYIUOdvWkJJlqoHeBlk2m2PaWVCQKv5257cTb3Mp1s
a+AVMRd1kqzLRAv6aIR6bJF6EPTvLV+THYQ/UZZsL6jDXPLTFoHUQ8MAPoojfsO0yTitvueCPBzR
Xo8ycR3uSQHJzb+nXQ/uqokUkwmv71f2uGlzeH33IcoRFhiwSyQbXJg36ygmqA1UALeFgODQAoAL
o8DhyVQi3tOTxSIWbqdtJrNreOhmBez0l0yJxjkK6hTiiLvWUZMRKgtxGpwvcyUYKXPrRvlqWINb
KHzC9ALCdp2QU71mTi/513yJaIdhGGrJCWPhQZ79ZxEgORWMotWrSvdr3vlUBkBob1T6lvcL+QTU
7W3/fUK1t/haPwr8z4hzlx4a8W+HSmZO5oLDpxvSOCsUHxx9FZOcyYt4VhQcurQ/c9hI3JFz6/oG
8me2yWvpYVx0IZJxN5Av5UVfWkaRiaICGmaksGXPn/eEQ9kUvJHJ1T91JslUtUyFFLTd2iu0p/zW
GrpjPm5gv6GKfdFB+UQMVL10eGhJcNE0umnuoG40fUN9o75hgvJmW5EB7jNoqIm33XP4e72e78yp
KJKg7XCceBEmEFO8IvOCLFNwbgbORtu2fRPB4TpKAJAaLqH9dLxMZV8wHXbTwN7I1WikdctyupUA
TRP6jRovdu+RbdIA1EuqBEgnc+vzsK45OTpd3Jm+hNHE75fMsPf8IMZTDzwE724LhgiLEba0P1h0
k+ptXxLoZJjimDWNL4WlhpDB86Ze2taTHwc/CHFk0bioiWXT5Tb/ssAlDAFVfhgSPyxh/TRyBfKG
2HmoB9vAx4s9uLASJNLq8auj0hormpY7+GGyYlBwmxDR4kOxvpgSmNTOshjTLbRKTREspJS8LqKH
kxYerN/3SVVBlXifmG4r5UVQL8YuV2tFHF6kQ4cYlMD76AIvKEJQoO19MIvHmqIT1t3SxYtcAhe6
4c6i0pVznM0ZMGLjFbunUwaoHKKPCM+UG10vMUtiRXXv/T+4bGqeRuzzYnCzVyLhVOBac53C8KsV
kT5zVagABpOSMyHdAglrx4ByGuoDD7nFmEjIPWlN1ZOrRoq779i/JNXFbZyV986Dz9neDwKM2ZMU
Unm+abkvKcOTG6+WziRcCLiqa7GdkQX13lmj6PAnR9KKF9bNytUtpQ5I1Eu1jifYtqmNcVyyphjf
x5geFbfK2fod/6+00m4fl//xulxGwe3NaSC0byNcSc6eTW+8MAUVDHwOC2sdIC/VXRXTTI+lH5xl
RVxugqoGYSJNfnoOaapaVLf+yUnrKfV+zNX4LcrRgP8pXIUqDwDRSWj+SxmGPQeA/7Mlh8KOQ8so
4Ir47VH77IwGaCQm/8VR0xk0+nFxGtNvDkHB6T+/Kh5q1rTGnCQLuxyZynC60onjujqo21LrcGhG
xiTkpG6pIQzap92ZpU1ercJgIO8JirN7an+Tv2ZzL/9+jXPDRjcl95ZGIREh+ngqWtQnol3O2Vyx
iHnRIWKTfmKKOhbrYrrfZt6f4FuYTc2xxPtV06iROh05i7/7gehLiX9Zk6SgzkaxaKQef1emLfOC
GQ4BcnGed4ry5r9+e12dduZzmT6INr1CYNb0gt7CkuvdLq9K9KHf1+1KLLRuH8W1QPbDimHQhItF
cFqEChKrJ6TcpPDLdDWWTVbwt46qF94GKxzGbUKkWHPEphHFSBhoLnKPmfbDuCQ4k3HSSSe8b6S1
K35gl7JsoqwyRaaR/pe7WFQeqKzZJ8UiJ8fK4TQP8A6bd5tZHbIkU4ja4G6GEy4gzVoeLcwiUfey
rzqIE0nl+jBIK2xKVjSA/PmTGVGRvybfCUYzuBSQc13WIR9F2T6rcqqJoHvvKARbs16EjchCejEo
WZsb3naEskJBaAF0CPI9TYHYguMSleZB33lrQ/s4DZSJPZJLc//+meeHaZQgLGpMIAYjgQXaBRAW
JEKBS0B0CK45ssG8ryqaSUjJF37SlBsArhQmkB9ZtAb82titOGRX1HkJEMj2RmvKLXX5+FBvpGgT
Ak44E+UX9b3AErpj59GEvqBuwzQk4E7zTy5i3wds5sSLGVMyfNx1v1CX++PekzUZfzgApnS1mJPA
tlJ0F3XqvgC0yWGU+S82Q0+xr6OE2kL7BUCLaX4aGiY+Vi65pIPvs+Tw4GPdQabuG3FKL+zXCVM1
Va2WBRoYvOETjlDsGGbyqAQjAHbh6VajBiKRnKe2MDIxrYGURMD1hPLfFUPd3CsA0ay6USGvaCPo
PzPWnhL3UxUnpBdW4Ym7hJlcacIGPI+Ru4uLa3BRWBhJE3v4r5o+UphiArBwKIClWBjmgsqFmHWV
7EBu/GbrIr0yUsFJ5tBmEgqC/0Hpvp2ff2hvcVEk9NWk1hT6d6VnxqBGabCF+rsR5mlYTKTdRa9e
lvZZfSYtqnFASk07573E612AbRc14sGIySYGf1gFkPP1lOh4WXe64vdlJ/u9HBRef5qa4caCciy/
GSjlolmGHeKyqs4niUIJMQw3iYtcMWZUdb2W5SdrT2wbiguPV7bWrXZ4A9a+7yEFFOGdTs+d3DJ5
zIHIRZeGItsW7so+F6MtS1c/Dw4bctl9WI2DKSHe3wy3bTkHRSRZHRBkr9crbpF8afq9psvqyoVf
xY+RDSxW1zoITVt0tzGsFpIufN+QoxdnCc+vOAIo76HzSz/T/a/N26+nkvHjMbfyqQcBzzpB1vBL
DfS80V9JIQa+Qka+HEo9yKDKk1+RwLPOvcBoQy99gms0/2J1l4jYxZf2Aj3E65GuwYbZ7JixISMW
FD64pWauruKArMAlg2V64CvAxeZlPjBTg3UvnNr1iJFVi5VIweWGEwQCE/Ix0o76wOIFr9Hq1W8o
UcM727bo/iaqPTD8urR3hLyb2jwEzJUJXKhfX9XcZlX09dVUqr2agpha6+h0lUREW6v1Wb/fDYHX
G3rY6NLG27Xn2MO9LXDErY3JUmSsD9c+FKoGzv4AMdsWib87JCSzl9Yc0aoFZNgG/e3+/mLQepls
JN8XCOMD6pCCVTbjaGBkIatB+eUBp1dD/oP6oco78PrWWOfuVGh6/fv80igzEXJEtuhgXnqubpPl
RM6uuBh4p+pdStDowmidz5ru6XnOBYx57Wpw90mYZkcvjbAYYyQtQqLEynE6j7HJzfdVorQ0WMtW
qmvDclnnKCfiAaJAcge6/bYo/IIunT9rby7k3vY5QkhG4PgEPRaAOe0l6pEts1sZ7CF8mfNcVUYf
+CVvWoyrdwmdd4nMlEfqMaZLaM33S6gcXVOcIa4i+L5CEHqK9BP5e8mkXASFzhYnnDzlnVO0X6p9
JgFx2cKatpJa3bRX8p3Az02emmGcp1eQuAP2h2CHDTM2kicrEiayl/9QnIQMnTwS0vAmleLf/Pck
FE76ByB51SzzxVVIPex2P6WiSxoBQq6YtzpVfA705mEYelapnxO3od1keDCt3hG1CxP2ShS1Fmpb
hGjsPeSEMHdCfNDACt3eh9tVbi+TVYpqUG8cRg/4tq5E2PlJ5S5cFAGwBcwbHb6pKKiVQW3BZTtE
BahswTcDB1pAYdaERNLDcQ85ebL6oPg2gx+d6XcEjdtFGCgfxIaiA9G8EVw/vlLo0qHm2ACBd9Kw
Vo10PjflUDr6PcKCpXApqgJMI2yrv/1q6ZfwlXEEBIK/W3AL/RpYwSDy2JcWUT94ep4bNIsv7331
VILYRLuecd6W0EObqT+sOsHHWzYTcTYyOl2kc5mVm9Gy/etAqAhgiuv3YCT+hNwzKVyv/4uit74V
YOG6/5g3LLAwyVtOZmlWtFN6SeVXpxaMqr1AMDrlvWOXHcyicCjLHum5ddEk6I9kLSQx8aFr4pGb
dWraYuC7qIQSmo9cxwsnzihI/0ekUJpstvdNwhvETGc7duiqQhRZowxEwgryERThMaQsdmUKh2Ee
jgxpMYAZbs2xv5eJJxjSrJ49klZFgKaU6fThRsk2a342evXsno56/soY+cl8Tbr8Pg8gg/bnplJO
Cr0gWUTX6Qxb75Fvta6ccI5lEGvh9DRHDlfa+Af+yCVD8jIR2Ung1YpAjrNec8AJ1JRiCCzxi4Sf
KNm0p/yI12illrhpzP5dacNbAKHfEip6wzl2JFfV8gvEAYc4cfs5t4Ff4wCRzQlUB6M1AnbiJc2h
IncANj/m6t3EkXgfgjPqnYuSRuWYgbWlW37ToFOVT41nu9Tvzcedf0txcJhOXylUKgEm0hSNBMkO
7L8VNHtQj0jrcl8YDZO4VkQC03/Jk6m3h5HcfEqaE/ieRIK2+4PYzP36NG8Ii6CHG7PmIH20Y4IA
sQ576tDrSz9GxvCU7IaVhDTD59KAsODbcjsCvSB3UGB7jKMUZryCTwMECXdrqcGaS9Q3xV/uJm1r
mTB9hTAST7wBgIys8onV+JsuYdypj33IDG1oUcPe+PrcqQI8c8nsFg524DaII6SKOk7/VpCcZ8+l
HH3b/SDGni0YlAh+DDMW4sJBKQO/boFUMVT7H8TRFRLCUA6XEFORbmSjmuT49sEP6gZTVsSFouYX
dSp7IZtFT38t87+WvsT0cUm3fRTQCucGhB7pjEiS4r1a9itBRxOQHXKGVz2PKKB6zz2R2JBN8Rf/
OLloztvzW1yx5gjlDnCAAyxvzopngccJ3I+RbVOmJ5NPDwaBWOdmh/nm8Z2MF0sjcyTLEWONyI9P
+qRrf0/xrbkYmF9SyAwZkw8zeTN0LVG64CFasbWrWI0P1uOlyjQ9fITX21hFzXDS+F5rKY0jEPsk
w37pbiW/QtBY78DjVzx6tJ/DAJZe6VY5cRZalJAXf3PkBSCVNsdNXrbmDTRgfEuj1KrfIgMJiUoX
a8UjZX8MzAY0nScLHc5YbOBAL4nzeLWKlDa33S7ybYHSuVJgQNVe2shmyOM+Ij6fmvv1xX0i41Pn
0Gy2wQHOha8nbN8+g2I8RL2aVbKyZzds8Qp2Y6aFn53x+Er/MOhkd8BfzNL6eK7zHKDHCEIZjmKZ
QYa7FAevvoNqaKORIZkRgSpLLfiC4WSQTSI0yFTyQokMIbFzLppVwMFNb65O7ddS9NPg9kggbphj
2kXINS3NeLON4Lbt9UpvLoHyfPUWjLK2hpx95GEQCjj13GRnfPVVTko6rt2q71Wf2Ea6gHpMzQKr
i7b+2s4o7tZ0x/vfaaq+VqpEKiOAGz+mdJQ8q+qHSSaYPwsT67rb1QD1PZOHy6psv5lH5z5mznlr
uGbzTxOKSNLAU8cTyfFvok5l+Hd8EyCkar8pVtDTy1YkUPikplSjig7wS6iGby3Dc1wecIipgqZq
hDXFrsaiJS8Pc+vVC9bOmP6y3trWdskl4gr7eHBmUdphEbBkX7ESIb/o530DEVoaADFSGoGSTMAp
vDDXFnPEymntS4XIL3XpdkPlUfHPDyvjcX1FZwth29B9V+N+qC+Ul8uHAsZT0KJA9GczdYp8t/Vs
qWxoI9CWVrVleg03PizwzQnloubom48V4hU/zCGnc7K5D7iUdnxyL7O7SqBw1GnVPXNwOkwxeugM
rh2xKKoet7QQcG+wk6DmEv6Qe1HTkHy3Lmb0ffaCqBOldtwZ6tmbWQQMdHosv4feG6KcrdewyDSp
+dHylQPwuy9m/zzLk+I+aTne+hQXQOlfsATg+JqzSAWfx4iUEb8lucfXweXBf/uGG9+yWZG+Yrze
6mkuWGMFR6Oj5RhTXVbuAKYE4PhJJEfSLCMH9oKB+76crAcnskJTmF0RVW+rm/IVP/kXkT5poHZJ
9kfhNE8JpX7NdYWUi9A1F09u864tS1wXH9bZv8lmx8DdfQ6mw7cKdJhavuWKdONo5MScV2HLKXAO
N/2nJ47IwRScUEaLNLFKb1zBXlY7PPtNa100vrtCs8mahwhCCaC1e57SjCNPHAZy7xv1xwsl6yWF
in5LRSF3oV7iuxZO1968zKoXH4UlcqwuF3hW3ZBseIhpl10WZI/0IHRcxBWuggki/dGc2J39EGOu
HJP81/MmsJITTIC13Ik2rr/rVW9F3wzdbj+ewR1HIwsZu/SuNUyM/0CjJR2V1nU5GEHMXOy5ZrV5
uLnvc96flIE6X5yYn9YPP8n/oJtfJ6RQmV8Kfh7M80QsDnbxQppxi4ovsxvZWrFrbAx4eRGzgkkE
wm+mDP/3kZ2d4Ruyz9mySBSYG3XC25Qph2IA5K4Um4Rys4WDULwzK8KMtjDvrLqrdonPBetQOvMj
+cGDcrtQl0ZbJlcDpMURHvVP1fJmvoVeCWbFoqTLHU0lGRKg3IayNPdezCZ32y0auuvtqN12Ll1M
RNyCd2Ny76fVaJqYgKKRJ6rcznsncq7TAShUbNPFqAUgUFJtitJvYwYiw+WNF51psepnM0Cg6YL3
ueGVTGtQ6byyIHKwSt602X/Y7SgCpVevPxXwf/CXSf5BM836H5lkx/Ho61uha9Voxt5wTuS8sxIL
OKyFHvf2iArzmeq85ghHLJjn3bwKyqWWbjj0pRxgLELB8Dad5AYHCZb9fnQ3PHPxc8gkEyseSTmB
h18FeBzKhP7tOQh31sZpKDPA7eHiguzbzKmK09CS+7IhpfXQvIB5JL5+LTM4yZXwXXCySReFkyUv
Ycew8W4Q7/w0I+BcKOWZ657N0Bt/0sJRAzx04V/rweY5DkrepbbhCEIcncociengn3sgtR8297p/
vrCeM9KOWRwzOCICzq70ftH2RBHkvLCsKPJ0DQ3/IV35yNBs6AbNPJK8zLAylzkbtlGXudfL2dgv
SMQx3g0/VPFo/4mcY4gP7ddD/L7eJ0az0VY9+ErBK3qY04YYJzmtEi7H1OUHL893MqEoe8HjD0IH
ss1VjMTBNS3MHSgonTlRRL65IyT9mpq6Vt8KqZHomHPGu7XAj3HnXr2YVPIhnyBUjubX7zJMqxMY
8yS9qA1gk43WLAG8ltVA0FR57Lm+//rU4wXLCgkr+3JxEPDjtEAhzxGMA30bY/DqNH6sDwHN9SLO
Yd82XU1wYr6keUH+7Pp9Hhn4lNjMICDr2LuJ+Tt/8noIFNtJ1TIR3XfCOKllqWI0SJTDNrqDxi6c
ESLywUV5pr4xqWuf3Iy3GXygpPT5YqybRcgmOqeV/4pRnMr/lTbO2UrFoO7s/0HMNsQNSyRwSGf9
EQiZ5Z9sP/ooHHzrbq+3XhuALG/3hBpDzGvLSg9omgzeTgS4AihRbpUmwjoPnDcvd/KN2+/s1kc3
VbZfB8R41mscaJ4QSW0jvgV/xN124ZbTi9eIlvMz/N/SuMTB6Aeq+T++V22SyLA9wTQj27ALEYcH
uPhNjLdVnEIK0mXf1BzFB+Ftxs5mk0mU4gbZoa33VX1btYbQ9jw+OWrO6w9BfRnPdwiN6xbbY3r8
iNawTwFBfhngrodQB9aqwEBnb4CehSZ6558gQk+4Dz3vTmCtmCUVQfl5R4CjzPC2ozpBXhPIvy9K
Gln4anuV9zQmYugfwQ7Lt24y4kogaoOZY/TCoW02I4izmOCTNelhyBpaPQhgLo0ZKuz8FrJv1Au7
iPYGl9DjFcUqSZozjXtpL9Gj0RtbJVMnqlxzi2kK1WEWOTpA2ilQJ7Ps1hGRvGtjYwIqg4JalDDQ
hh/CJCpTkMrUHxVvop0Re+xx56vvE8tRzSsH4heMOWRkE8RAKkkayv0MgGNzK4hAvDML2aLsrWQ8
1wJ5pO+hgaNSmXQQAJBn1Sn+Nt4OPmNoVysMTO3cnE2pLmqJ66vJBnPzXUwG+Bsh/iVfRoNpR+Bb
jnBz4McZjeAoG3abvsIBFc9NHVeMctnk6bBjYZWMKudfzFMPOPwCKkU1Ka3n84mGjlBb4AUllXof
xZNbshb20KaW9ncpK0me6zeGLjaJ34yQB+anQ2+qijP5Y8m+H8S3hffKvKQQWt1bk8w0/h/8Q8UO
rOC/UgfYng/1xozLxjU+sHMUes+DgCl7+C4GVKdB6pZinc46jyb3RFaBhjws8CsmtHlDZH9+a5/M
XQDwDmHhqMvzbgXwOdBRjhke+mK9NEA+uW7dWSz1ccq9dE6tBzsPK5fK8ZD3rHuBd9jB18UB7Mpx
Y/bYRnrT231MhlfvjqZrojaYV5L4jluwWIG9VHHFf0cLbqsNhBC8cFhLPTwP8R2YQiKDEIQerm5p
gn97GOQnYQs96rsS9aShvJAkfgMFrlfqSJps5m8nlfl8eBPGV16oaOi7xUBJbj9EuFFH63aH+JZ/
rgj97/LjbeWue5DuYmfWVPEyGScZTMpoPAeyJCYoYrPv2VpbWCDog00PHRKTYOo7t/08UvJYw7km
uwdHv2Im3amUZSWypNtx5q80qkfqjXg8087gaMX4juEBdf2B3rfEXZiyjT2swsuo/mbFdb0T3WDR
2cjOpi3LAh4WnQ60e8QxAMuHkE1JidefsgViOLdVGxpI3hgA2WqZnOaS8cge878DXs8o8OLvRMfT
BSWHkT6j5rLmNB/105bQqhn7TELj83J2y3aFZ5gSVSlbvoImGELh0K87OG7pOk12xcW49p07b1QE
UdI0QMLkzfjHS4PjaHlDz6PI8HOKIGcDjHFv2JdgutmINSTslec5b+9TZpdjlGHSQ1Vw7NIYatyM
WPPfaIQfesoYOyoic1qOnXrlGTWI2pMo3vt3tjGoXxza+hJc7IqKhRyyhimiUNMqbIRDt9bSEfeD
PxfW9JFKHgV9zDYGERfgVkxY/8gbpnbpS3twTmYvpdtwbMkMwM6R3BrdBp2++VGMh60RXTLxHxEl
LKWCi0Q9kOhQobTDC2qdP6FbHbWP80fIfMqzUgaw4+y9KTDTt91LAEeFaHwWBCircnf99EP+gJPR
QTEQbM61nE0nuFK1Xuyd2YxczSdyO+SlrudH+l1AYVJKt+dSRrcdnsTLan7/lzjxxXqK6iZUTFmV
6GekzzKpsHiZG/d3G+cRcodLjESCM94wigUvbcCEN9Roun1NOOrYp0SKHeSuMBsy0rzzdAGqJUy+
BnbbApFCDWHZTNhz+erl4XIK3EH+Pz9hKkYVj0D11VQp00cK05dkT5+jQLadSr+JhN5crfhi0RQT
KT6BuXYqIQqS8do829sOXVbPsHPzz7NZOFEscWP7QDJbokuqaTYb9m0I/jdxYomSWWDehkcACXXp
LZF6zCGVr00NewhMlQZdqk97vmUxwFBt+a1Mf2gC/PT/2JmgkGft3q3FKcZ7JbRcDy4K83RYYPoG
L1KAewqGzvTpc8kcfYjsJSreynQXfCW4Qh2ShEyqA8h+XsJ+Y18CgBxu+bTsGWKjjItNXxlDEOgy
NXYWBM8ulzYvQU1lCB3AbUdtfoNs7BwAUDgUVr/XsNBxEdZNaR8yZ8jb9/Ick1+QgMBLE9Z0SPJT
GqH54iUkffV5TM9m3vHrC57ZHCiOid2VBcmZhOadH1kdfvEjWYuy0JiP9ktRHoS1I9mPGJTjGdKm
6equ36sOxXtR/PfDuAPdZiiySv7Md2+5Tbflp87k+ULzuSJov+kueyEMybnfcC/dOyu5m/cB0wha
dp0Vp4XvUXGh1hkqO3ifYEO/w6IW+e8ljsXpp4e419eNIzwAF67sow35x+hk/WkbSIgCswb8abWj
Au1Z2F1lkTQG10yiP+T4XelWxPltmX1TWM13znlIn43HIk9DXKTG0jCHxRQ80JMd6LA3BR3ZZ/tc
UhXn0KyQkKIwI4QY4HR2HauJ5eb82MPnQ2up1LqzG7woolC2l5d0pwtYUaNs/pMWI7/S/y0LRmUM
BZHSXBRAyZZvp+ryE+70yvhn+MdYR1uv/PSOR9H6trwdlK/CJRdjkQHHdXpqSuVX9BJcDxaaLFop
Yt76ZzOmqK8DiJ7EVZ1VKzzDztGIqL2IDe+vPS0IgAEKROTn+RUAGAlh+qmlmQmRN06gYyS3vDHx
yjOZ8mQ2cabNIxfK1gDFCaWewcRmNnl7R2T1g9QCZTe5qFt8rZbWI+r5y13jeOrBgKHx+4dBwRZG
ZcpcI9+pJF8DSz7zqG9n5LedK7JY/IZyfzv2g0i2+9+EoGepmy322tZb8Qg1qHE198/CMl2/91ny
bXfRemrFSywdhaHWXv4T4c/LKOB3SrHnWXbUsv0gxBMX1Bizp0STOAzKH/InM+zS4UG9apmwud4c
axKiZPVfHWlb/XcmVJ3rtCq967louOi7f1N733JwKare4RahSOpPw7FVLdmqxxkPyrvPNbyjAgvz
JBXnDdLKZf9tBgn3sjYOQhue7LiSSqg5Li6tsPKPNGEdSynqiZND1qVXtlfbzxooM71ibZP/Oj5a
XyqGplSvfnhwm0tCs5iv7oqYfjVGn3DIRmqVeB538EHkjb09M76u9V2DdWqtdHZhSylf23Io8LND
CS58SR0zOco/IlFyBroqZYmThaUfHnIp4kPhrbZJnKrVVZ7ip5vMb9/UOEWHrrGw/64xpWSE2dr4
iiDxivpqVIxUiF+28BlG2xbfcAytABuls29tHF3eqKOcOpQSRMSIIY4A1loKmrUnXhUu9BkvzdfB
d9I5BUy2h1d2wFij/1caxbHgex8d03PfKVTCl0iEAovAAD0e90ZicvnDwP+6OA+/J4WMsVbZLpqb
GB/bTAlYK0bBvNti4kxVhXoNM0lqZ5Zi+26HwZ2nZdT+9Fph252M71yXr4iuyTsKNvHpKH/5d27w
c2wgvpOCydGQEtVogJd1oyGJys/NGer9BDCS1TqXjWUc2t+meo+NI93z5/mY93VySaj1IT6vnvwq
braOzQE8EgUKvVXyEOSE+kCDZXNC33CznkKmv6H2vh+HMfNkGsUVXxUFZSm3tspdQpa6kAW+qSxE
02lI9hx/2uU0WJ9s6OrXh67Ko1njOICXmi0mU7WFbHdwO+aUcgFAxVRFJnwwDTOS+KS88x8DTpog
kvJAfCqibdqMamjtdr8OLlCTSV0/yRSDH0fn0tZJyZ5FY0q0oi/X8vhal4SrtU6XGletft4OSoYV
wIeOBOoa6WJI1A+oeDvpdPE1FkPvOHetFrmvQqw9s74kxD5uOTz3og0te9QmLVuPhKp9rsdmWTic
LQrpSZlaDW38hrWHB+yyoA2jLSzWtzQL7PyQpguz+I0eJ67HDqANxLejRr47grHHX1haj1Kn9xhT
AIw91gaROsM4nitkReH4yj+2MX4zV2Puk8paVp9neA20totZRHamPBFMRNTo9h3d2t4wh8NsThR+
q7c4VUK+0ncuU6WHhn830XDkFg6iyMcNhzSAMz/2c/W2+cz/bJG8rpiJuQKCdcMSIM/I8gX2lgUI
szL0pWbvHiUlYzRFvr5F2PibrmT8kYYois+xVRFeWD43ULD/fihcTKG55MY9NtUTC9B2AO298j9N
jQZJY9fc2X7dMMzZqmyI02nZkMNsMTXGYr313scvktDy7UWvJdn+/ExAuAVgKS0h7sdY5cwJHjV9
JwvlNhdrREBtfxVYZ7hWKavdiLCdBPj9QGnp91z88Q/o/C+hYajA86MNu8hvhk7do9e1qaZ79Rw6
YB+iSEriGLVXyI4fknyyD3yNpMG8aMVws1tDeDi4HOHhUlGqMFjqh2+vXFOOkgFBBYxsbnRRitR7
PMT2BbxoboVQoQQnH4BSi45gK9+s0VYpZ094v7fyA4HnIOT0wpT/Ce3E17X9jTNbpnFgIp9wfCrJ
JscsA0UBnRQca5zkaOTNXiZbFOwusH5jpH/s2leI2/lpLH0mSu1vV8BLFFMKp1SS2Rm8rz7ZMccC
usDSG+6Yg/Q0S/E3j8wh8E1Z6P8wrwpbODna05Uwh7WMB5rhbUmKELLSdG7R2Hc+QUc5ow7HbwzA
Ay3TaftpfG8MEe/SUEHvGXWlaGj3GvdPfk6C2X/P0C6LRZtVniWFSqpMq/KafncGXcrUcgt93Qbj
vA9MyRyFJACItwfWlsF5Dk5XAZFnb2XZhMmrHCJdXlUV5UPT0si8hyr/h8a2dYEXoTg9vAI6eWMR
CsSjSwQI7S8QGzQ7you8QdHJfbnS7uGKxroYa7aHqU3rm+fdXc2WCVL5a/iSLlTWjr/JtCRPZGj0
FuSll7SmFnxagC1wQIQnuK4K1/1b3tWxLFGZJjtYUbssrzQoN/ds2kO4/Et+lffv7dp8VMVqF8j3
C0hroYt5Myz1D3+wAVSAowhAZ9004TtpDGJ/oy4gjPs6N/wfmoTunJqat8X7py631nj/ap6kr6Lt
UDKRu3FvErMDq0Kvedkb6807rshRuBG/tSXnZWa53NkJe0jCdeldH+13n7LncxYHhmQl1NGigEAG
6XANXlo9Sztw87bU2NGyvk6l1Kajrdbkb35+zsN667cRsPbuj1y4LVuOQf7fI77RZM4WHAHTvpoV
Y3z4oHJzsCXESuD6LAMxQVyFsOIfZK3oSO7vJ5wXihSJT21u0PnR8fM9HTSemVneBVJVF47AYJ7Y
3vNHThNwchKTxXH0e530dZ86oVlK4rs+EPTlLoYPdnVPUj1KY72lYFatjk8x2JdIF+Ze/f3ix0k7
bHaOcy+8N9ZBSIJy2B/HNmWN5Zgzd1RssVUVlSuqcIPy9dhxnp8gqgT1jkuNQmwt/BksEoy2WvqN
CCWxCdET6k3j7BSaF6dBVH0qHxHLj0FGXpCTq7TAhJ2faQe8wbXVs3M79o3p9u36caEukTqe1gP6
x4pCUlQ3M5NlgvYkJ2Bh51MPpk67z4We45MhJywYhjxAMYP1yegGCrvhRgzt8ZvvM8qkloYLLDyL
3ymuFpCdwhit2YnM+IpA/GjezNL/QrCWf14PMeQ8foqgAfRlFJkBd3/fF0ceUZ/5qVMioP9pF0dZ
mqXVCf0sa9fbOEuwIf/gU8Jk62ItyxQhUDqWyKg9R1uxXa5Rt/un9i6T+bQyg3Z5XaOELuOPGq/B
bJyMB47MkKkb6x8cPKVvw8+TSzKf8Ygg1z+yU9WUqsLMxeMeEybIVzObGrual0haqnypuTLOHB8+
Ukc977USgx1YSYhyLbtTDoRn9/KAnZuwCyLTu0RgYUDEJJJvkxUgM7H2aJTCEms8DDegGaZ2eJ9t
yoaNRozuFpbDpNNNMp8Tgq/NdGoApM7jV3/dsi2tOBLw00KFNdDuhQIStrjKv1uztpUso+/HSYaS
4F5J1m3Uc1Db8RZEtoGcp52PdD2e1Vpr6NGxPiVJk5AiG0qMjtfx+Bw9S5s2b/vd46RyoG6YqQrP
CMbgQ9MyJomRGU4CdHq+Pzo23rxbcTmU+ylMd7miCyI+Jrnr8j9Ut2Jc79/t7ILnenTFztitrIy4
3PUZ7hImLgJHk5qFuIT+ysPZpdS+78HtC3Y3aunrBIqFqJKtBXJ2v4S3o9DZcY933o47rnsfb+MC
zMKbZdDggcTkMomGVzj4WP8J9UkIiEevHknjo+NI9jBmbZ2tUwjQdo9B4Q7cq9Zyq/GBzWcqx90H
0rt4OdLRlVjq5D9B4c5zl4zxFebDNbnJuEj0E0FxLles2EnMPZaVS8In4eoc11k1P65V7Yi9ABn2
th0dleCOFgI7u+c2dJOTODhhZTB8tH+1IMoc5kyoLAUdN5msIqZnYpvEfb/EOnB4zE2ZEErTpsqA
9SWhYftQMMAal/TyJ4oGAdNuwGcHiSk56oDmaWSfd4x9Gj5LYwF90yRCg0zUpKcX9UqHFyctXfCi
EYRh9IeTKsjKXokYv9HrHunfTvsGZYjy6Gou3x9WwLt6O2Aw82ABpYYQPIg5aAnCMHQFRxVe7NjV
5b2Fiee9bXQEyvUlf6ZUPOHOIOw6ENMCuL6uWblcJ1dg2JpPo8UMTKkri5rHzfPQ8JOAzILQtgX7
1D9lKy2NvLrpbSGr3P4zLvcF9AvXDHUZsUWVwhFAPFS22c7rKeDw9zvx6TO8m3vx3Up7bVOwUMxV
5VNVIsgcZNS3nzLX3wh1X3tGbKfucHcTn3I1+OBbR1RJfZDyrtFrVo5MsRBRO3Ji5eIOclzEyWwg
MjSVdMC9ymJkX5mJTHrJ4KkVbGAc4M3aLI5/VgmFTUQ2IPOpdV7qH63Qs2sulakSJ3dXjsrBbbMk
sIpd1fLYiLtjPKnjSLpeazceMkS/2ULt2aGde2bXA9b7vUlaHWiWhVDc57E/PtM5mGlBC6WDH/D3
cvtTMf+pewrrx/+6uk+fryDaa1hdhLhGuR6OnFqA9N7fIw37pol9kZ2ty1Zu2uv9WlnNiUx3uxIM
HBJvhn/pppRUlETiP1P7bS9IBDHfDr2rM8JnZIsQl5hH19Ikn++ghnCS4V6iDJSNey1qotDtI9gJ
WHIryhvv5QJKR+TITRTUoKUPekvp4N3qzKMOtERi3YaUM9XiNNnYDl01gJ9MWPQoEBNEZofJ9z4z
T2GUoGJR25lHfztRzkUiB5iXgzC87sm9aqVMOGY9rAGhK1mP6H1SEZ9jzaMz4cKOUl5c9mP/PxTp
bUyWMfeX2ridgFOOIosg9vojDqOeP84Xd0VBFNiyIR4HijGJIaS7aiZwKoilUJ4QZ3zqHyjQnsOX
I14yRcv54Qi0tLheeG0U7VwPI/KsVmWwvLgMvj/LUT8hFwPoFYPHT7OaffXkfTf2MtxEeUWX9Q6B
6q5NG73PxmbwbdZbdwtAOxklGHzmo7C4+ypHe3le7iwGOEOitIjKk6+Ld25zQ6+V0qlVbSg02rjZ
L7dWHCsSUhcGJDJJc8l++Z8lH69/D5w7zdbx6a8FnN48xsOy0ekU6DGMZPMyfoxNEkm7JGozk77s
PzSciWw1sTZ4/BbW2fM9folRW6tvctieoqixGvc5tMfGQDBm7tccxwhpzazs//gVcFTy82SUXiPX
u9Z4p1vU9nsQ0s2qHSwX8XkHLsQep6y0fBcf3PB+POTQrVaLgzlAh/Lwg+CSzkkbQqsufTXKyGFc
fDvDDM7DF9Zrosl/Sc3V/GqgVW97md2H364NehBsl3UEoJ4gy57GdaRUppYrODBtLKiByDiEqZUd
Or8/qdPHRrcroXfp8lhFkUGGlOfP5Nd1Tb0jruWphqvpWqlSc8IlauaSWcQffxNKrqJI6oqizEdc
GcnuEy45qzUFJVsMoCnhL1jbCY27yJ6i1H52VXWHnWXHO9HeGJEl0VO7IE/zu7Qd5Q7TkPEVh9wK
xYR7ktB9C2jMZHGOAYPr8VycLEh7QzokbY5Q93/POUTsZqtbWDJec/bEyFKSOKh6tSBsPxl0sLnV
8ba9871UBtloTW1f56+bhrmjIebfGggRN9EAkqEUHFKELdaO5sIlXqlVnvUKX2jyMUyF4F/My+mh
k04cT5XVHJkHHlQehcyP8DJTCWG/a+UL9LvFKUpzn0H+Sc/ii5MQeQ8EaqNfj+o4Fkb+GenwyQra
qc82fhNYw0eI2JLhckSRUcARfgMVIH3+k6v2jABPU4/mOr64FbtO/au8Qni4fL7w/kFqWp86PAE0
pgYuGM13TzzMPPEEIbMPTU6yx6+Mj11SE6cjtfenuXyDT4GfCO2Ef/ZLenBD1cK5+C2s/+mklgym
jA1+oNHzXxrMgIE5Lvxmo5JSuQK26H9IuKKKuxEdjEo/zQW+srOiTC/v/vUoHRqNwsp/30MEhWuI
pomTDbcpyxUADwE8kv8oRnAacZ9s0/s3j8NaAQ6E9JhtdgSOUo/bwJzsG9yz/XFBvYc2MCDJyqfT
sUkh9HYL2lz/IIaue8Ilq5K2QxEVKpL0xM29lCjyRxfUGjn/wavQraY8M2yCCx/Px/17i1fWtTLg
CCpr3kCYdhq6RSY4vNNh0m+3jYJGFHAaaeGdrLHOskGQi6F8guYKSXu2EoK606JStWuAzwS0AnQG
lZAmbrWcPQpNd/joQCnw2chqjY8JkySkDPTyCiC0HoTDI9UoNfflFO0/w88pRX/yxGaUs4OFFfPK
4apStrNpFaQFBWhHd8VYmX3IBjUL0H4IATbjBqhREO+gvY87DB1NCMMe2kfqUl1d/Z665P148Wga
ssDVxWzrWt6l7vXUlUD/FrOuhk/L5PwTUeDudQSCiyKH+fmt2MVY/BS92malyv/j98vELnfTkj24
UdC+R0Dgd4NVN5hfBqwF9MCsNKD3uOtvIKucvuF4E5H/eYgG/KybShN3nSyTEwyVcHup+Yw3+Qw+
UZyCgsXc+DN9DqEKTIrGChmtK75bGLnHqrIArPI8tnQPSI97fHr5bCQit9rwgNP5aQugfr866qxO
ZE0AMZPJIdjwsxSR8Sf0/oZt60AIHXa8BIBn510yt/hR5vKly7bAjrPa7sp4+B0IDEqBRrhokzjB
nhiRmoT9UKJCc4hWX4qopUdoWx/MQF8nvQbjfKE6xJrS77fbQTZp9R4o1l/ZIJ1QctwkSC2yF/ui
4WsVY1aQAg98SnwTTiWPGJixJ1dEN7H7PLrnXDq+J1UelDFQciSZ/Tl2mTG45LDAdQ0Q7mQTEZ4R
BlBz3g7jNreiRiv9cOZUHLdLYiW34tcHm6GbxJFQfBfp/sHm3bJcBHxsFvBhqNfnt2gyNZocgATZ
o357qHDs1olu8I8cznMwZuU8iHezjkZDjwTDivZvFkwh3aphWa7KYqlSpO97o8w+Z9Wrt55ZMknN
JOMz3L/kb19Gy920xrd7Rz+dY7TJJrBJ67L/sCCcs+xIaBS5Agiptndu1nZDNT39FNcTH4pBCvSe
ualXwRJMrD9lkqBXD40cjyw+V3TyvExqt3mhmhiH9h4K1ZDQfmMtdIbfQN1vZA6kvx7IRnBevuWy
8FWc83cGQ0dHpOi9mQu18CTSguC6RrfdDYorTaqwnTWzIaP2qcONaNYI+EzFz1p9eSLcUKdbar0M
EUAHe10je89YnIb0gKJfQmE+QlhF2I1DKNsFsLX5ZFWlqnvv1/QNU9aNvuCY66VhcJB04mLHxBsf
6Io0U5NB2LTXW8EOtGnPu/hPTqwTEg76Eev8P+iHgb27Kf5nHDxSj86LORE4prKRLbiGbXLY0jqt
AVi3uCnJWYie6/wuftwKMXENB3hPv0TAn8keoyEka4zsSXJ9MznXdI/4YQbps1rkzUQiXivSaldN
ECzUiaNucst3oUZOYEbf1hQ01DUdNufO35wg/rvE8nnoN0o2PNJ29HnjXj4VoyQb3bpQiVT75+1T
lPZIqO3mFowu0A3fh4GjJse69wWBasWsVlCiSvYshRRv99UGiAI/YHwFb0TNxH1msF/Q1FG+wkbL
/DbhRwoW736tgexVJwEuuF3WJtgRlt7zrX7ud5qoUT7n5zHZ8pG9N/l9dXQ7OPXAqiYxMgMIcDx8
Mn16+KT2d2fZBZ/wmsc+TyWeKHy2K8Rz27VuvGQGnCqVSDFtwXuSHQ0CwFzHK7WIzoMEJocXjj02
lr08gIEAbw/4HWpZGl1CTYjPvTzzYCUmx79lVQK0NMwS+rFEcptOdjDrYpxxb3gJRIX0uo6bT8c2
/ozGenhCo3Fxt4b69XqAZQ6dcCCsviyyyeYmTEfEbRp9P2Voae3w5ph9anxnJhfJtrE7XsBOHlRv
373upo4k3QZehENlQwXrlx+82PDbjiFPDJqlg3vj34JuAjQcPAdXMgcGMZQjLKsG9zlfhnx7eThI
RZHUibce/T7+X7h4PZU9gFQ5kEZa1eljJXboDe3Y2mYQn1HYWmPuqr8AnfGPdY+N4HvirEIUqaym
u9MMY2GW8Jk56fVppO0GYOZi4cP6Ss7vjkEhnGRm+DhZFYxLxDARvcma0b01omsq5BSS5r7oFe7g
qZidpWdqlbv/jRQcq1M1gAB+3ZRTt1rgdTros8TvUhFth58NuDgh86kBsYNRfktR3pg/iMRtCS1G
5NdBGXfyg+g+LfGOJezXtcMGksmRhLF56YK+vfoGfWEzGFq+loryBb3R3cf+AHHq852w2DdVzDZA
NORgPErq8BKtifit9T1Q/aii9W9VUyt0YcSFWl8oT/HmVOpL9DENK1KyyvbsUAruurzFfYVGIQBa
tbdOeH/0Py0R892fVXEei+i5KWIR3It4gercDfL/FVR5GtJj371T58kYGkZYaeS2llu65ZU2g15y
sdYOF56V/ob9UgfAxz480af7bmtA7VGLxenPeUDCEQn5djYADr3d/DPmhgiWItKKqcJzLgAj+Ly0
p1KOKpSm6UB06JSo9CnabUUJdahXGu+yecMzt3ai7LPak7tLG9Wo/3zqbZ1P7HmQ/1rNW8hZd0hJ
tf1HylHLNUAJJSyzW6+xN4+gCQ8r2TI9Q4O0+CszJQEhRzmSgBTQJsY6WmcC9Hv2plErEXnX/zcT
AUTyP0Do/bORLReigBKfwvch3yqmq7GTVhFUQUd8DNJi8gmPEdl3/LOwul0PLEW8bw5RWHSU5hZc
0yCK9nck4NZxcunrpg53Y23fNcz+3U2PWkgWZZiC1D6vTV/YDdVx/lwv/dz6yjizs/yMb6axxyjP
GreCNGfXVhRYGZ2Bv5Yhz7fIZW0QgiMAbwGa9VsW1ho3zSdaai8VrZRUhSWrCKFxLUXuyqIq3oJT
vDk+CbmAE6S5IPzu+JfspdX4wuUiKA2/12no0sjCzn1jQtO7F1Z46IVgS4QEtlwtL/SUVUaCusPd
F3xoyWr4SDUew3S/lq7p1/pBMkTX2qnvKMRkG/X9vPyS28kqNQo5r4NE4DCAPhnhZA+NyIJLmXTg
rB6fyxbSlgzHmDxBqkd3ay7Dsv0uuw+0+eIv14qnQefxzybNNQ7YPEhP0dIxlYt0Gt8GsOGArZBm
70h0AhaIg6Idd/BCnUeKrCADYVsT1WoxJAYDv3mVeosl5n2u9+0ebC/Q3KDEam5uBC3++MhmaLFc
zUKKdjUS5DOxOg6IQEB9umTeSX4fvjqbrkzk0inJ2AQD31qoLOz/K2PGQSUnUpdDgX7Ibjzi0QDq
wzL/aafPtRGiS91vBLv263VRFrAPu8TzrWAQ4EFizSN4gm106g0cxZFhI3uDvgA9X07W2SXeULgj
JGxB+90ZJVU3g+UQP5apVNdpv8wkndbEEuU4Sgy+prB009G6GFODeSZimrBg51QIOsL/tK1pqaa4
G0Hg3tj/8NKtpMFQhynAys5x/pe87wzUyvz2PWm1SjJdhbCOx0HSEflxnzdfOTE4cK1HmrG4FA/U
wCcOjYwVbiwX6pCrn2Bizci5C68YbEXBtgZBCt0wjX+r2s3V/W7BWNwsYJRPbKD8EQeqvCurCJgT
so3P1nFiNFQ0Ud86KLmfRZzPGrzBB1kDAEOjtfl10yoh1DtfDxWQ7RTHP56+fRYbd0hTfG00h2ov
Q//KJTFhXWvH+q5L2iGxHRVlg5S9mNxF2+F5oVOWgnK+csMejudptXzK8uiRaUHceG9rIFwGnnP2
QzEk1o5+Vvn0oXI47d+64GUWdVVyFdRfNJxEzf2+u/Y3pLN4aoJR1GRjule1zk7mjTXBilEHOwlM
gz8MwvoXnXX8gg+YKFUDGeHn2SuNQlGk0hTkjZ6i15M0+sbhToW+CRYmwdf5YPEHMqewgeIxeTcH
CWGWIq0lwOkgTAryn3VDTrrMrjOGXC7vXVa4LqNqdyeooystmg1x7fWjE3z8BOsfKxeJusVDh94e
6ZqAdwVCo7aL7YLsuCwmjWN/c5OD0Oohk1ry8FKuZ9LhimkF0OAIl+oSLMNB4CYshwaXrRSczcPO
oG3XUCwvTdytvTkHrDgWUBf+bjBc03ezDiGtmbZkiTNetZosoL3/GIOPnaUddA6FhROq7mO+tIC7
cGVzcdV5D7nTlqu2d0lSmEDv18kQMQ5VxfvRT0p4tX5gfGhG4oWvX88U9rEEeGlfNzzx4zE/3wJZ
QwmiCjUM0ijoOG278eFTxw314Ms4PGqd82oRpqDYcogcvUfH/TC1AQOti0vrC4IvNYn+M7etA0Zm
GjsE4T0q+4vIg2WN6dmhGZ0TD+QVFHld4g+hjeMq3lvfpD8Pl7dhCIdR6uJN5v1tYH2DTHkbdix6
fA+4xMd271Xi84hwPCm9qiTn/trRLfNcKprf9vmA4LOvthVzLOhUegtgcFkwEJHhVgILhhcLKNGU
EshBMZQ6rIbjifEsbZVyyjh4oUh1nXCpqLIbETN3ilAKO41JN2LbNM0paD2JI765RfzO816NHSFr
FjbsrG6xHpnEHemzWOdpwd9cmcAzdSkA8MDR+xWwzG7QGC1gKVO9b20wFVYCn6CbJ+P7hSWU9Yc7
INsnFgP0OD/kkeY6U+9fDwEOCffJ+Caw91xVfG5QjZcH4YB4/NXMcgaogIjZmp01Y4PxT35ioTkj
GaginOZc+/ubwqCY5NYG295CDaPxKqS+/sZg8nEkatBv3L2tciYl0i8XSUQ7gwHk23SSvo9n63yh
4SWqJM8SXJTJAgMdnt/v7lJ8sNaxL5ZHXwrW1g7eld3Ti+BShZ0D5f5BkUOmRylS9UMDMOByLnkR
VSTgk3RS1g/XlsD24P9n0NrufPw+rTev7mbuYo69kLCNNwoJo4xURQt7tzmjW+dqmXfx6ulDQ/NL
RiFpOJmZqaXhkkcj7zkIEXYQ8jqaRMUwxZ8E9AKrjf15/NFCoCohmWehkHLXFGPlvH15NvVCeIIO
MU0N0jF2CXXc7IOM3n+A7bdGD/FBFaGJeeuQ5EbeWyCFXCdVD5aHSu6nqGDpLovDFq3rtqBYYHQJ
v08ULp6eJmLUf6Bj5qdhSYvUBQHKcW9PfkAr0gdFNZzdAoB8GZFcUzmOciBp8Q0CSE3RM0CbPkVV
6a5p/Q/HpX2VxFtHS4lL/EIymAXjDyBnFQw07r3+O6YW406gQi0LpxgthoRWnYD1VAFS7eEGj/K7
niMYNPwXk9nsJSJH+CNakrcYrUbMoW4pOom+j6FhWiw+wGQPOK0XMscpXfMhfSDXYwu9Z0ktNxXP
ULYpb+EqeAE285exxZfdZPmso/2m4tR5NAVmCYIOvHrMVh4NJqs36+LuxoiI5fQBX4qRC9dJjr8j
ZTJw8oRfqE+sE8/0FbZGmtURT74EKbBRlfcUci4wpFLe8FDk8XXLm2lfF0vtLaU/aOlsltk49BjS
sImTnCQF279CLpfehM8Beb47jS8vGysfdtTri7Z4voAYliwEQ4WNm1C8Gd7mxRCOaRTbOWMaE79z
onZEUkCIbZ9w2m84EIF3vxGXberZBftd0RUpCRErlHTh0O82Uyv44sucmIa+vNqfuV6QtnLBEuRT
3RQEwr4GYg6ecxMcv7i5BD6anyEmfNc7Kv92B46o4+rxZeLlyVg4rbc8Dtgen1DDGNaV1/EoJ0ah
Z/SF7dA05jeseU0htpqDDixiGBkbYH7INAIGpfauweP0CMOcbvNYBczZ+3tdh8VG8K7JQurwzkg4
7yUB7rA0Vwdcyyy2JclEm1kvieqyl7n/Q0XuOL/0FRpkBxxoP7BaqxmSF22K92OAg/XfsIBztIoM
JiqNY2e2v3QXXM062jWUmlyS4o3jc9NZvCsFfARoIrBwG2urkCI9LDn8snKpspl7zxFCR4fUCSQ7
C4lBGSV94P39CS5RSLXGJI9NVdhfRR9exkFe6LFClOpF2fwgFDS9Ds1WfMs1DZo2EfixXaUklz0z
CdlOe+v1Z7YnUMdvAsUYAM6x1SRbQwf9e3QLsY4QeUkepegHVn4FVQDgsIDwvYM71fSFuTFht/nj
sAtdGlIWJQWx6kLhXBW06+wea0VxfEDxsgvEJJDJlxi1oXMSR0cpKvlLL+tI+LlwAUwM3ZY6RmrR
htKY0Dl+kjv9cK8GxwkIaD0ukqR3lYaB0GZhbONZiaG5bIxHqizlVKB5e1tDooOFCPYtwmXkB0hm
HSavnjjFUJj0ImIJjNnj270510eCBr53wAQOFQRwrcrbZ/qDMyPvsbnSjpd0dAeSDV/ljOd8fmrq
kSufFxpagvS3p9X+XPeFoFqeSrzbZo0v3jzvr/iIRgsV7TxNSTAp+44a5MjLM4Gq6ZubbxJHopux
BNI9TcDzsyuwxm+lMHjXwkIYTjgaCVcjwPKaJ1CEfnrPbz5g5GVBAuCFddjRPcCeIwkdsCxoMqcu
fIm3ry4kfz1k+0KZuhVYHgsfbUDT1r6yGzbxF4MsaV6lX+SkBZPCASwpPv+UnJYml8uRsrGcTvzI
zfWWn5VTEDDzHdOMXXtfoTs0qt4V71m9md8bjZSmOPaDFFZD4sQJGoDi7N338CAcs2/us6jAGuOe
N6mywaeLQtaZVBIF8yHHTWd//5ycXpbd77b2/4rl1rUGQn13YXon8Eof3pKO8BWYKPcmf6Eq2yW6
+Dy/DJA5J3Kb1UzaI5qwRJCVJnEOy4Awh7aJTFHo4VHez24SnCU+w/R8+o5L1hkLs2nNP/XQhbc3
mHGv9mmc041VYiPx/qF4rdN5A9YekEI+al+xhVIEhks5zh6fio1E4x23ksMO6c+olXE3GnRFIJjb
snyIhhKu3y9bH+uKenwiGMut7Gn87vwKAwjHRMyvbobkCOLRXbHKCivRZQ/W6RoD9d8tsCFXGsrp
EM1UPG1zeIU4UkTUjmcFe6ZixRxDhcSHa38mxEKNB2x8cz158s+HaroZ0N81NxurVHRvsGZUKGQZ
r9k0wfDFR9Aysv+IVIFqyyK6F9Z8FA3cglak+yM4HASJKZHFID+3mL/fFfwm7xfgG/TqXHABeDRT
+breD0rQgg41t+Fdpkyonp727odMWa5ntesGYfBLACVFbJAmUgNC1MdyBpt1B5GxhL9Qf+U4AHt3
68orkaF8Lhdv7deZzAVnzygiXxinYOWdosLwamSRBzoF4/GgB5DJ6vjYbsAmKd8fgiTiHX+FV2pA
g+5yRKCyj9gW2/qL9hDs9pt0Le3x70fo9r6guO8BJi4qzDwqM5EWzIIo0oM5v7kIz5uaLFCV8XPg
xAlIHDXWb5oorBDcpY+d2yRlWiHP09JVT0kAjEZna2Awphnl4HTJu7LQVVNokE5taWcfW2fF8X5C
23tuMYVdmDLJMHo1cCCKtT9jEvZWg4OBNFb3V426j7zZp0x3LsBxR/3CnCLp0IVbi1zQ28SD2VwS
8cMCc+XTSYLZ6PQDwzu1BOLVG9b015l6HRVYW3mYYpMc5SZA6KwrBh5r1C54RiBINVlKsTD0tsia
wH6ylKuIqY4Q+dl5z868MdSOvDHJpOTeUqXXp4Yvc3R4PDCax4jFcFPSsBjRMNtz8zqLaPl9WHh4
xJ4j+Hjgvy33kyhIWg3btq2WYKIOdKLyBSq6Bqjh1dKA1KD/rQZO5qwcFBNOHrvLXAcl+w6J0i4b
63SgvVM/rxg6y0gV+cnFYND8yE7NMYZkWao9CVFlGUlDUVK8F2ZCQ4UfmRAwsuevLqlX5ULvU12g
beOSY1WT3XYYNo4Zl0Zrs2slams6B4VjrdzWNKByv3zB29sDUiuI0FQTrznJ5LNhf14O2kVJAeKi
TRdVl0AmfVNuv/7li93xaQnQV21GeNr8KCl77DaaUYt4pfSviSKjF4NjmoKJhOOF/bqu2sn0H++m
gMvD1mNsiJLXBaVJN/j4TLsnnCC+8N1w68nODKdGgFJt3cPwBYOm9DyVd1yfaRoFdPDaFLgBSaZB
m36KecJN5QzXI+ZLTlZHbu8Nwleep6GtIFwcvXXAlNMvpoCAwlwm81zBgs+MiL9CQN7yglikjCtd
nva3xd231kkYHbVbML4jR6fzM52li3MH6DCsBovyxdV4QoPEC1Si7SLD0DjkiwUw4ioTujbhQ3v4
NGtLcQdEKmxt37p34ZzT8B1ByWQVDA14dyFdQ2r/if+SSwfLbrxtIcTC8KFr5XG6Wo/Zw3bWM5MQ
74AV6XFFSFP90/86BgIoKDa0lHoHGgJE4qNkB1uOQEnHFoc+e7M3IwRbtB7z/v4nvuq5xtZWQ7og
65JsHJmRQrPKgQYyb+pnILIQBaVfGn4wJoNxr2iggkH8uxxt8B9uG8DG+vhpzV8GWiyHwoIfOLR+
C83iai2YUHxB+VUbnrxGTf1f28AuP3PCygOHemIRvbhnGyFXyTgdtoRp1DtvqYhgPQNNR/KYAFjn
zX/UYe6ST6ZSl9TeWkduHlmpLCM+zoKsH7Dl1kHxPLRh+dUsnu/am9vNkIPaZ4BVpSYYAi+tJnf9
roxgHFeNSQWzrln/1YevOBJ60frEANx8gOLZai7kh85dMPvLXUJL6mLpt4aFXquylHxUcU85fGRq
DKbQOYtxyEt0ZZr/AJcRHacyAwISOoCn6avlqEUmY0gH1IqO5LZFOzYYvCpZm7DDM9fHqVReOmwr
FrCXU/a4n17aWQtVw+vYzDL0MH21eKxb+HefZ1j3AfP/DhIzhB0Iih8w1Mzdbq5AYadg3nICAEUb
pgGBDiU9u0O38DCCV54gCo9zAURtz9xoZmzIzmB8+CvsFcq3IQLsg2Nh+qLCXxjwN9D5rBhpjIW3
vd/onKT5RSfaO7BDsA9g0sVjfUpM+YdgVlKaBUIekEiZEIKtVgrz70UpISCUD9iA0gp/3YeFnv3W
bxz3C7+ZTDv+wuI+X7nQCSsib1hbEMYZ97qe7cJ5wic6gtEjq04S5fuzUsYZBFPcdI31rIERwO0B
giT7oADrqWHJEcOk0Ug0Cz5gC3Dz+yUFyLavljJZzItFfjsRJB6ymphZLxNbZwa5qpmH0TfWxN23
mDPvOkDJV/KIors+fQ/6jW+MBULlIz6ueu2xHAFbS8Kd/cWbmtZpIxTFqbp9zdQNU78J2ppBCzyk
SmlfR1SIR2KgsioA2MaeYxlf0cZUfadtB9fauGukRfnpuy4GdI75q8T9jw7lgXELgRP/Wmg5kOCS
YYQpOOS3xTbDPzw6fMVhHM6S8S2fqCmlclTkd233z+IQjRJqQZO129iyEValChpLDh0zHpKqq2EL
fbB7Zno5ojoSFpODtzy75ZIPudktzCTZz0S2G3Frx+dIRK3rqa1OA0dZLqQCdz6WIEHrT76DFWIW
muUR1WzfYbYnil+3NSaBzWXSPWWaUJFIaY3KB7AVrv24HRNMnF7hw+kBiqRiJYwzCL5Gn1xqZApy
jgkLviuigoNeWVKd9BxNh3LzW8reQdMiu8lKTXuC7eLEqL6JZUuuc1WbvxurCdRb1pDFe7ugOguU
NjJFKvQ7gGpqW4S0ajqIntplqR4kvHXMPCu2sDUc1D4E2lOPXO+NkbQDGPH25EOHVOtf9VBVQNSs
OybxqquzBSoZeFMuUf68z8iHh/N27CvInqPxpVS1mOyKPDnGzdF/pIuHpVS8GQl3/zkkzdrxd1G5
Ykx706z96fkjrogH6O75ChZ22LsFc/qu0Q7nZhP90DM4Q46GxQXtYfF58kGKnx82vGUPCNtC8PhS
o1iBFZFF0oiHWiPXfsH6JJLFc5xkg5zYT7HA7J+nmcH1JFhbqloAayKZQMK5zqenBgRquf1k78xK
Bd5RWb38kr3IPih/rS5RYIqfHPvBDYqCQn+nksEmR+eeDT7R9W6Ip8nSb9kpRhxKxc1o5wtD7nIO
9UAc5wQYj7R2tNKi5vTcfCRvFFbH/BU+wBD2wzwGfTp3uMw21ePcymtpEZWOkctaUbXLIvkxhE+L
0XiFmowcllQLlqQzKKZtdL9QbUGJZRWwt5OFupiL4sECHKBgaxn4V5K2SB3+QsUFEqYMHBvlbHbz
4AhJrBYTwzIFYNWxeFrs5UqfR9p6r6l+WyDDJh6/6b2PBPxyBkK5adWJEARn7Kf+ZIfPJdszQcma
n7jvlpecYQVkzNqZO1fR75msK3pysxmn40A9KVXWhDO5buTKk+I21jWz79I4Vmxllv9OJElU9F8T
1P/DNdme8XEhryL4YbuDjUyrcCav0r3TKfPegGly9edJ6K/7vpnN+vcvKKJMKbBm+h8CiphniZsv
cv4OlvOeKNrvwWIohVMzSzte7/T9NZBENocSe7TSfgz+OTiWDNG5tWt7AY7lnoq3QTWZMHuWemRj
ocCIhtDogkDCUlCR465CtwYsa0eB3rVnq7uJUZNRIjm7e5Qx15ZVYtv4Y55KONO4KYTJMMnMToyD
Z05Fi8KbMRO1Q3DRjgR4w4nWQvjukbH1OdiZfx2VRR14ZoQzS6jmQFWEfvf1XCiWKqXu+Oy74U37
zHQgSEqSzNk5qN7fLkGpZhy/r0z0dRYvKzwcwJPSBA9GwXPXeEKnMd4EAF6VyaDwAoJodmsSXbI7
+K/zQ6/oyb56v19SONpYIKbeMZ1HcO7W4uqUO9Qt6gVokH7Ubwh42gMsjM+ZYQL85Y8SA+yelYx6
rXpM5PFJFw7rAAe7ObZZ88MM1CIWTsPyUWjT094GNwxf8iuIZf7ugTe296QHII6YrQ4C9hYCDp6Q
F4sQNfdCBjP5/YE66EVRA+3xYWTcFJrB68evWz1xX6uwMu3K1wkhVI7GVvtLQ4GHQN7v2cOQ0ylH
qZkr6jHLMdphDZY7nraXD9nKDy1K+HKl8Fyi20Wr4Q8UMJ8bAU93oBPl/vNgFooBEAeBuFtga4sY
YWLIP3wZnWwDdc6QHfAfV+xdiklWJPa4ZdHslP9PAKbFGydPecwhyDtaEuZ7AGOhc4b3bLtznLVu
B9pafUiQN/AS6PFi9uoC6wvPJoW4F4VhU53Trag/gqHaeVCPny6V1rBzA0hYk4Z7HRp+XdlQm9Kh
ux08vDPrfeFy8ZYfyMXslw0rybm3ihyezDi96fxNS5Dgon6KVl2t13OKVISqYakUlez6b1t+NQk/
W8eqpxcfbhfC/1OT9jBFMYrc/H3sxFfJuXs7YOvwPLHXBSdQAr9Sg8JoC1NdmzFdMFvUGe5EaBIh
ojliiS/ROBaXJTvngIlTApNRXmQj7e9403PJMdejfjJDDiT6QF+rFawdNZK/4B2D608xO62MCXsv
88z0HCvjzWaqKPaM6BXwypYG+G9wQUyYdhioDfI6kTjGfInBaQ+gyWAvdRC/uaJBtnNMbhIUp+R1
6Zs7d1gZWikSeiG5v7ce2U5hPnn7bb/A0ABQ8OTsGp421lFmVI679wgG+lBg/SNlYXrZs/WF5UK+
1pIobQgxzphKf3CW6Axbcvq/izaPxFKK39KwRVQ1KAeqpXjUD8xeBne+PbNM9JTtN7cirTiwaCpD
TUVt5Kxd6dQdsI1QeHRnPGZQD5pwn6OmLEumlOhEdRPeZ80s3+bnj6irLF/26d4JZbCyuyLxAIJ4
hf+ry0NVXmg2vOysIZb5DffBj8ssSHb5uH6OQg527phJUgORK6vmpRdqXOXQmV4Q6oYiwMCFHnpZ
1Kpv5b2lAfOIOGbSheF29oqyYG9LBiXwUxVHAtpgAyPCZfM5n0utT63fcrVjMhHczOfynx0oP691
9ZwqDgIGieninQVm4qLfjU3wrY53BXZyS4Ky4gLNEUbsS4ekG9saWXz7J50INNV7P75TnaWHkne5
y4iOrhHqocLou6uV1Y1L/veQjiHjAgN5Ux+nzmoEM0rZ393PCyp9DaowHnqLA05icOSsH87dEzuU
kH/ZrNR69HsRJ2Web/KiR5sdvo7gBusnN8sEXcpBnirUOJm2HpLbq4JdHXTiYjqTaTSjvqzzu/iS
dExQyZL91/HqOUHeMU3JsS1sAa4TgfcOIrO2T88o9WzcLbAixjK0PBmczPIrnVPcHYCIRATVL3Wj
D1qVKeD3quOOwHOMmZJsC1JoWVBYmn4qPa1Xwe0BvP28bgWg4x3hH7OmBSfXSe6/ZADcInmOwTX5
X5YjmYZHNsIlDEzgtpPoQ0dhs9noqH5FpdVIfYO2am4cFK7iRZD8zBAUTMk/7ioZjea/d7zQZjyn
1AzCRoTeDXLQYoInj6k7RtRyASkBB9MVAG7yfOE59aP1zxQHbzAmZqjEkjavoxGwpQ26DjB9TjK3
VIRNN+duy7ugBBudNru6b3fg4gpmN7bP2x0gcUrYuP54fw1vAkTWNyXCGVGENQGmzWXeCgvPmqeS
A8ULAQw3Qddr7XFyu3ikCdJHrg0hPLaAg5f71JvepUJ2fp3zXJk9+a2iJzyJ6R1xpr3mXKlwamGM
xIzrhSGmL2ItVY3tWPcUeueul/4W7pZ+tYrdBMd/6gtxp+wHwuQVOsrSQk3ojW/R8BzZpF81wc2e
7IyP7tVsjirDTdk5xBlNaOnwQ+wnZgVCiabUwUodQq8For8vD0XpLnX2TQF1V1Wc4XWYt00MEWK5
x1UzVEvu4xdFzHtLCCsPPjp6L1hJAQRMThtZI5P/D+efc1E16jXK+c+zSV3SA30xpKrTT4W5yJvg
FWeuJtRDMZ5oyy0GELhjqawRm8ALZwyvHTk20gz+xaoXqzRVg4npzAIRN4Ku9okYUbu3RYb7sV+B
HcJ2P8FqJ8ky7EICr1XL+JkMTkHaFoCMa0Yqyw60dHN8eenca7YGVZ8rgM6w6k/O4b5+4gDzctnR
FviK5yCnB9YkfApDk1P6ZIgNcknxfp80sP/g6RURvebpwNri+qfWVrwZpoRcWg5pE4TdqBovEf/h
6t5X2IkYiIWzdRQfQ7nDSd+m6LWN3Vb9A/VBHoJXFtBmI9oeKnSKT4ZZrCyr7Xnn2hoOpRUgrgCH
uO3hil3wHBptst2a6oiOjdJfO2KqoDNcEHVwFTvxkC9pmAgObEU3VqNCL2HbiLCt3OlC5gBMmI0s
hVlIINAaUb3I8aw5OG69y7KHl6td7MB3X4SS5bAWrQYZJjrbH1yxcC6ngh1JxwXIwvs9hsUMvlmL
zgXbTobdmOv14TH6vMhf7OffOMO752aDfWg/R7eilm1JMU9UibbMije0TXPXi6D0perCWfl39brB
u/SPKuvugqLUnUPiBp6kAj78Ah9kNFAV1X6/yh9D5CWovumWIIm0kc1dKIxVT5uhxoALqkq+SV1+
zJDtZnaXNWjQXV4LVdZSrdzk3dPoiYQjUn/3oowUB8bLNcwZMwq1Gr3zUFAnjGIp0bKAc3wltqyk
HqgAL/FrJR8p1hIY2Xd9GE3vtDxaifMTz2wvpwiFfFMET8FPKiXXvy6tbM4P8ICBC5neQbJj3RAL
saiYdhISvdto9qUYtmVUbjEMAXkaDoEdKnDiW6MrcU9QJmVSAIMGeqsGO5bSa6+gYtrD8P553NkZ
zhGd2201D5oQonOb5KEoNA22d9K/nhYcbLQ7tuX/Qbbur4rIfCDVXhxlCz1q0uFiLBRVvWmd4KIC
HuWWiCh0tSJ1PdcDEYHzdVzfnxoYgSC/XJNjeEE0xIWbmkW2NUNmZajZ9q2uzoVe3SvWNNxvqYyj
8E15pTX4hcITow6fDXWohbYfzvq67IKmD8HN8K2KCMSM5uNXgjkx3TbM5hyrqCa7mCr6tElSJzvk
Bn9mJpyc+lpmKHLa1K02SfhFr+RJpk1wM1C14XqGyhG3qltQhcM5LyetW1RaLFIwX99FYWthzgmB
OCQ0OMjCTvuQVQ6AbGgGvyxEW4ci1XmZqP/P2tugipUWJkYWkRYBrUva4l105Eg6L04jixj0wz4f
QmO0j78ci1hc0hhz5DX8qRbHwA4iLCfCZD+tp8BFm9GJDHVBZHWdzv5IwXhrK/QrQnywVokw1tqM
m18QqPTMgJ0nM3noEJQ14xR2T3E+aq52w0sYPbmF7OW8P3rWhfrSNCzFKQdYRfRS/4cCvV0taBTL
V7CNBTx8boLunLdf3Gz7cOBBv/AIQ3wutawfR/1DYqSA0QygHTSCTKXDBmpmMHha9K6qbRAiG57h
c3yHffIRpZ2PTPTr2FwDYUHx9znUE4LogP7xyJGINs+ojKgUFXx0Aq2w7mQrMKZkNsoqMJYR5ntL
Gkk/+Ynoar/TJSYsmNnRMtRk1kWx9GSG4wj9aavXUjMc63Xb4RgdOuLVEDb4xGz0NTM3VwR6waFW
IFZtJ78SFggMmoRcHjxuisesnfJDWpslTIke9hoYAkhAbIiqoki3xLlFQLQdLSEFbyPRv/3IEj8P
ct4MI2ZjC6ralsesjXkTFdZL2O0cDjyozUv8z4Bu5+CIVbzKhciIQlupdvWWeXcQho5X/CS3jPSE
Xmkp+14kk0qqw6yWN9/foQps+jfhqFINAfDmGc2tznIIRVBTKgxUnxXxRBgHjkiDfuCqOxaUf/Rc
WGprhVxk9leOCszvrWLdTn3TstunV7icyBSzgowPcmwkQtCcWvEG858M2nVJDJYtRlVJEyLhTrDn
hlgRgWUBLbV4OeZYrK+g4noSr5ZIQCQQ2T8bSe+IczX5X4gjOZPa68NNEShqRx46L40YZnTZlL4x
9tYYOp3b489TkanMN49xslQwoe2/mqAaoEYvtJysPcNaGHYJPhLkajXUQuOmH+xsh9Ix9TPt043z
8yDZnJwB55fwkVAezJKGp7QtI95DLFF3saOgPLPlwtdWNWnjeOPBVhTCUyczVR4qGIVtKgWjUXf8
3QezTIM+YUGK54dhKURCCsfUu7IHgZDxVuNMMM0IiDwdXVsfZ1EjdbOs/5u8WqMABAsJJ75WU9Q9
ajUB7/15ak+RwOku8Zd16H9J6qMdUG2OOd2CvUe2I9y0CEmLZLtXMNFRSfMt/FJIpttrObKhz3aO
mY/ySHumeh3ujeW0SusfJt00U7WhOdY91k6wjChmCIaqQSw3mPNNt3o4ruJ+UMDCq5VfbmE47CRb
S1zZkPn4BoZuifAhBrt3cMFFQGWFUJ8Y7dywyXYzstGSMsXho1t2vW25NDNwCaDsW03mbq+eDjEz
zkIH1vboslolqGF0P2vvFyuN8h262uN5knAM1/uGYeLNYjSE7EU3ynqe3b2PbBLyHH09Qpj+Mlm4
lWiI/X9sMsfcSehyIycRdEssKmHKOXS78zKh0pL+swefa9UA6f6ufzjJZm6L7CJdDiwCcSkn6QPr
V6PUJe73Z4g0IuuVD9lQgBq8oQWPRIIYyIkmPvV7ym76fKw/dxuhfU46t9q/feJq32hXScKcx/NJ
1yvfdYrVvIDAZJP5KRpdplU8GjJCapQ6H+TLBYKMXjL7lPS8ccVBz+Ey6Qfad44h33lNhc/Nw4T8
BLCIDTLR8yHD7h/zMi6GCq6r+2umjEU94u9y8v2Slw08IcOwrXMx84JL1LU+0+EST2sC9467y1im
ySutVRBm7gjAL++W8FKr/i8PPjXpq71vgnOL7DG9wrb7haEtHXEbC1ycC5G1OSluh6NTc8IgWB1o
MEUsu0Dn6Xlxyb9enL1nDoNWTNELEkjSagBsqKLpQInvY5Gt4cKgwge83upnyHDc+A880pRPBhkQ
pFaLM6mqmPG2WUkB9pUtbNN1+YPAA8ifxqsoV3lwLJjwtc51Z9ic05dAOo30TAdUaR6pTwPq2noE
4ZKSW85VnQCcAHpeC3PIAeN758PWx/488kroDsPzpeRriBiy6/60BV9bSdOxU3WDNciLiyIo9BJo
iGZ9WrGd8Ny3UrZK5xaoFlJwG4XFAVhxtwqk5eBFkGE6v7hJS1+GFqyV/q4W4oGnlWq7cruu8D3W
FA4GH0Gc0XxEZ3gXWBL/D77OpQMgtL3CIe1BMowWtq9dTGquTriz/2VR++cOTGnyH5QrvIpiNGti
Lh0HW3Cu4ZvOjnGliHMOaeAlY9hqbDFQy/cVv++kPML+HfRIjPeqrhUyshop7DsGPc/VomDG8fJj
tXW7G/7I948FqakWIYD1D8VJg06QUd7SPym8/u/xeZ5i7T9Qi1io4dlaFAlGCEvCiHgt/d+C9Lwr
Hbnu6cmdJ4ITjLEfk93JGGg5R6a9SCsKg+HMq9VWX2Scs5aUac7iL+yXD4qe3tOeHP9wwaDldibq
Zpk+LovI8feKjI5CVIFtPATcPojUX7mJjku2XHVtwL+Ar87bKpuPqiQ3ELI043KHcmevaVXwDfjf
A9Hs2rWPpf+gQC3wStqaWV20ctKYDsCAjsgANdFfxsLcxIf4hCHs8EasnzEnuawDQQ3fk7msEHoS
wOhgXNN/xlnfqlVC5G3I+yvhDxK2SRRKYTu/o1D1i/S9HhBlcSQRmJp2PEgTREPnEezCcms+0kqu
OYzYGmZ4MJN/JVE51KNRIwlQ0Mwr9NmaFPx9L1WdQ1enzvNg4uhqkyT7ZRaOY76KeZ1txTQQzmAt
flEANvN/e5XScetM+D8wafxlbrYs+PqG1xARhO/uXRr8GdKAXJC5O0Z8j7Y5GQKSa3f0Kq2lpjRw
P+1G1bCco+/PBh3iaib7C/zlPWHr6sfxBbZJ/EEeiELMA7Wt+lXgfHkfzawH0OsrSYMoQni4/kUY
U7391+rFbaNsvCylg7Td/SaiZnmB07U6HXz4S/CFoCf+eLNuA5PUzX+La/A0F7frTIUb08KZkLxE
PxaBMSFBjDZATtNUZk3boLYvetvkExegPDaOu7kFdH6hi+felBBBxLLbSvkv9IH3zpL4OReCWJGg
pujDiqZsgSKH56/FmW3Nb4EJ0cIo8a8Xh4zMGfN2xmjQR6J8IzjBUl3OGWEspAaYwySJLLuWnm5o
L4Rk4pZHlydmFMl5rnvbANA4ByqpPGsS2FKnEXrQe2wznYoM+KIU/4+XmPgNeEjSPuQjv/Inh1C5
uiLVp3AzIvcm6FNMZUllRs50KS+iwUHWsjcssyT99LlpP6yIY07bn1SrA+87E/eQYCHGhP5sdGi1
YsuFTt3QuyShKj888mOUO7Jh24g6MVZNaIxyEAlJz6XckeEyyfQrTwFRza97TEbLM1Pe2R6c8YbA
+YP3ExxcirIhhy5Z012fqlJzCgwaVM1tIi4KHpL9VuN4jyHqhTPba6bmpjsi98THynoxi/7s/8W9
Vf2dXKeZ1cV1hXZuFbA1tbDxHXAHbjrVlnmlM2VFrywY0SyybZ/T4Cg1icYasYbE5fOHoGudi8Fk
hLYh9Oei/zZtrkxpIQtA9QYTRWK0ZxBAinuthjLHZUt+cSHjtoqKWD16fkC5WSgxjdkzuLfudUlK
V1MIuGmDVwTnwbpMrMCjKp/iq/L+5pLi6AbufFQNuD+8bqKhlGSYdzrn2a0EttaxK4go2KyKfJ+j
giLzxftFock0pdbWVRUp3+Jxv5ClK6LvgTLuuZdSG2KXufdzzqFYMLr9GwXapgu6c9rM8tllQi/d
CkUoexlrCCxBsa4SRNmCXT3D4Ni1Ks0PetLjkU6L7sBbxNUZ8MZlbmcO+SZAJ42fIWr31JKZpg77
jGLm70VtZuAv+vrnMxggRm//WGz3vTwknlmRJ5aL7tUuBetnA93nRQ9L/D2cxB66eIEy/WJV+gdg
V1NRT4Zax1elu4ruUVfLpyEUsuSkHg4t3vqq5uiM2Uke4g0yxfNe7gcXqQt+Y3WruDcp2vADuPvg
OOd7zf9BY3bwrvUVbQohqXmnrIjyC5+kP9PQWR2pXDqS5CKFeQn2UgSYDQ3mwMFP1Rtz7rAn2yzD
+cXsAEjxQp80K6sgEBskFPi1jDvl1PtQIq3N13aDE3AdJIZMhe1F7mg1Txv7LngFPu1XdLI4RFHO
qh5kxrnjvpZB7U7dvQCW4on9F2Wz2o+ZStu9LxOOMsv09JtGzZibj+DiuYb5zz6IMZrFIDOXtrpV
y4fCc8SnLaY3QkQVqUL6eGw7x/6o507+fYcaAZeWzJf7fnKnsxJebdgDprFQKWkl8APqhw/MJupN
NR+fWC1BSLPS6KMdiY52e1N6/rx9+Kiwm4LK9+TUFE2j4bq3TjSgYMbc4iiEasV7bHN3+egcsnS7
S/A/eu4oedW2NkEV5ndz/wxNkKg8OgiZKhpgIEJh4zyZL4FdAhCmDiXJuGFwc0hy8H1p/oDJA0GH
0Woua3wIPIw4wk7ZYkGrnpqhz9g7TbafA8GdiRUaXGeKhtth93tfWrlocItpW8gPibohQv/SwCiq
UkwyGbxx/lyUqBW481pZYPZELsNtdNXh6BwYFcVKsyRfAmBHUZP+dVkm8MQmfFKfHIyCpDF4tsXt
gYW6cKHT71a07fRyQT6P+LJWMVkkVVJ92BXXnFWvzyOa/ZxvMI69yVQsc9r+1KyP1wN1cFrSd0Fb
FR0MZLooH9XjMoImadCQwyBsGY4ZXdeELeYKugfmdENrazur7lbcj15njK97VyPyxLjW1J/mMsZy
Jq/PbeUQ/9B++R4KbWrRD6dxEmjQd+quABVel1jy9s2z69wYrFiRQNnX0l6QenEPKM/vACGc+ZAK
LaDUgRZXcLXBkxWwDM6nVb9AGdBDMnQUqbEPEEvsl0O3ltRup7fMpRDTIfVaL8UgKx95MIu8n4Eu
6q3iYFW1HexpRXTraHC3MgSVbst/AC3C37DlQJhKB1mqyKYwySG2FvmtlfXWeYU2pbYmQlSToLYQ
U91VCS/mCsrxeSDnNo0oA/zwYWM1zQwiXyIENyAJ3SYmi74cpjLubhQu1L9jO5ApmkXifH+XuryJ
2yIPvYT4roDQCWWskfM/MQNMXF07J+j80mHvafDp7TqpsttshfWKesXdEJgDrfgUUILHyFoH5MPd
vBv9o4M9jHbIS6zi7h2cE1fpK3QLUuCHl+Hnn4aaSXvBTtd9nszZsqPShNwiw6f/4vXF8vQQQDZW
B8YCd+66AG174RjgcCJRSRa7JETuV+Nnh9PXfwmnSeceD5KqxbjgejWvo46ZRiuLYSlgJ+5/I7n8
jZEd8pMtOKOYZKFz71pUe3vWbMnk0HWMH7A34ojkfVUyTD+lHZdcGA+cGF3UT92j2qHFv96rQN2u
Sxb1XqAWUgvm2RBZleui4GDhJCmuKnUEWUCV5RTnnpKJMSngyDK0ErFKu6LHKq1hmHCrGGrxAHJQ
soa7Vo6VmONaEjMOr6IHpPhWVuV6mU6BZcXa6g62B7GcyEfzjYTAx0TRHbIZlpfFTQDaqYOUtRs1
q5Jr1qcGvtUG+66nszkt0rZJHXDMQO6fjcKulNb1NYznggxqo0OnMbWrETAeS3tjuYV0AmKGUjJx
7jk5Vd+y8Vlnz28/pnEEIaZXmIqSMcg+n1Enh5oBP74CNpI9HeKPQhnl0StNHjt9MqfNPVQSmZlo
PPS9mXcoFxRd4V4u8ZsdDBiTbaOSdOVmshPQ1rcLLcVU2Mec2gcJqybmhqfR2SyeF9FvC8e9K8ch
YAlVQJbI2lYBHm6iqi+jbTESsJaeFg3mjTd1Jkp+NY4bLsksM0BFxnNXFJTu/zk9KVxZkuzksT4w
DZTvDh4AQgV5TsFZ3cUZaB9r02MXh3Btlgi+cq8eUeg1wFjZvaFIpuShUhzDb17RZp8w4ulYvrF7
4ldT2oQ0FZVOH1vu8YOkKhHB2HlOMCIzvxbuRd3kG2+EgMaY7c/pTRYpmeGALkR15giarZs+0Jz/
E70ZPd8G/Pk2/Ns/cQU7fuh+A40PSMqJuozZSBcrgmoDd/3VQ7n2QDNlhhUqQbuZh0F64SHPEY3Q
uAmQy0ePcqkkeEm3dza9l4va2FdnxF396N4bC5vFfQNXr6Q+3KX9BSg2uyko19vbCaZwaJSjZvDp
40PqavrlD453XmuQQgTuVa2qG/iKcY6Cp0PQSEJxfTy9RDoCaySwmBxAObZcbVxs5A5Ken3HCsiZ
GE8E0gtd9eG7RrBmv4OpVe5T3YlwGKhJH1xH9T+3q9pnE44EEfOcF1gIvLEdobw6hdQ0tr0lPHe+
EwPUvfZva9s6HMKceO4N/W7R9Gp5A5/f0lDduI93mwoqsHOPmMNtCSu43HFsQPS63YNu8MIfQ12Y
gM5qHdx3icAqc1zCS9hTTBsd6WA2JJvXgVHbfdAYrzHHQI9R7fSiwcnTckx9koo29IQGFcvH70GY
h9196INxMkaGwIhh8FelsdSuTDpF024DAbzi4NsUVn3lfhR/+CYxn+p1DhvK7VienpcmoxSC3Kyb
Up+gcAB0Kb5fY9bKU93X+ExqvepdZJxId91viDb1yzdxi6/G5VXeG1chJ5wA/+1DucTZyexHmxa8
wP4O93/DMXd+ItgXqzqlDjrOcjy+f0w+589roWMG9qq1RjbAKiecC6nrUXAv3i8rA/a0LMB8r70Z
ZWbWAxslDlVpAD/ADldZlv5xLpcAuw1fhBtdF4AP70HzH4iXwYgSRCNA4e7Gop2/eRogEz6kPoJ+
fPePlxyeJbWDG0ZT5uEsJwCOEMJ1icHNYkv4dEJJSAYg+bST7K9BvUrxVzwvnZK9kzSWCjB2eOhS
ew7MvuuIBMZgFpH/GK2D5WEG3iwFVaeQ7lDSwucLM9zm8A6PJiXiR2TDfRJ2teabEv6/D9mWzrMW
YSgj9nV2v5W2PzUZZQPKvec295shmuQJ/w04EyDXCFJycOMo+gapQ95TXF/hj3Rjwx7GoYLPm/hK
v4KF1niUWsM9ydPJKvIs1p1sXbL8nX84r1/whNTDnMnUz/pRa3o1JFexOxHu5NRR4EATZJZ/ze+d
qQuZDIvlXVDEv/afXAYKXpDUf94d98TD318bmwfuNqYpVbrj+7qd9GTxg4mG/MNTNPTJnwtDZKQx
rX7E23EldP2ByijgVIpdg+oyKJ65sGgwkBzMCjUZhYhAEtz9gToGTnO8zlk0/iAG2BSLC70worot
4hMws5bfDhYPYl+DAp5qOwcr2vyMb606z4W/ItqV1kiVPpPQekOHdcwbKM23bItI1aDkMeBZO0c2
VThwSRLgntYQXl4+vXgkavuX5ldmSzlJiikL0frlHH695aOw/sDBoUIteYdVoBcNSWBofS5TgiPZ
UpjNCyFUntI1exy2s2YOwg39XN0UZynXuozbmcnS7UFmJwXYX10XJ8L/a2mIpwwPNqaxs/fmQa1/
gsl1Uu/CRSL61dIty24vSDEMP7JgaiQyV0OuATdEpy1crf6whOika1Poe4Si9t0gmsZUye/WWTem
VCzxlpb36oOlorq1m2VPJOggxD27HHY3fB1jx6h2p4JB9nnVnhSy4iRsOayHAu9VvjlCkr6Xxewa
QD96n9BlAk0h341s7xhqiapDqjPbLhqlrzlhro/TkzySv4gsf/JoLFE9HJaHWmx3L7auuW9rZEXy
ZqyWXcdWnNUfSGFFOCO6jMu/tEijJTB1P4mA6FR5rDtn+sNDu/raRMUCaGq19KWQFTV9gwf9MeNo
GktxRZP7GaxS+Jglt2/NkAWlElt3CuB27DT2wqvfKhvvZeY2N4VBHeu9yJB/QzDz1JaW9xn1r3XP
KAXfE7ylN9mH7w/Q/ysa4ry+odIi3ySQLj88d9BufopSuoq+jtZlXo2kE3d2pwJSxXCBVRWEIwzS
le3/g4euZSXeVNL96u+s/YPFSfmdqoBFcKlc8h/qlNmceE7XwdFH3Te13Wj84TmgZNeID+Rp05Fe
30QBrSoHpJqHB8xYnken1LsPA1swM/6f3XQ4ViGtt/tFpmvI1yI9dNCdlK2yTzXk99Cz0gDZClO9
W1mftuQeeoGFBFCHSVWR0PFqdf/okdelPI4cqBCAqczhur9Og74Zno1w9ufFgHtd300EouJK5d+B
N7g/IbeU2ceM9IrIWG5Ptk0ts3/2oxbd9mmDuiZBt2OfiJbKfrXzj9IID6nyW/AWgdauELzj/6hA
N5FQBv4QuNvGpWtFcgWzStyFnSj0AinIrWn8AwUwF/KNLEcITRRku0/5AMYkldM0TXQ3IJvGADDw
SavHk4VxwGxsoERQdTGfx33Mq/etbDzJpHz0R1xED65CrlfOQk2EzKtd6jDqHwhecOwi+8qsIQcD
oTNUp1Gh5v8Hq7Q7k3wWgWJa3Uo+NODem/zzBLpWFAEWLGhkDKTtcDVvL6LCqW0BzyTBXQD2+lcf
Qc1oKXFjSxlUhcXLVeNtzwqmPeHRYtWkJEJUtgx6tuO5+V35lFxulGfRu0FWJ5vJlEebiQZmyH2v
OJ5UwipLslCKixlEeVPkFHm0ryLVz0Q2xXXC1hlMdMLSVl+vTbuN2WVhN5pH+hWQQdcPwGC+Xusb
y8Z/wbANHuADVHA1UJRJi4rsOzcCf/GtfqFOZmYmYMQuOv0zjwV2FdIBw2LcPUheRP5nqUj6xD2R
DXdkOcquYHZwg7jIXncZaOoGAKPslftmeseDcf6Sz8HVP/5nypN8QNRXimppmDigF9CyfbkPp/Fo
z2llRfIO3LKJhzNC6oGGv692sX7DUicoKwCp9sZuK5kRcRGlbETozZ6LHwasVNJ1sLqupxMYzWfD
88WmHWeBAASFRpwBeqy3arD+41azpAr2wuTtt02jkK4y4RJYtpmejnaRM8jgilKIz641SI7xVLO8
kMMDF2kjQCEJENOEMHEtdh/SsYMcS6Fm6rTTL8d2vTvUgrS4fbFnWMqoC/9+QnehoUlxHiVQSBGN
IVYDeeO8vepVOIYmb7OcTy/sut4eZXH2pJoUg4WnH1R2XG9axD9dr20V8m2KfycTe55xnNtDqRM7
VpkvGyeX6rKdeoX7bbNJKb1a4uWQSMb0jmmYOIoT+rT99cf4gwJLVFyGD8Iwchmj16O1ujH6CYKP
zYEpstRTnv1GIEWaRkSLN5x6g154P3LNg6KtkrJIc0dgYalbPawvbkhthd+AgTtNZyHC64ynyAgn
bWoeoARP1TPL/mkbaFmKNZ0usJh3q1H6c/RiCrOfOmpxCf8x7Ib9B+L9Kg2PugcpsxbrLaWi9rFK
6Hhpu1cjB/C9lNxufQJ5X+jqHaX+c5K+QrD753RAmoz21qHaH6ajo2bFD2w+HbfKXTBLgke37RG6
ZLnszV61HLdAjtVqOcPAUSeUH/jf7ebjLWGR00fzFsm7/GjoSRI6bTBIPt2K206Eu+I8S2uXF8z5
FcO6JZRz/bnf1Zr6ib8rfQZCrqdDKa47SGMJLhIVKWd3J1m6a1bM0PQ+AtGBkNj0ric0SbpBJ0a0
hvZHjoiHqfCbF9Rd7bYoI8fqABP7cmOAGfgkubD4+ddpRsDZf8N2xrohIU+yi7j/n4v5gBVqj0Wb
rZdTlq2OBjpbbaTVwQDN+EAd/EBjFGf1k55bTdCKOz8F1UkCprmHrnq+wA6DiqnlzwMLsH2+4Ce8
jKvPyDas/S8Yfj9HWepIiB5DlYug0aqYYe8Um7a5LdAldTgFDONIMszxUiqxTdQW+lXuzkMaWfIk
hSDeLwyMZ+TbkkuQwMaR6oKbe8Blzuex8ySbU7QpN4p7YJKT9RkY10lW6mXHJa7ghSm/dZcwUtQm
D37zPCDVxrGXz5H5U65s8aFXFO/l1yoseysck8032SG89lOt+XMAy3mLysiSOzzbyAWfENFYfjSD
bjI9c3aujPjZsbdG/IQgfKdCNeudi1vgeplIozuIdjvm8hzPFTHOPqkzqzmB+QGZjnMynNn5rmMu
13aZDCsNwxNRHftv/002l8j7d8Te8Kn/tA9vomQdjmC0xoeo4qyPdPO1etjqh2QX/XBRdw5cX9N0
GSs9o6eO0hh69NOzj396RNujUwaar1JfV1woCdc4anZ8RJM+HgrUpIaZd7ObyWZYS5DmWeNffc9g
uY12z39IRKRPxCb61q6/Ryoc/TZumWn2B5xI6KZtwhXzpogCdu81ntNq/0zNdxgfrmw6wohYyH56
YO76t8eT+A6lCCH0SbilGAKpr/DK7TyfeHVS9jckwQOfhY9yZdijDtlofGNAPiyG4o6BxtDcVE7h
oaAKR+/GI0f7cEJBEzCSLoM8umvUibevRvKktI2Zp7sgz24/SLgffZXu3pWBtHykf4JQaRuFpuji
UiTKFw1KKGblFXq6GnjIGji44ranmOL5SK75G+Tjnavlvf0YNAR+yjBsTd2ZhlQcKcrh6V90vuQU
p5fUMVWjGqW7meULHIToMZ/VhGhtUmcxHXM4nCmhW+3C8rjeHDqWgREHP53MXcgWr608AEdBXDNb
RyrWU5cH/hksHgiBXJJVGGpTsoIA1jnrabDzU/cH3ZRm1m9neHHrdsmeafV0M7g3YRjyJS850E4/
xSEhIHseVGGhB83rLjxbZBzpzPZYRVVw08G9GKBQwT/J1cr1t3HW8OBGJCVDHgM3yI3nBilb5SAR
P9ojmYAhFPys2yD9tFrs1u6x6KkHjReTIWfgk0HVBEo21ceLyxZn3Us7t6na5Dcluxk3RCWDjcjL
gUhJ/I7bAJU9Fe8F/yXJa70lRQG9envPOh7K4swo8oPNRE7M4FMiCGswLz4ttXImaX8BOWw/G7Ow
WpddDHycCCbWjfSLpc+M+wk7lwnDk4ivE9iifEUwe5956sDKzoa/Y9qgGLViBW8A6EQQcnbKR4hp
G33v/etH/mA+7Zx0zHCC1998L4ZAVFas2XdS6AbVrCOF/0HSyaKG1sosiipnciT2pJKxsgnjQJ1K
lyRwT/D/OMUrsSq68bAN1OTrr+T/RiumYR53jKKEZyDUP01nBeVftCCsO5jYG8PdWwjTpZumk9q7
4dMQ2CAKw/93ZAOP8C0g1YVpvB5+iJCMOYPcUsDqbdSByk/kfj5I3pvUYsZdD5pasHQJdY9i37KH
oiAXw1qT3p0IBa3Vv9SlpYXP7pFYUgCRD2TAwJ+b0Cn1qxwMVZNvNeGxFBFGoGsdBeVUnF5VLit7
JdyEN4Kn98rWZ8guJEHIxKlN+ja4MwGBTrLOcDTdnfuUn70/Cj9XEwy3KBMUtt8kJhBY7T+1wDZA
CMOGVkOj0OOhJN0iiJmM2r8vgWCIj7Ef0vJAedOD0Kfr60gYRiabZ7vZkxhcakBTGjYJEAfy63+x
18lPdoamfMIA02aGaRkCx4sqPPodhI+6TP8ZCtk6OMyuj5ezAXGbrbutLeE5BCFOBqfJGQWkCup1
pXlGDLlSpgh5IV0Z4Z2lpXIVD20AQzCg3RKxwLaSiwOy0LEfVJ+TFYblvJ8ABuMz76hxbzn/8ca/
Zkm5TCkJrPWugaEAyWCDu5cO9YhXg5D5zStCQjU1Tcvl/+0mU0zGQlpOjJpg16Y8h/kNiNjAoF9x
sU2vNlflFElYzj298rSURTL7kvbw4sIh0LdEXC5Jvc5bdeeoYzYDcL7oDaAiyIuncfzRgrMhycor
GclFgcjAHYy1x4r3YwlHk5yqtAeABDzZYKQEp2FfmvOrygyX4JYDP8RolKUjH/2P4I5BwttIzTb/
cqSPiZffTr6AMqOYYygrLtjC9KlKaaaoQNDHGb8SarBpqI5oKarjD6BTegGFKpX4m2KjHXtC4me8
sdCJUN8wMxiN8Yz6GlmRBKYvG2BXKd/mUvwXEF3D56Ps90ktZLQNEcxx2vwxv4JVPye4Prr4fKrz
TbO/oUSoPAzRgM7FjXuhNYYnEEMy74bAyeNRC/hTkEnm5zOZeDvK91BMG6yiUlZ92AQ7CHDNeG7x
1+4gEUgYwexUsdHQ63QGckVan2J49poePJYmjThOd8tjn/UjmEHFY/c34kCp6x7T/PTNpPJaxpin
b1/DQmWWzgtRPHCcsBZwIjJrdaY8XqUuU7vQzVbhaRYQ9FwUMEJoBPYLeahEIz5r+1nT/E6snUst
A3F/kHUHBjLuPUsJZiSJD2Qyf9colClEXWGZwuDLOFGz/jvCmMEiIk7sYYPVFnu2rWesPtTuCBcB
YWlmTf71qonSIo2DP/VXWmRwpU5PbHF+wBe+4QqcRy8wGFh3tux0JEF/aNJEbYcPpJiFYu3/8kjr
envnNAe47E4Yuo0dFBmymTIz0lBUVZO8WiLqbJ6ACHCb23bDSlGyTGEGFRZ0lRbx9J0t2D4klwRc
x9vJN+nWy33DjajlJPXuKt3oqdYazwBYXENaUKHJkc6s9habX3JC6VL/yvtMpjY/ngN543s2BTZw
I4FJ8r1jx0cmFnDHWOfB2CRS7r0L7KBA3Q+V9ZRGPWqTAMbbFtGpvQSkP8mnIYabHr2zGaacnBDU
X19RVHi0CPZlXmvyY/dWws5Ji9SXTjGeiwMlJCQ7iy7qEPNmSvaaqsb/y1MEvR4RcdaqV926d36E
sVPF/0fFV+zAEu59314VYzAJ0Jm0MXyqRb2RfFp+D0ibtPIEkCL/EgXiChb2+yh+iZmsa1wkFo8E
1uzZE1S0wzyBfceK8qZ08tpsuK5gZs1hCoH5RRMa+0dQFki5AF/myMHqKYFgf3kThjvTaV4ri4GR
p7DyPz/6freFXiBQ1F7Zcc0OroV9GT/74XrxdOw76rV/U+L0PMQzH1lwSRUWzbsNNG+lAfQe6J0r
9RYpku2JhFfJ8HGnwxEmgg+wPndXFU/0JQ9wv0nBZXA67u2VmiyTDBmzWGbTNjDPFqREsYNvYrNJ
/n9fgTzHjgNUm2fUKhth//uahSridnfWL6zsXGb+zPxRXzrraPPwgSJkAxx1rtUlht5pPwxskWtd
wTzTfbhuFEeBbEzkr1QJgB9Zyoy8d1fzMZ7k4OwehjtaC5kXG+weoWVrzCYOcTG/627bG5QWY+Vw
OCksvI3W6YOc8rv/3qNAGj2dCZp5UyJNqvya8luo+on+4NWPRUlVRMp2/4tYa/u+YQLGVbFm4VrR
xAm3fBiyRov/nH5bQuouyez+FU2ImlNUZsJekoIpkGk1JBe+fSaVaAEMvEdd22BsvqCImHLDeCt2
/x9JQZT9scSqToqxjAtBvbfZCi0vfNqcnuV0pg9tusVjUj7UiCG/UEaQsLbF4fW95D+D14W10Fnl
ngUvSQ6LzOIlb8sO26aP7rxNgNLFFZxtuKq6HNep1j5RNROqgO7vADFCa5l99NyP5wOvg2obX1fG
phkqvoaM04UEG0JowO0rnKR0qTCZT3+JD2Vx8DH+DmuuUMvAB9RGlr1naM4HkYf4SH8nlgRvoV0O
LrDQx66gxdFfCGnJiYVt8S8wgyQGNGqY3zdvlTG+Ro99HIPcbDcpf5k7t6eCayshBr+gHdwFgrnp
3cnZ/vgXbEPSk0waEiu//7Pwbd9PCrMiEiE96pSYdXOo8w7J4WgCYBNwxTsmixFM7lI/Au3u67lw
S2W6ZCUwTaBb1XtTqsaJNvK7eE+9XANxCK6U3VQWCcRtjVruh9k3iDhgqmCNRapwwjXpdcywlSyP
L85cm6+QynuC/EnpVnp6vyoni1AveYiV5hJPFxj04+rm+GOc7XlGNqILx+K3WskUZ5iGpEkaFUfG
mTPcNatGJD6R4TjYfXXR4pG2ahlkG9QYIIbpxgGuxDtI3vqCMVeKgoZoSA0g6imu3FLKzvxDVLpz
i3rWEpD7x9tP/8o1UtS2rx/IobEvtEuFQdkHgfavsgywR1xEHGOW3NZ6WGjG468vEUeezp4CSG9x
O6AkSERYrGXtWGPl09Ksc1GqrFjbnLjGpzBY6x56C5g2x94ao+xIi16kI8xltZ6N7SdKGW88zS8/
dzNi7eaeIUvN1qFur4jY+yzBsLlAoVITao7R9W/fuz6Abcfouh3LyW457C6jq0s67eG/HPDZs1c5
z6EJBthaojlnafQy7UiqZA4UO+ngyuYT62JC/zux4MqoXI/rOV2VbUQvzHLFRriw3+0s93pLwx2j
5a/cZz2eBtcfDrYy3a6j8RGoaPKH6Q9qPhd0JSFnlP4AWXYmMdYySpwfzT51xemnIi2m9WQu6JZZ
KaQIwMMuhE87fCYhy6tVfp/4zkyP85RC+397adoF/BbQBw40DPp6mZzJxz3NBOtxSDakkx1Tmxh7
5J0eYPIgRV+z8B79nuTkzXrxd8JsbMCo0pi+J63s10fpYDnJ8VdKxRwioURdPxoYTsGlyhJRlyeC
FTFemgJ9qcD3OyL1jYggr6nbpcsB8yvzLK+N9l2ekeV9yJadTdKklRN7B/23NlXqzxt4HUePnpZQ
BEGCGhDhE1LznSEbajp6RTKrEFN/brgZ9fUhhro7+LogSA9ACSUwHacXclsabLwyVDU0bEG0fmcb
DZ1pv0dUhUDO5jI/Rypz7b2AsNfxRiKHDVewIh87A6czMJkQwCoc6fDpm9fi4JDf33u8/1RDr3Ml
/1OyoYCTyI5ICezPHW1lsYR8qSL64tg6D/h+8Y0UusTmAU1nnoaBJ7Pgi4RIgbYHrePqaFsI3msl
0xj3NXhBrY8/4fpRZUPA3AAZ2Qpse+P3FZLMrChQjdL/quz8NuQCismFdLc/vAquuUT+uKDGC8hh
p+ZXQB0ABLGlPfWwdWj5EinUNg/kX7nVAZBdWlcoOmTdetZqLCLGCVQi/bVwUlSaUjPUorWyjMY/
2uHJCiVlRMtVnbs4D01KwFOQ6xET1DnaFe0oosMMmd7OFqmtCep69HwfK2HpH5HdEDqftKfQ+mau
WNEXRZ9KErV+f4aQ9uhrSTpn6jhP1ZFkZH0ld/7l5iDc1paWF1rd03OVSXt1cRhalS0MYGHocjqm
7eY+AWcoh3z3nOtdfGSFe/6+BWIw72j5pNbvvUeozVfMoevy7cBIa9pK7yyhOXmr9aRLxC8aDnTU
fyEe5PiwrpUkea5C2t7QgyBhBdjI/hV8S3m1kCz3Uyn7isTh1GgmOaESw3xFVk8RaBkXF59fDDnw
VfOZPB7Z83GVCf2wB0gN2wKuenzNpkbv7yxoP7Jrj4Qi3FThOBQS53VgPoc64lQTcWCB208n3jaC
rBwdMjspDMdKZxq8VURpifahWDmt2QnzMzK8akKeYqFSulWv7C3aqf6FvvD/+/sDouSDyVk1tGTq
YRM9YkFYLqb+sqDjX/kvfiFSTRBeTnqbyG5E2vET/q7+RlbRVrA3WDbmzi2N+ztj8aeDbI7TAveo
ylUbzgc8+Zy/ApDcw0PpExjh/PvgZxBrt6QFx8c98t0/jI+Om/D2WSyEh1pndJl2AmdazV9MITJW
wXYTOLkzDO7UhMtowenTLY/ymGK2VOMGVm/v2jKnOqzelPWLU7RvIaV7NpAX0wWP2h08p76W0AgK
xP3exxDOe06LMOgOqFi+T+M3NaYsV9LBS5ZcrF6NzO/PqGuwT5gzjJJOYTPs6G8r7bE3Gn45uZAS
mk+X7A+7cnCvNBos8hAgaDXM3ptMujDIfHwnjo/S2AZeUm7j0pTk6R1XH8USdcZqXoMcd6LxVJSU
7jYC0rVeBNiCbC0sFahEO0/Suh1S4A2/BsfM07uwgcqv0R0MdlTr+Rtr8ZxFxv/VvwKvWnYIY+3/
70Zmz5YuxkTkhJMNvztGeNj1xTFoT0B8soW9CujE5arhQzef5fPkjcYhRL1XlZrwtCvJBdh3c0zd
lQnKk7rcD6MxhowaakjUrBs1xw1P3HEkp2MPd9ksKbAUp+lE+EJzA0O26vh9YFjwlsfTytDXm9fI
Vwy8shKddyjAz8wLootG+5ImirsghRu96VodK74q/SBTrd2cgZp/pu+d8gXQJ+189K0j0psU3RgW
auGUT5qtx8/UWRYth211UuCNgaIDx+osY50XX0GPqR7xHeURh27+vkD5gb+cYXAvgCjYqMKUfLgZ
sI87S+lPxB2Ue7WwIxEMnZG6FKDtvGOpkuBPtgy3bsr/hWn6KU5wgKKQw3XcZD07Cgt7S7j9+viI
FHbCMiKx6b6zg5b89ri/yQ2J1boCAd8gFw6MIBIiGx3RN88vjEXuZTWN6u4BuZoIo6S3UJ0u2qJe
J0LdXADiyQH9g3AKVCprkmuDJG018eEeak5tZ0QDXGivqopIRlwjaeHIa0yPgp5S1911BBo6OY1s
22mKCaq4Qc7rO6v9z3nONx38MyfQSRSr6XEvohYyJVt3Zw6kdIflld4S8cKhfgN89Io38ffQDxMX
zAbHkf6uhSdWXEV6oNV7/0tkWED27/1WS+WWKSQHrfM6gERmal61vhLRYrWKXkg5tuCmlDfx6dq2
TZWyhEOZ6d0nkGuDeDbTl2KsYtBtDA6vxrJEI6cXyCqwvNrM5TBUtdvE3DUFOVTgJAburRwW06BB
6TF+TTszBMmhqIM7IlvLMBGTUbsf1kONScWI5BER3BWMupvnEt0rO9E54b+7azjEpPs/u69uJgiE
CUe45bzSagq2kinbxByL8IPE606VP84/d/1CTGKKq4DY59+ZLTTGTkM+gHDvoJXjw/eLA1Xaxts5
agC+iF4g7LhRotwC+5Yf4+YDnzAg+p78xok9+RiYygSacYI2A0Bht6K3PSmecVXar7OFSqWcTzpV
ScAAzM/P3fQXrqC16xk7k/2KBiOvQ7SPAPZzwBx6Et0Pj7NybNlVxcAx5jDOZ4wOd5v4wohJE+6m
MUGVgS42rvFVnx2dy291z7vZ85Vey3ilFNuOY2jB9bk/Dsy0Tdn3mcbmaNt+IXPlxWDJ0DONbCnJ
oDwT5H9hPe60tsnu2B7E7N1hF1G0sB/UsTYXX1eXOd24lNE9MDEeLBOGglQsD7qD71SsY3+hfH/Q
R9dmPZMJvBsgUjV4W6T5VAIt08wV4/a5BddIctWajb7VUPcnn7qfEosupl9rxvNZqLwA8jDEGKhq
H3mlRZclEQq1rPJgMxgTFlmfbG08jML67k6KsVKlCBbisqEZsS43R3ByGSCbMXmrdO8cUZkihBKj
7A9FcTWa7bcpYnlx9fpOyF6chzLnn5vFVCk3nrXUs6yKUTprf2VDmbQ1jC0P4/nS84imKwb9PGT1
alOE1jFi7+2SUHZB22LmVZRTi1pFCH5MkZcdxlSXthZjkJ5vG2gjN3FGcYBtq6hjWusoi+wOEO/i
rI5msffjBylFaDEAIya27Gn7fb5AiffDBggA0E2Z3ZZm/VokjWZ2DG+iX+RU0BVjlP6Kc/D3r2aP
VZNMXiygzgH3k9SuiYy52UtA3O1ogwDog3B2pULdzhR+Vbvfe3IzRFwdODLX3NbvAjVZ3CLvTLt7
txgw5ruxvEC09rpA0Kc3P9g70z0bmixPq3MSwQXoV/FvURAR7X5YwvgApvvZZKHVwY05x08sR6VS
VzM2xa5vA1/LeIPWZm706X3FoKdXlo/s1AYUad93XNYpDcUENpcGX/E0Ltr/+InDK5RzsHyXpWWU
AqAYJfldaUXZTmDQJmbOBJDBIJImic7npRFRze/A0xwLUo536uodzTM3lDt5tzyTt8n0nHeJ4TiG
Z4Fvgc3z0CN+7x+pIEotjhabclDRuLRPzN+DOi/GMGf8UlmqMv9JQ0K6+5sU3/CPDgasb910rPdR
4KWWcaDIfLEeD3EW05Mh0RcaZYBAnStvK7JWfchtzGOZDvLi7zQb0Bk+LHTRDEEBuUxGrSgf0TRO
8cuRnjrAobzhX6ZevAV3/pBpfsIGoxvnJPWFaMErwknTeYXNXfzmYjOoALqghB/h/o6xlzTjOWDG
H716nEe7Zme0jb+nWDZ3VSQyrib9wHa8GzLvhdavuPCiP7MM4PiMMx2Dtf6SP2IZUgGl4tGdc/sp
ylmPAs8DWzbJ0a1TG2zcXtElfb3kfNI85V7rDEfulMGO6f1AkF9wY1NcKle+U9++aDyEtniZDmwh
b/cnICYJ3IUaNbnCgp+8jm56G+QIHSaNyf3vOHb/bIKo4L+A1dCaXmm7oPBDDLxiJw2ASdahU6WD
xP6vxamGZEg+qRcCZSp4e9O1Eim7k78Mq/6REaWJRJGPiyBmORDgFb3luHN8gA7qlyIY2fc48zGT
GytJVlxuOMLoU1Nt/JdlD5Be2Nfr3YYWqNtC5jl7cbzOxDcLPFVqh7gTcoam+u4L3FZj/1Aboxy3
/5KHS4zlHLg9aVP8tt3jBxAI+b9wwUzW/OzpMBRSj4SlwG8zs5ZDJEtULxNZ6Cwov/K/te3tD8qI
eLRMJOp0RIjT0gyi0zYoVJdNnpwxYppv/u/9sUlRGKfMsFZA5LXcQMOW3nRP2POXhy7qsYMWqhwL
WohhOj1HXGuDeR8NAjiyF3r6G4N8hKPZ2P0izhhhLdpLA/B2/IwVj4myxUT/NFq/UtSP57WxLnAl
zC7OJkFv0JOlnzBJtP6HJrYTKRFE6VjoPZbSegATf3UG2c6Q1b1c8lUDFBRcTN92dLUvjcJ1Ordk
3ZbUyYrUb3OYdzUAaueczTYifYSfJdpMrfrt9CHJbqk5Qi33COw8KeIb88spOpKOyh6yLYjpuZhk
AWn0/Iyd8cVQ2Ly9WuKu9Pal1gQL2F5c7vrbqRtkLzrK1nVj6MWhUJnMciADri4xhJh1t2Ix4p96
yiHMr1SB1tXap/wJ45bcnD4uHE3Jpthzix+kbwZ/XqTTlD7PMeSdiKjVvKV1cESePrI3nZeHX7je
l3xCrpuCXB4BMzPXfAH7E3ZUdlhhowrzrrS3mGd+SrncSbn4So/YQv+EJTkdnfjmxhOXczpcWYW6
arjJNHLWsPIa+Zk/QmeRSGTpKUS+kKMVC3hAVc+cP5Tqx2TKEnaXClfr05OiPCB5zIsBTQV5DhhT
OX5nMD76nZVUkLZ4hM3XV6JwJViX6k2x2y3HnCQbawsoTD9BuVMli8y+37tP/P4OFw127n9vLMRk
pw2/Gyrd7yE8BgheK5zRjcozAXo5bjOlxUaOaDiFeYBsbpPghLSuHsHKjqxMTzSksd+NYy3QKUdC
uW2ljVZsMJHNsCjXH2pML99SRxZYimBeyaTgxohRZcLyFa4oEOZBwayjQ3TNByMDH1WrwIXOzNh5
Fhhy0YKhl0Q4pNBNyrAhpOF6H489xxel8lg/IHltJX4dw9A7z5q2ZiOTwuBc0lmrx4kw0GGkCbZu
cJn3Tqk2VPch+mz8WdyLfEMq+R0pj5oy0+hd86bMiQB3ELNOjAXVKc6VgU0+cmooTVe7vK4p/3y1
MuDo/xZV2xv+zyM3L/SSiWyXmL3tsKBA9vfiL/0bqSu8CtzP7Gnf6jqc6KIuGOVXWClI8PFaZLiz
sphPxt8RbtpsqQIBmFkrrSmDq0iWomL6zlrKueRn6N9JvqkVNirk2gsVAYZiNidkjkIh0jEFxwrC
hQawOHoxUkWgV6GeoEmEwkDLYd/bcYCRZF8PO/MZBfAeb71S/LnPRgxFXgIavg8pYXiCP5EI2pa/
20HRmobHK3xwwzUswLWLdcFomsOgGFDxZBO3Ir3oxm0sN5xWOsBfPYHzbO8kRa80hM4E86C+XeMd
ql+2Ov1r3k9H+nTTmySMbj9l1wb2Xs1tCjYRHIqF3R3dmLPGf1m83YS56U2JC3l/gT8i+q5CTPvK
Yl3TkYJNaFRDlmrJH0Z63AgNBhljkbJ5s70bX1/1It9AuF335mWC+Pxu+B6zkl4dGb6PNUb0Bi9b
Vntq87bl1SZVq8lRcORtmFDZwzFrpCzSde5/olFW0TMeBpijEziqaaWyr0rHzDcU7ITylAx0jlXC
doBZtoiR7Sl35ceraqBH2ZHyT0NQbu3XPakBBkPE1y+6Allo6ThiMtaXTLTlTm15H+nDoIXtoelw
oRlSgHZxqK6f4+Vd75aYALGHuzcEHPEOQUaXYLDHHPaejGw3epRDf/47zFEIW1klatU4T60wEgiJ
PccJeqUfgfQh73zrNc/5TH5fNj8jPDvBQH/aPi9fvDtdOHstJq9hYxt+gzSSqI35/3Kc6JdL+Lk3
TowtK3q1shqltgcYCygYHHGc6IFh/fHh8bf62c4YcdBGlEhFZ2zQ8MIPSBOObgVJpHygtS0JW220
nPX7kq3oAfPtmQR+j2blaf+8QbDC271XWp3L4Tj8Gv0ZmpBsq8lh4UXPlLffu6eYkNxZ/eyZ4ZK4
57YvDZ96FVIg2Oqx4lJhgiBEasj41cCSqXbXT/IBVgQPhl7FOt0xJ61fUT5pKpHMYKo8pCOLILEJ
KhEUrkkRpQLZTbD6a9zrNex5sGxCWHY6bweXcxD8g6F1+zRYb01D4uPaPCS7jGazO6LqcRuSun43
5YRQl8LwOurjNknTiCChj4YHnasoJs9fSPN5j3J+GfazhJfC8N78tPYhXT/9VK7i6qRX0j2M+CGe
YX9lCtjdsmVPjPqvot6O+I30HNLnuQQfFL6S/rBOABnTEwNfjEQKC8QHqxDzVPB99g/AdZ6xQIVX
2a4T9deT6pqrriCUvjwtU1u79EAS9CtzxvYjgFh5inXrn1rlayKW4p4yr7WfgwwX21yw3q39cYaT
wHXhLWo5Mi2qwKO5cYgEZeoKNvJmDCLosvOk459hGsMa4df7L+pElj8VPMectBJo5frB7XhLtudb
1QTyHGFSGzAIgOMpmhA8kZfT7hEmbNQNp0m4XztyvZ+HO5O3gy7/MK/hcSQ2soPXzdRXuWSUEWyB
EYimZ8uzmOwDlv/fU1hpK+QjhV5Eb9CUnlXwKaPO2AuzuIKePOxDyL2DB3kjj0EESxCsiovKD0Y5
Ty9vfNDnMbUkcqqQp9FZeT6ToHwWraIVnHpXnFmPn5uIdibAWN4M6mxgpnRYzCNVj+Qt0LAfIImV
9Myla5H5Zogwh/0Ib0S0/RyzjPm4QKr0P43CvZH/Ru5nkI5+//NprpMkMkiHHpTDVCC60pB40caw
xl7kx2gT0ow06TDij4mfcsA8a+OwqYrG52TarbNlB2l6SoCAGOpE51Bqq9QunhU0PGdk6S0KEGFu
tWQYOJ0cue1INiX77mc/0IddNfLps/4Qw4kiPCp4nWdZMOSZyx3+oYu6XPMVP3d0urFEAJUDyv+c
5VnsjiJ167nrrbuOWg6EVJ6HrUb/EqVuRQ4CxQwvN5R7s30EU8DCH8MdaIQztQFryKyt3i1BwuS6
YB+AzHkgnxII5sp3bSgjZQ1rrTtdkjPfrlY8dZCz0IYIRSQv9eamRBiPfNz84lGF8mPT/blaYOhG
LXgPNTj68ZdjPSSDZGR5oLx2wHAqkE+2pAXRTrfP78B+pGafBiltrbhiMByYkKQjyKxNJKR7ALkC
GYayz12yBlge6iEZPAmN7VBbhj/H2DNfrww1vTWoJcK3f/Vq0LzXThb9S2y4bzZd1X+U9OMJsoZF
pBM+wRdAExUPJ6hylPG/tVa1mk9YvrFwf4cjXlDbKhkr8RgG6kNF7QJFt4mXB1Y/N51YRXjB1htK
vs5m5cavmfvb7BdytcmAwniUO/vdZBy4ORbwCbuHms16DnLFOwXqWrZbmCgIQ9GPGP5jYXqLjGUz
WiEDLMZzAM34pX/VDKnFVgFV6P/GmoEjwo28F+PwG/J9QKvhRCvNqGko+Qem1HHq2DBRyAjx+Y0j
6gnaXEsIMymazVVXJIefs9XGyI24Mg297OgZiBjEF0TexiNk3xJbWbYYMemJjRq8QLoilFKwGzcO
p7iPdU93ofZSLSzZ8pr9ltjq2seWc0Kp30xmqWNQMevpCuDPd9xoWc2AdEV/XGcL8FuRUzI9FYLP
6m1lvsRysrCi50dgkCD2z4YTRiqRNVcr/NHkQwsHBGnjaW1JqcS/Xew1S4GBhITiWc73lVFkJivt
MbuNV9lkn/uGnHZgFxxhJAFvB5iu6qPK53M3cEEwOa2XRVoR+1y+g+vKc+ZlK7CNW37LBY6osJ+S
N4FwiS50B9Fe77iBT6LRpPe8EtuMZ0bk02ADl4J5YnPksMC8fgiqn2u2GFlJ/4zyhLoWd+SJLz/p
5pUyrnafRjnej5wZcxYUcc97o+PwMe3rQQtnzl3QxxthqctZuRVaGJ0Y7ECuDr0yzdE8H2IVzrNA
9WAZlaNL1RLRThPHRPn2dK0hUZ4obt2CzV22LCObxLd5AzXxyzuGehXoibYey78f6nSpa3fyGWyE
+QwrwGR/0Ze8ZoDKZDA3J5UfIXCwt+sNLIiuhBRf2XS8Wz+n3AjW+tIKiX0C0NECZcg1mzfVtToq
K5LeXnYWVX0B46+n356FnVGSffosroAviYC8mjxcQneJYcPLUCav/UPRxbd7kFFm1zU9v50L4fcS
/Rj2w8hPsSFFfWyF11CmDbqxRhqlIvse7DFPcFT2OFwQxQpMKWqG4VrVoOcVa3cfmFFUboAiIIUB
kpCccG3mupB01IAKxx/2ncBB/2PuZ6d62ZtUSOrWAY+jVwDIC9Cik/GOo/W1fvzurezNYTe9Ia+2
1jI1mDBU26u4OBcBSzy2eLizR7m/blQ+cA95GOdcKNWI7BrR0Km2Dz9leZGzgBTUXkaP0GCYBbpy
4f0Evz2pJKackixamjBxjjk4JqB8V1oDgMhj8J06mTHu2bTex6NZ/Xwj8cTNzOgEkUpKu0/Bclhx
pe6GPhco9iSEkRl8TGIfJA2IAMV+xSspuQiw/J327mQoXaySGwWIIo/zme24e6ejnvfSWjQn/Pso
O6w1zYQqosUaw2Zf6UA473WWdYZl5uwfQ6CXF/hap5lm7yHsZlOU0OZXVIMcSw3OxnAw/CPRg5pl
mpnY/Ps6Xbf80NAikxGlZRmdto+Nsf9Qux4aLbjVc3EoGnItkDwipX23yrA8pI/QbWNTuIeAUxFH
srqUFjk8nGZWr9I2EiOQpkzz1+ucDic0LRcz3g2AcGC7JQhBlaEeVa35ETrBUCeVLAlT+5FtV9pu
T4BhPU/+5eBuAOzmi5gqQg3rOY+ELsHIBFsJmHkPtWXPhuRsa7xEYxBjrvSXRuWI75ec0YMs+J19
YOA08UXs+EIG0sTFER54mVaxaHtvVS4DBVOKlaGAzQgeoOHg3onmTMUhro1U16ogIN7oP1SNGRmH
ubU0dA2XD6UcVabVeqqfXMZGH/PW6zGIHtK8BSro2T65sRcjO1eVhih8ICMUWi9jyt+MSzJJi1W5
qeiP4FfLZjZ9Czh3UURglfXy58LXQ6GW6x/K77fQ1t6tJ+UU9V6797O23kiRoNFByexrS3MaPZIp
us56VCZvZhxBWmn7Otj1Rx0YmM4dD06cmSO9UcpViIMgBlo730zfyyc3QpXnLQrGTeAKftb9EbXb
RZvmnGcGuy3J5WSai6KJP4p2PeIEsU09GjFEF+EGcVIWzl+XMPz9GyDj3tkh3WGnxYxPUbJxcgHE
ajvf5VrKQD5giOvHsvKFFubwELkCCM56ii9gRwIBRt9JjUaKTu1adMJgODhd3MugKYK3imNx7aHl
QUb3CrwPz4dld8AxJWcNIxBPtSZNC0ZxOzBKVK0k9Rdq3SajA3j24hZ/DdNukgsmLNMaos9A8c4y
WXSgrANGpKPnE5IPjbl2fIGvN5wnQp3uTBic1S9twGYg7t7OubDU1IgNDcgS3uUgo/8AyxbnTRXw
0fcYdoEOHbMJKG6KzUPVF5zhCk7rCNLmdKa+nzA/Uql5CFqNO+j3e1I9pBmplm/SB4nimiAzvSiL
7PAvhP7iIg7bBnfxoznuKrA9PAIaI4wCQ/5tp3D4VuKFrTCjQSjGePNUuVAmp4CvlKhX6groyZZW
LrlpdFowpDlJ0K4HwqUy9AIZhU642sBcDrTC5Yl92OMh79ZVDsVjoRMUdr5dx8lk9NeV2OUMMgWD
+ksZxib/q1Mgkklg4n0XLROcYU5NOSm4ujujjHA84zXTFeKi+/LjGYPQ3hPFjPJ56xxpMwUUWfCB
YG9HukH9snp0mAi5dHEyk56EN4MU7shGaoH1cwAQ8vuKE0NfosAQgikHpP0FmHxaczREwSRXOemn
S7BiN30xRwXajj9dNwvOJEwsssXj2aaMDkYEWvGW9/Eh7Hgr8ecuwvgl/kbbi7ttmiRGfDm5tnZD
KyUlQrTRrF3u3V/TYVysfHHe5JE1Rr9xJTW60y8CeOS43LDmOVwVgK/pLKy9Z84dXFyulqWsf06f
lodUpSSaZuda8FyMRtx3k3UqLVDpFFa4+S3mbJcm++8Dp/Frp9SniZaI5k8e6NDSDt7b2ykacePi
MIe2vSspbflYWCPiXmuNrPdCBYOw6ghOGFbb4hk35DXLaa621D9wUQvxDnimpom2SdQclHVPOy9g
6EXE0A2n0RUcvtCH/+DedbRAct1QldmsKeWnb/tcmaWcYf7S703iSaH18R39anjdTox716XRCE6y
1DImhCrsOxNMatYMhdqfigNuQ2q47Eg8ceDaFOlERybKLApDCHvxJGkrRbWJj+ShUpHMN0G9cubi
gsDQ8FYoGPFvWxDRmkysQ6Wxx8mdyD5tqYc1UoIPQ6CcYFHyoKANMkaBVv1WVtTZGJlDtCrAaURN
oY1IjA1RDNfQdU71BSRukgStRMwTI1dk++hQbY4VwH8hlkbVSxVoJkvVKlK1Eu99U5HPL9yZqwWz
7ePh7jO8dLrmaWkd33DED9+6bS/l8bvskpSrci7NLsXc2JoL21UC7eJKTqc1unwIW02rrSmhFzm+
FKjwzUyJQLMHDAaAy/htXs0GNAR6DG2123rSbdl13hwEIG+KuIS3QrNbaleHOmPZlfSlKVh+ZazR
9BI4uZlr8yXk9rD7P+97GYaimUh4T+3vMS6Ag4aZ0jV57YFvqQfQ1DNSZClUViWQmQcPBWSy3lUH
29X+amo+fqkD23UJL3qDOoAzNNR5u9JXTzLc9DfS0CfcSoWhz2F5jyOsRRQdUUja6hspdmM/ANwy
KgpKbhgGK+wk6fIVvqt8ua6sAbfZG27qT6pypuCzNwgjO9qS0KYyJA0huzMeXGSzxDdUNrzlizBr
NoABaGE07IGE8KxfE0W8F8CMDPQtUdLpiBrARZFVAfoLc56EAK3X+2qxXJ6XYLwfhGNT+5Z5GqwI
zlnOle++B5rsar+ftKweWnOxYwkwzSY9csYS4PCt0hzYD1l13tMJm5yCbyjaH23eSVG/WbF7WoYh
QilSfvSv+BoOkIV2CUnvmQayCVxC/zN2VtntVhMrSIdHZODzUwrZ9P4VFDlapY9my2MBZVUDRxmO
aES2TDVr5UOIBiuMCujsCg0FNRHXJ66NSGJ4V0iDrZyAz9ZQmz45v5dRTR2NvCsEja9z9FU6dWaI
tEOIK3j46hK+DkXwp5Of9yhKgHW3TuxQdJboxOiYniJaWzxJh7JL51eXi5xfwuMIj0xNpRnvRdsH
ZHLMojBGCBfhQhD6JlXPlF0exe1tXLtcZDLhKOm8hFjQCLpWLrnwsZXQqGy1cULz09azZJc2ticr
D90+droaFuf43/sJ8QVifUAodPSSLiMmMZzpAl1AxuXqxHh2dqvlWLj7LLaxQ6l1lSuJstnF9m/b
FGbSxXvfAv2a+115aGjts/eKr5lkfyYoyHzGBjgSEBlIWDx0vyPSUuiuwjZAW/qpAVbqapj4S7jb
jBtTWNWlOjk0D/5PHB03ckC8fGL3MczDFd3ejuHn8SzV9oMFfW00CV+82zsa7KU1woNx5xFSYWhq
vPIpJZ9qgpkulVwPrJ3TqgJM3ECX3/TV7+bQCNITHbV3IJZYiaZl/Lo9EzPbxxBZVTWex+Ks92az
lo8iq8Q+mc2rSsnSscefs1u2qstGmvU7QrEgJrdJqb1yxQzqSKc6LTo6BED1xWjYJcnhvYIui5v/
sHHkf/OdHun7O2DD1IvftBjw2AmT0AlCrnQCYVBx3TeO2DT5SxOsfTdTbsAQ9MrQvQ6mLKK3NFxs
+mEW9kke2QNwvRtcXu7b2ZPQ7jz86Nt0XgbnbAmaQSDNeYOQCeIsgzCpOHdMGJysgPDJ8HkUUEI5
9K/ngI7FhQIaBvHrdnGNFKBEXf7Umkb1WgcSuSos7ZptHpP6i/Dt6xkW+mCmwt09mDH33fFeL47H
y7CQ0Ns8PZ+UtgrY1ne20SL4Fy6eLy3wp+K1RObeiUSlbNhvw4JEhSJs3FSua15SFzHhg+T8mkNA
OuXncJn6orcnoExe2ZWSw1LqVAeyN2qCiroWVSNlrmYDp/OHPyPXdUJhHfiw80/xzeOXwg7ARf3X
ew27m22/TRktRXj3r83ObRX+LDtBQSs/UZBtKeOSn2SM4dFOQWKYEaht8+Taev9C5v9/Gh+o1wdz
ZdWoJzz25DcdvlfKI9uNuo3G7orkWy+dnf7/GlY7JHBUqnRbR/JTZmm1IR4ycIULtd1xQKfjCamU
XHkQyI2PlR7cuUps8C+/4mMe1cGTn/yKYzywV7/VkbpOXfioWSv6vZnt6SmT/6AItXcI8E7AqVtO
WCIhosCZbSVN9zUTp6ok+KthUlCA6+jzXUvrNNladdhAOPbDz05pwnOwPt89HFFFc3SGR3w7FSO6
R+TakBQ+HZvbIArCFEu90jPZGxDWU5NY7cQE4CHSH4hSskSJwXsoOAqzNh/eY4wZFyEG36jk9pXf
tnH+mwIsnJKOpOu7fUJnIpWQSRwAYg0yNC4H4U3hb4/6axNddDMIJV+lChEJg+8qN53TrWe5gW02
GCU1t83ddtvW0yjZY7awckou0wsX9u+4mKYCMMa0Zing2pt5Dgnma28D7Z7n8aWE0ZZnv8BoezxP
llF3J9XEB9oLUA0Xtx6Jiv49TXsNNsLGrdVZnmeQw0MciKvnveC3GMRVSKD45dL/uDa2DLTyWOUK
afy2HfohAHpVy9tGHdWhbI5lstonk2PQrABdvHC49w37ayfp7GeHHpLSSvbDpR9mPT/JJEVIDccx
vipvoQs6JB34n2yiyiv75UhMjCJIBJzB2/6uQHcA3PbedvqsejI8QM6tQHJFKoW1s3u1l0OprMFQ
tecRGNRQI9jG0bBZVNq8EQxqkDjE58EFD4oF6AtAJCDF0AA6KfSNwslRM0HpelBcvtQbUv7+yjOT
phnZzt+G5zAH3rszHcDlIXDksMnbJzMJJH9QGnqrvRoh6ZLJZYZj+kTcEKXGt1gwH2qS69LkUTaM
llSTfiBR5m4+KTxJEx8qDIPrjZi6N/+zB8NFxSpyezpHg4a58JnMHqLL4nzCdvXhSfNQYEo36wW4
9i47XbpGznyfIE0FCQgPfl4zRkEbO+ij/ZOvsWtUdmM+pgGR4Xe8B1ttBbm3/ph3D7t96b9XpNZR
XqP7rO4QNSaGnJd3EuQY+AR7NFhI/4v2j/2j3KLNco7+daac8sXnlQ1DsGN6U35jf8JpwDn25s/j
1mv04V05YJX8jiguWRdmojqeaMXa31oaGn8nRg8+JR/+zKiMOZZqgjJreAOiT/kl+36LagA+trzx
Eabn/bzIXbrdiu5m7eZDEnGRL/6UbhoZZ/n8PyUnKcJXhKe/fJtARRqy2IZblbXgOKUTbyA23sGx
XKj9JXVSCFoU6lm+hp3Bilw549dcQYflPT0d3fUoj3+N95GjtXL2zDNpKDfoURatQYzd2pRJGcbo
b5bWPC+/Ry5/nuobGWGoEvCs5hT0ucfGUhev6ZedaWlG4ovJyO8yr8G4umNxDSq04jjZDCCOt3Xq
elc8dRM1q73YJJ9S7u+vAAI1Z7uaS/S0csi3lrVdqNJsJe8xajDocOgy4LmQbN4Z6xrWxKZvsxHf
DBfvhZzER2FDTwsauLBQnRl49hJ70Zq+a5MkHfz5OVsmY8/2ocuuWt5xTt1RDKNLo/W6G2MxCFuj
F9PLe5oAzzcgU8dif8FmERe/0DUBk4+05z1q2er2yumYLV30voeoUvN0Hxf9wRRboFltiIHP3OWc
fRKmf/n4DD0wkkeSN10uAOGyNGWAENApDYjt1YrVr2zKxXnSzMQF8lzDg57sN/8XLzbgv6iv9fEK
xuO7QR5VVxFVA5r71g/oV3G4HBdANxXcBNQSd1nb/eQX1YdK6kQMJfjhVuUh5biVl/NRfjeLRU98
64oO6l9b3LFJotH6s9SBpez6EKsF9TIPjEpuIMbMaISeTjwoxx2DWZhHqSrCWyFw8tkmY/r0217n
GnOOJf0tsVzAorZ8a3XUqMWwVAuEeh5Prz6rdh+ae6qDBJt/LXun0dUFJytPbSAHyfXVwgSS89OB
CvuMMYLjGH/tGNPGbPkaa0piAX1/pwdDoqQ/bc14VwLF7je1PcG1/HHBrltCMG2NkIQuSjyD9orM
sjAXeb/m3H5Mw1dXoubt4/RByu8zP34/8TGFYkaTnEhx1Diz/2/kFCY/K1PjVFxwyEqKkCTZbXZJ
HfKUW4WXGfrxYFd2K+YXu72NaXSLifcfUZnhxn/u7MMmyAIWXJ0gZixmcbTYDhZWlf4dEfy8lV5v
vP5rQ0VvvgxwQkn3OOhqfoBHwWe/tSqljXPcVv5buoTJX5iSJRJEARSYkeXrB5k/igvksqS3bGul
dFQgztqQf5o/sruT7kzlszCLrCp77BlkEiat2kGCMc9QfpFCpK5gqyzyzN6fM6/e397zXFvWwvcs
A+Yc1SfLFDCROOoLW/n3BGHROopeic1iznXwnKbvqhszOkf7LZu6oWzDXSuQGCH/tD5wO3hMLs8/
A+OXf70ViHbfoBlH4dJK4Wx4nF74C/ZEBVG3elOVnqYx9YfBYcDpZpgPnWQo/uur2oZvMUHJ3bhV
Qo+4DDwa9LebKbgUjnQnK91BP081qsuTJmSsflQRw/sQ5fcPxeDeIPQCtNwCniSGZFeoO1BWn8Kf
rdrN5Z9GQFTT5t9kOpNTFcBDeJsB4CzOUBBjKrsfDBpKSdXm7EXo1Pa2z5pbZ+aoO1AqpKb0x35S
hAc/a8SG2AfhRXFLXi0gGT6MVjiD1J4ddb4uL6s/EYRhg5/VQvKfIEyKlZiCle31rLFiem7pxDei
FvPfpVmvmcPsI0pV8FNwLbYKntrKBLGOpvGtEb1DQjWU63PO8SA7rTzCuUCrj7F4M6XujnNJI9+s
qJmHDcJm4VghQDu50pTcQaRORU24+GmdmFDo8u90cF5KaYnd1+VXMK6l5XYC+jNV5ITWDeUWIm0f
NhrR+KpLEh7Fko0ilUX9LFe+zRuuvIEPY0FnWMqcUBHmS1shOsbY5GQl+NWdK9OuPyMMRL9hHJUE
H9tYYPfW7beB1GBcybDLSF68E2zLh0mtVeQr7mAFml+zonLmqudwB+FrirSq09XsjVRKniWsL9HA
3qz2nuk93/5nTG5Lh+rGvC0/8aQKQqI9XkHOtR1OLEVGEkXWCpHV6MSHhZqNsuL2NKlEqnEfRjAd
c/VY06OmY17SCtluiCER6PMzVu16BcXH0sGiBoFhbqSb7hXIMfka+E/EEcB2UISGTuLx03crgpGs
k0E2No7vf6c/twWoijO5NdkmKAnIYD5cz4TSZ6jKfDiz6uOerVq3tCO1LE8j2/nrX5ilEo52+bdi
gPCr/b/+Iqhi5ESMGsLT/XAhvIQ9lMVpdDC7CnaGAkNQY3UFzU32DBZ5qpvfHaEar7LzrAiYDh1p
n9Rw5nErzLypOqh53NKkgXs2EDZRl3HtZ2FETo7xbIgcZpMWYNe2CQRKKveY+4jiQQGfOSJqNTn3
ZNxJX1r/Y1YmgzO0N7t8n2KUH3g4RV9pEgzHS1jSUfm9x9frVXLbvVdQYI9KmKOfP9qPyZ5EAMKv
7YGlEzKgxJRgnk+ziXbjMDOT9wyBkHJOufL28Xl24a1OklrO3XqEC7fpoE30g5m7FA/LvhinVnyn
e1PHW+3Vg8+aDyaOdMGN9ooFDpquiU98YboNHWsRJqzGhFioK+7mXgxdcAJ5FGoZ1tU9E3HLZjwV
SBF3FVN16SdhU0gWGyLszx9GMscO/EYCn/2rVCMA4nLCN0QsjWLPHAAD5Hm8Ji3hNG5JvN7PyRen
C/v3A5CIcA/1eQS0fZMYz7vQY5K32891oNX0KjDNb8r1ANRqQyTs1KKB+TbTygQ/WvmWYL8zhgxP
0qtsPvCr4nXJRSe+VL6qtjV6c1KjjYlWuSemzYyOIR3SuPxK1TtHvAhW4O43Y8gQajf80A9+/hR8
RIghMseDBH8n2SkvZE/vTicXy+EQLtgfSOpDOUqTr6zlKfV16CG8cYskDwTI1nOOvzbn8ZTlr0Fm
pHD37FR7dJJzOoDhGgO+bTGE8lA03pW+7UkYL/100DfjCFDrGQx9TnXxMUYDxqHtN6Xpqmjj59+Z
gGRu+wGm6rznNJC5oQpcmwzbVhhGUmpn1x8CvfCb070vHePQrS7UrRl5Olg/cza3mFwxfOWCg3TY
WEg9p0rSOEXwNyEHr+6+Y/sIKbzhdWUOOvHamwpBWXBNPi58PtZFT5BRLWNMnLhRLU/5n8aG/2uX
Jzfbbdzjl99DRTtZ7LeXuzOOXkb3YECqg1B4X0a5lyEExp9HQHfEhBYPV5yKdNnda3Ue2DvJ9OXU
MLsKFHYZFVid3A5MWJNczNS9CaPJfkl29NN3teqzV1b/YrIIqoK+F93dc+VJw/6Mz8sVovLQHVrg
O1nmJ79tkTnoc5wkSCIkko5bv6Ma+dKwezYoH9JCzRJPdkhcTi0v8jFwoCHkJL20lnrPJxIlnQcL
IbbXsz07bv/FYL349bo6CEtQpYF5DMk3AZ60EB9uZ0+v8o2ew9/rAeJszRbz++K8ZVbku19w7Eh0
LfGUdEA+Ug270jmrcO/wRCHlrhI/k03ulLrYUgc9SCycJnlAFrWkbV3afQVf5UJaw0fqZFEZ9nVI
bfw1SlsSVyJhuUFDLlgpqQfkTePqIa8iKBRqVYNgUyCSZBXzRl2UBm6P9oDJj8ogaDCp2hpCzyam
M9A7hbOho6o0/QHeiXmLHB9QhZaPLzVsI/dm7deeoxzeBjxysBd39xlvvnbOcomPawfh/WS4k9ou
XElrbyDO2mHMg1ffwV2c5w3Rj+zCjSaX+YhLMvJikBKV8M5tKhQyg4761gUleeZx2Vgp1f6FHloo
tPCZr9Ma8yKBJnPH3Kdt7yo/DVBOeKQQwdYRP3XTMTUywoPP78E+4rD1+cKjrSKEZ0g+g/tEkc04
VxyULQJcdNRQgRMhVfDHcqnO9RhjFYPX8ts90UJe5sVa3XOTwyHYOjSi1DK9d1RdtVd4CmOLYpFH
j2C32/8H51K1+AIAvZfOo4/iAQT9SU4z144gzUV6UYHxuMZ3WlCyJO6u5lnG/DEp6agTip4KYF3T
0PuOQIZkBFxDL9R217ehIiMphlJKU1wPtHi6iP/9ilE/WMhAuOLyZGLvA05DWt0y6zObSBwN7THv
b6SCZo3a5wO41yauyu3pqF9FXdTdfi27RbsZ3Z4j3juYk3Wf53HsED4h6yhkcpLDWLrFGNv5ACFn
zIAUYl/igH7zk5vOSPXGqVKcCZwOc7V7Kd3glM0sEYoYQ6kdJwx4F4ixRHVkyL7lipE3HlkqlFQI
NZppgdtoOmjrX5OSjM5ygEHgLu5UMRfjYA0aB4Uyl3QdpKBR4sy4j1lakUbETSv5JEo15CtSQqLo
b7ocwMEfnOzu1KGIDCVOyP8EU3Ke8+ewDhCXUnwhtF0nFtfrq6udSUzoBXOZ5weBLaj9qfZViK1p
gmLo0/0q/4awy/GFrBz1AeACR3kyOwqP0Hm4VJ0CGpnoTHfa2mmx7I3duWmjo73dzXWTj4yac3tt
izV4i42dYRMRdwqCJQNrKdjwaQ4jF/qd0V0tseIsWGHv3fNDKhvbRuANKUGASwSWqAIEtXzWRW5K
3KW9xRrXOgGEeHo65V3JJzqWKQiY9+urUTkrVQ2felX24Jz4pXwW6ujr5LErJMBI3FWsxxlQqUif
wb8IFGe5s8Jxmx23jq+B3A54ii17vF1Wgud43Czt/1VlTyct+RjOaMGFfXsNM8QV90SLniHKnflG
nvHxdFPrPtBNne7YmGhRaNZ41sLfR0kggP1Nrm6qpV7X0DDvR+I/NuiRvByqCVw2l3T3x33xE9kX
24n94s2r0EbLSNPhwno0+y0P64lqWehvZtbCDtbIYI+7vefk4TRQxc8LdC2AIDiaBe9cRUp9Posy
ztbEvswXqZkt3OsZBu8g8+D42fPAml5z6oRvAFJXmYkmyDQtJqP4Wxn0yz9yCtc4RkAdSSQvfhOB
SSYiNJHZ+NXt8fVYvknoKq3H0IWNcFSZIX2/kvkGDbfIgyM0lf1I0UZd43nollvJfcwv7ZtdoZ9/
pAYtocdENT06LLUwyFI+hhyub7Dyh1r8HUjqFBR98VXRAXzMbSz5cUj54+opmjz3hm1nHOtwSh59
IyXlS3PFjoepVqfbdzRVYO5rgBwBj35HnRZAf0xNXuYi3ZRdQpAQ9dLSA1vpoPX4VIuD6RP5W8mS
8CCZ1W+x+Wc/OboJtft7wLlOHxeb/P3pwBq3b7ZFE2i90L53PApfNzLnYE71p7p7mSxjrl0Jnb5t
CvdjcmAPj3K10Znrq7AjPLo9MPDYCHggWjld0STYRH4OJDow+FKleWLrFD0zV/b8LssFNAD1vd4t
1SBnB7U//TTrrK0NciMmqA93r5HSNtop+NJazJ6BNScFNVBsnHe2IQYtAvupM/SjEv8KilQIF4Lb
jeJUdxPvhV+jONht0BbU1lkqROzHd4vihGKLp+DNrDUA+ekR3xZAvl9UW8UNx8W8LhF2eoprS+Gu
oUuyFIyofl189ktefAP5q4hphus8xkxr1AhPDJF9EcI50TMjHZuSorpy31T9U9JyEJZTOqIQl6Vq
cd9oqN8t9nEYc3+WzT6uISvHZo31X8jSuWM/sbSwht/c0Y7wfz1G+15TiV7NMDqUgvJQmeduvIAu
82x7eFUswLONcLQflaWHSoM5XAcnNhLNNIzyWOQau/gvixwy32GtG+GpNa0PAHXMbqdUnszrmNDn
FVHrvTOtza2ZW+5JnUJ7GThMvJJZVxZ8mlCQTvLPRTU25LMTCs5rzmoLUZHsTPbO7qhOdJ7qPoO4
PdzhfXm6NTzisxKePhRfTwLY2toeD49epRpw23tAalPSawqxIidMQ2PRoBWs6nXXTv3+qdQ5K7eg
gm76uV5K83vA1vdoEHGOe1JuCfyIy+bSyxdcjRLVRjwnU+UDZTrEdyHd7mTJYZkKJnXRTDUnCTch
t6I4OkGcGPdgnz+IDy6iwRi/SBe6ODOnQILKmlyqWHn6RWGfojncMX6k51+F0sQsVUJVgPINoZvs
QaKN6UZ9LaJjVKrZE9m5pznU6LFz+boxtt/56tcvLPBn25U3n19oWDuZ/l8HAlF/cf1BGR99GU6M
HfWBaDoJ36A9fjkFVESF9VDBSu8D+kOkHmXeRm3drIl8prfCplCOJ39EU973hbcFQ/5tFPXpR6K1
Tp4NSZsjtnBnUT/ap4U+YiYeMg8wT1lL1g8S5LUW9QksjrVliZUrmdUZ8fQRAqDhwKdtb8+YxoAN
3d5gN7WEFc8i1UNmg++xXmbxyhFIRUTVRgpdU72gMucs7mbp0SKHYv5wDrfm1WrqjfDbe1N0wpyp
Vlram4TapGpbanS5omPXk/wsQgI8O752Fj2NIdWNVGN0U1OfE7jjIWhDM2Uv+6ItSTLE7wZSXtfP
79cJ2eoceQvkZOErMzHo3teQg0FRKYb9r8jrVI6ls6JqmwipOtW5KgRl8OvyhMltQXBSLV0YrraM
tl/XOQOBXoSiSd9dlcGrjhCPJyfYucEho7xbCrDyQDxPHQMWxf+550HLh3dz/zPLHf7aT5/DmHGe
S48O6vfRd2hS1ZpN47FVA5T0kH36x3fPn65RVCx3IXvbYZ9bwxesrrSXLTSmnwT9tydNksNlgVnD
PQPpt8X9WHzw/K6eh4fHw8+gctSsQEZ23NrsDggAlh5lHbHRBp4fZPUfYZXmCgjw5A7mxc5vujV8
gJZQi641eIkmhsJF31ShGGBSm4LbX4LRDZU8c89YMynJX86LKJMOYlRe2FcEwe2ACQ1TT285qFf2
I8NZvPzR4oSfECVDje1G+E9CJfKp83HiNCGd4r/K5Pk+8dawIyIOJO1hRFDYRyFDcqUvC6KhpUJn
dqpo1FVlumdeL2HIu59ps1+MRZToAV7UVK71dVFJC+c1JmEydTVGm2h70nVmu8epGTkxNuSh8HdK
KjcW1QRGMfAiRGHa1DgFpnIp0XO6oXR+cgcuTlCFBLG3NCSnCCdCshPlvbuKI8eMTPPx5L+F0DlB
2T2TgvBKDYkIB+HqUjWU4wnXQTSVkK4a5KJxLVHpN6uUVeQcWjDcPRso3OLVDwM8ljdBL6ZdsnRG
KQs+6jbX/M72QGONZIFoYT4jmpsQmu+ikUY9bEY10ffXfdCFzx10aIY/X3mb6oc+4sDbsW1uR/B7
pMguzW0/MWr2KOsgDLf/ZNms5EseRIZpgyc6Wl1jB1Ytpbdh4DT8+VZBnhALMSfRYt7DjtEFjW+n
YjgOtW3BlbGsaAhPsOAy5YQR1Uwh3Z3N2xjB/5SNHqD4i+fViHRHHDRwCwFYup+IkgA/3NtZeum3
NgRBP366XnGRCE6v/8kvu5k6pE+sM9FLyrgNje7X4nlO83FvbT8b1g9ccl2GQKum2LPqiy9tCMGR
z+r0z7oORZHoNEELkINGhl5aGSm3m2+YSMY9qZuQ0/lQycWk3IdIaOJXt8Mu++zKPEohStClYvj4
Yr9+8/W0jZrUSOpQ4ydcnOQ4tcapYEZEezHcCu8nfsdELuR11QlUrUKHJMt2WLsSQIuPQDlGLMIv
OY073BN5wCfW6foX3m3iM3f+eN6Ad9wxCJn7YTnYtdXzq8VD5eoIxlGvtTyfaRU5C1H3ZB4ZlIMc
tLLG9v09n5Mo3M5MpS2XvE0/+IQiUuTceOoMVcN4rZ2RKU+xEISotVa3ga+cFY5HOxurdLLtOBCf
iDxteH9jYP0gDkTTEsylYR9+ujIgxcWRft7NNfJUiVs8RW3/m5bzMpSNeCMOb0C/uZ07Gv4oQuoJ
75gTo0lVR95V62Me99q1GjAGi9Lc0cPVClQ2vgGbTeznPUCEC8sochd5VPCFLOnmuQE7fDWV/lgE
EhROUCTlwAHed+H8vgB9c4S3ZiQSC15DCO/h7aswXhbvver8L7Ne/GimTPjWs7d4raHN1R/Xta5A
zn09jOMtnhPBsrvUlgY23vuy9O4okLRJRmbIQ6l+g8TB4T6RnmzAhiV4PlO2UJ5uMbmgxmYXYMmN
tgIUdK82kkuND9FI8saonSkuYcL1yxBLiLl1Hzf+SFKnN4EEKbmgAIVNA6HuCfxQA+iDAooC+I4w
vZ3gwxMCVUpCDA1RX963lbXWdzzJTQpy5hKQlLGRWlObf2Dt1G8H2coCkTwTkOyGqA3jcdgPf7nA
f4pScdkB/K/m2ajswoAiX+stVrcQ2A9NAImYvuTU1b7NH+euLEKFuiLo9X+wPPgU24+Cfri5wuE6
lsgTsTSczm/pILW0CuxU099bvDjZ/oaig3dQylNOYaU0xCjhnLv/gBRs3WAyES5Ko/c5WJwmgbk6
fHi71dHwx0aBWwsWp9JH3pQWz8y7SbhQ2ed5ELQBGQNfAyGErWPHpseL6oWQE6x2QRD3wjkrPDFT
WhsyhwYcGuNd0R3ZC8YXDIo1jksM+chc/+5ny0xas75X5eYTfUE3u9zL2NDS9OhPWBGf8KcddfRc
UooF5kl4vYz+gD07TQm+nhKYHHmPwq1RcMV7sTNXR3GzcTOTGzJwHioPZQU52ctpj/WeNngdUn5F
ba0dfi/9GlM8e2H7awBUhQVTk2h5BJi+yayQw1YgU/uOzY1wPnGVHP+y9WsUR57yYAcsm5jmDOs3
FOnJ+yjlhF1GhFzl5OaSC0F95Dauk4ER7FZFdRRPEf5W4748o5UwQoFVt0EdurLNNXhpXyuhQAvB
mx8FHAc+jOWaPMYL80c1QWsLeRKgbISKsdHZf2OvI1PyVfcZPK5qH5nBbGlgB/zjhW/SnlOmMrX7
Buf7rmnKxNe8Y1oEu0IbPloitzHneccq80QL0y8WBs5unIktmkVLXEPEtTeW5PyhFHaZGn6Dmqy4
xbjacwUOSB0bqg8FMtywrZdkCvDZUCED2iJZciyqudt9mrdeI5MjZi16kKGT5U3zbtk8K75t2McY
T6DHZSEYji14UMZRVxu/AoXPFu5EhC8aBAwig1aYEx6qSZhuI+YwkPh9GMsBQUVtJvMlG4BdhndE
pcYUwxpGS3Nk7NEVNtpkE7KMbNV66xaBb8sB7aDLYnCbiXBzoAeu4yMuf6suA/0l+nlGDmKuYNyd
Ue+729NwJVw3rMNmvSqgBtN9QVuuyTSqmmb+m60ZQV8/BDYQlGAMw4Oq1fg0dGjAzYiz1EpfbhYr
AlPpeW66wKqgwhN/Z7QlMK/q4OyNPAMFVupiQZpAbBAYabZ2E1n4NfoDnduEoJB+HNWW1r7B64Bh
TDNHVXKXIPldev4EXZbtHNxlC35YU305A6fCj6AZH+tob8TbKQDetKpaXvv4CuazbBn26BRLC1Be
Dzb4rKTqpI8zxjO+ZARjZJ4x3fFZe4juQ010SSPe5DdL0ZaqLULBe4p+swehXb4x2MG13xQAGexE
DfkHiOzNrUNNzpyelHcRzJ30IDGKgU+r4WEarHDml0cBnIXfvMA9EYoZjKQ7BH6v3kfvLuAPQDME
3cGREBvrhJOS640k1dqRJ++LYXE2SIgjRHDXSQOGeSmBomLFkCmPqtCWYZlj4GzdMdI1ymA2y2Pp
rVmYHgBb1J9N7mI2LA/EETxfPKRHps4HMNvXnwpLyppYtu1jo/oJZkS+Rc03LJO/G1ZPt4MnqWJH
bJlfYMM6hQ5Nn/F/EEyKfw/tOCQ9iS2p3evjrOTb9yo1iRO1fOPOThnAk0unDP2nSCkk1dxI+sLH
q+JJ1IF5ttEUKzLJRBsfdOkr1S0tJPX83yHBWl5QP+cid2ezTQRVF+yCPYi3amhOmQGfJBtfXxLj
dPzq71WhYHDFCRMbKpoUS+Zr18zbUgfxiVNj3PJRGyXwb9ipE273jnjDdYkIvKg1xZtaTdveTrZG
7RMweqUH5JiAcmW5Ugvc2+Q8D4ftKB0c88eVJA0X8seV0Pt5wLKk+gUkcM7/txEFK3ufKkFn3vbA
sQUaXTsxvtj3LakRJgujONon17x29Mw96kJclvycasT7QN/D+PX+XSK9UhZ4jmwaY+OamoJiW3vv
84Msrx7ZA/XGdJsaT2bJF94oM+JjWa30GyKAbgWyaYgXoP25vD63ad6Zmq/JFrGwjijxLPwi+i22
HNMibx9UYDZbwJXHhoyJEGKPZDnl/VD+KCvms0s1cA0NNxyYEWOYJi3ALQdR4VGWnPdZk4nO0KN0
FiTNI1x20EujbOY6WGPXRg4E019i3B2yVLN3cl2sGcwoR72EJtuhaI6Hs0iIol+0pLUPqBf7Juwh
ZoO9kjKk71Ug3Ka/jDjHJOWXntOZVBGEp6IFs1fzpHffMj2IBzlsMtjjdXtRbp5cSuuuUk2VVHc6
9O8EvDHAIsJ+KOOGxjP9xY+8iRukeJGVsm51qGW7oGXExOayWlIHVyP2D7pQF1XXfVcfLFbr/7wt
w9Bz4p7VV6htBhRhMyUigdXIASNtA3kYoCWepKNyldikKAWZS/vGUZEzECWFNozIYy56x+Ds9O/b
b6LQrTN/+pUgQ1WVid9IkptLurdm13IfOAEoIHSmdHOljMwIzYwzmjv6xV76hnuyC0M+BssvrHK6
kHR9LW6CsLUaVK6ptZccHm6T5agRktfvku/7Jvx6EoM6sRLMMEUCB8I1NIH6T04J3fSY+ZSWIPc8
FzPHAW7LG4mgWmizoB06tlfogf8pSbAavmEel522BVd2FtLaSOBZ3SNh5HDcjpFDY6f/31Y4/ebH
FD6wcpN483oHsiUZGtSzE7eG90jIJyA3t8ta53iH1lYwCqFH1xjzayRz0HxcM20vDeP2Y/goUqqQ
XRwOATLbPsT/fdOoe32m95G6x0/dgEbe8M52GMVVHANeLPGnnJepXPXW0aXqQ7jTgJ8qfx72liJL
uHLnkXuhJ288L2+uVkcrUr2woO73kUCJcArNdSM+vRdo8B8u1wqqQ1d7w1bXyahiFMRuFc06r+Sk
HaWO5DxENU/acBJeVMCc5lrbeNLuUCi6dQbVdAZMLxlw8stFnJ3GRB1p9Zw36pUYj/YQW+WSmxJc
Bkfly6CaUtfJMpba4kLqLg0p+JnwbwtaGw9W5z1jySb+TnJ25ClUdUU8f/sODEQ1/1lvefEbGsZY
EdJGroGY3iO/PyADXy4wzNHT3QOiOCtJ0GXvwTAMU2IFbRq7wRe4BMmjpALZUAUMUF4lZQ/CVgVB
3q0hUUZj0kdkorUZBgLW/qTaR9AAcuYt+MQVgaHaX9U9tsSEWUKYLuyKueX0xHuVuZPszc8NhN5E
2+hBeoTd4MD8DfmwMHUZaL0Nh8XgjmI4HuCBdtd6AKyAEXwuqG8DAutNIGIHrpjEctDMThD4cPLP
HQruXF1qInhuJ8EaJ7VO3aMLm5UNCXWDkMQxmSfFPhVwafCx190GyO1aqm2tprvmBOUu8GfDqtv2
HqDmnNvCGPUoa6CtlTMrJ4ymI45WHANI/u4DJjBWW8PifBE68z5hABmh3gUwAN8COjdLv7P2JxMX
WeR6TpbpapMT4JjDePOgCkO8KsmmFbZdFLzqaj4M8G3wCU5aZ62oCFGda/7YLPqLpXZaeQcRXhfW
Vqf+hbX/If6HSve/5+0Vgq1FkwIGXJDA8tGl2mUB/MSed4fU2g/+VyWYXDUobPUAS1y4jvpW+Dm1
oRNgA3HbFAsmNNX9sTijbz6m/HGbl3H6SUHHctxf/RwesY9CxoBceAMFH/FYGRJdnEzXs6xWEFuk
8gaC59eAI3bIF8pLkSUxUmHWTitPzjxUw2MC1N32qNvoff7AnGDgGwamuWC3mEGB8DLshZYExOPN
jGPWR0T2IUQM8epJw2nKYyrb9/UHaOsEVJ98YZNGoI/kcE7P7UUVYmCiFi21VGFCgIfFN/HM611m
DSrbTKlcGCrbNpLZ49/mBNQlIab3KjdZWgBNfjtMfo7d3q96DVLTvEIsRGId905hZ4mq6AGOnJBs
XXjKWTp8PokdNT56Uu6WxYBywnzTtuOOzBYx0rXDEdeTTUf2hzAHHHYmr7xRHXEsKu8Gmkysrfic
7WSzhCFtYGqdA4sRde4ZytwSi69S16q1H1vRkqEuS1rdfHZzA46BEwzrCy79Vu86h2fNzRdfgZa8
ACgRXFsOOhg7rW8wthz+Ff9jwDuQKJu4kXARfb65O8c6Z21MtKPnCOkO4MzPpOstUxdJoU1iyVB0
xcHYoYBZiTRw5XIYwhMb2ESvA2Uu0qKvvgfC8hpamMWn7BtpJnPJbQvqz6htxqygQkDxPQxD3c2A
mmTooucQdfGaz4yGzBe35qv0b8j6NmQ0UHFANPNJp3DIZmLO3TjJOhVPw/EuDsKbxQtgDQNCYpJ2
D2JIMGVP9lK/fTgyxavfbM1srp0L5aylG5i6n1nadw2qtvOSTj8EnDi7K5S6l56G0mYV4erHfy5o
IKNZg8wNibWiAQnLJra6ETpONafaiSLW1V0iS2pOIlP+iv7yq/RmNj7SvZVeTtHVPXPpKL89dnOk
CeFkFo+Gj/DGmUNh/qHOwW1+q1jx0zjF1NTxqNiHh9pf75XWHl/dBLHwAlafjO2VgDM/kOF/ZPRP
y+GWUtzTbRJOZmiWMEkQ6ZtEtw+A6bxWtv12F8Hc8GO0rRqMN9gmBmIh0QCeCohFrptTRglA0Xc8
Z1DZsmW79GG7sfDSO2ed/8FCod9jxDXJaNRLa/g/JuuE5riopfxRNVSU3rDbz/ZffJkV00uJH1hM
Tz4TecCqBd+db00qdF+pFyDf661axykUTMNk2fptAwo/Qal52tNIrfiB1zfI+zT4ktnz4ETrf1i9
m52S0BUIrXqTC+eCF95pJrAKmvyukbssqi5ATk94u4AVEV93QHRy5JWIrGw3XCl8ZXIoW6649oVz
9YXCb4/NzuubbvObsVDotb46Ekm2fdRmz5muX8gvTHlYXJU7lLVGm7ocBtpdEcmkGX5H/YfujHNm
7qwtUbrxF83xqtRsoqc0pFT9LjzwCeLAEkyNJjXMUlck2KpIK0+62RF3AeGq2kSn4r5eJb60nU91
JFyarfBFFtQOh6aRP7bUcD4b3fpjd4fWtAQJB2Q6TcL231VunmSupRJ4KywT7xyyMweM2EmlKpA/
RUJg1rpzjhuc4V5B6chLIje+rppa1g6UYHaHztt4zl0ht6D3DO7ynly6eo8xnKd0TCzn4TrQGlQN
TMfb6mBZ4lyoJTjdO2uzn3ojc4t57BzURUJ9aYtn35bXrlAuyRqdAhlpYJdvFheaAl+IR6aV7v1I
9B+/pJQUUIdN+gS/XeCpQuXAHoaMmBYn4ItSy+YqPHhyaGSdeJxSIdxywy0ZVLPkGDPUW/DjjXvj
tmp4dLn7k9M8tWGTTQ6alCSnHoS/2q5eWFGxAuh5qINOC11vKXK8C8dzb7nMJQzAqP1SBpDVlpNT
xgGib8DBHdWr+iPd0PfvrwOD6ix7IR6wWvMS+UYECq19s8gNROmwwQQt69wMO6eYiKJ1Gdu6ToVw
FbuL2XOOzfbH1hbotf8kxc3LYNkmZBNvNWAIF/UtY1iX1waxaoos7H4DfTFyeC5qfCVwGigCdFJA
g5KdAkUb32VZPWsB0YB+WAr+S5GD4MO8KunuR2Gc3l/T5/GFqVfdznxt9PkjTVHq8wnXBUKecHT+
aeNvpAlzTavxQ1NPlz+Y2MJOUVO1bdVU57dm2ggbwzGGNku9V+dL4bmAeiK5fGmv7WfRiCSbvAXA
rG8jqsaG+Z2mimshdDhqegfx65br+2n0eQx+jcy6mRgEgnXdNZfki8O1HeOov+f6eJ3baPIUgnD2
2l9Zei+RzR6fM7/eMxrSc/HhJyOaEAN275F871VCqjHDtUMlbq/oF76uje83T4hoBJ38/1SFiTAr
ntqdBvy8+aqfs/Zleg/XqfdZ03YLCzY0eHPYnUWzAQpfFRaUqQwKF10JuHJ7dKHJfhuhYGCmsbtF
Or+0MlefLIlKfXMKXWnj4fQegPQZUwo7tju98unwHQ7aYBsS6USo9fVgPj13iPIH3nEazsgnzeuK
bG3Ix+mdOrsm8/eX/7+gEEsUn7GAZSQXq/+fOa0kqf2VbFlGXdqnUkOo9lVpguEFms02As04gzC6
Y4LYfcnc7zXXo0fbwajQwcMG9DMCN7/e6sf9CvvKNWwHPzzh6mGuPbNOX1Zwc2VfhwcQSnVsPeqf
ViBukdSFi0ROgOZZowjxUn7+9J1VlyMuKkC1mDUq1UpFktiipwUfjSnKf8lC7j/QAbD/gcT+sW6Z
DQJwrCwd7wAyVhwbdclXdA1wVX9D+/HQ5qlyFQjZtAcEg31RFe48HQhH819IFHqqJY/GXxAjl+vi
NETUKUnzjgraXB+HtxS6B04x2kmnAUtyRcYwOJGI/i3Pym25LnAPG3bd3gyCDiCfQ3ewxB0Ix7CN
jcquY48gHVCSD7fuDRO1O0iVz9LwaL8PSmNkVQ0dCjkVpuZLQ6OJwvkGv2QUEx3raSpP6Rj/4h5w
7NdCK/TxwSETiblVlUJET2OFOSFcLbjNNjufev+g9Y0h2f8abzLiJdBtc+LOYRIQVIOqo7bx/64S
igpzMTrqDF00/fxag6xerQR1jorPzlzb29wIrt4JtKO+m34XJIhaSW7cqXxT7yqBYkd7Zi2O+QVG
/yETOHjdGOFZ8uvO92QicE+rjex4X+HAW+9iLBA2Hcq3kOl35VJl1dTmAsqNEzsk3mgUZ8wtfxoY
5XXi0H8ShgnTF+dYideThkEPJR45n+Ap1T+YVVrHSxPQVYeC7hE6VRHiw96KB2hv097m95RuZCzH
U0ymp0O0oHO+0BXw2TvT0YIjY224iRi2hql+aeu9WfzZzhX5xt6L8geNDIX1sCfsUuoVJmZZM24E
nMJdbLO2+gT3LpC9Ux/bVW/20wjIfxnr3HFVHzO4b4Totxvx/5DpxjXPWd+cRFx30/VpwnJMN8l9
nxk/eoo0RmTKBrIsXzxj8BvW9E0bdsyowWkl+Us5Sr8+g73sVSCYDymbZA4yEEhH3soLy+hH6+hq
LqwLfU5fvP1jg335I3IxIBM6/ScAyTPzB/DRmuDzc07A4oHfHDzcAFEEOU0ZltQ22bY9OROF/Hxm
PHFROJlhgT2S5u3V8LvWrnRcw4Q02WFPtE4ezl2IRb9ahhgHw2XOXVW83ASXzZZHPP0xstw3iKGB
gtqomHSoNFZsA8YbbaoXuZfHcbQ806SSh5M9ATjOk3ay9ZxDj6J5gPouqCjBdvozQqhKp0qeXdEX
p3nif3SP7deHLp50akCJ8cHb0gIcHEc/q2sWkZqDJqIlZyJrb2N7t3GkwSEaWjg25lnmG/w6mAHG
SOPPjIYgz/rUS1Q8lVExWDhrOacJD4XqQiC5rCvxtDJ6bisqKaNlkOGChqSNKbsx+8mC7K707Rnp
MRhUPJTAXY63B0wROHHjSDwPO4zQLP6uhFb9YQEBAKfSPor1WfOJkLK/+WFLQQrWF0i+ckqGrL6i
VzzOHgj0ycI3/PgSWp30CMUWz4bYsNNEIcZK86+asNQjh4h+eEuPX5pHZym3l5pU5/elawZ7ZB8n
nMBbUTHOpcL8LlGoc7HnfhLooNbvx87GUV4MYcXvIDr/NoC/ksjszvrw/h5vHKwSeiU82OcAGV6S
gzDm2NH4ouTLMwjWmTEZDPf2IPRuLNRRrENrgnR2FEoTg10ZV6YWiHd8cW/DIZK6jZhREuY05E2b
ZYhTZ4tq02yPxRd4RNGVCDCBoms/rY88I0ui3I+MGB5hiYYjNIdQKe+ILue+3ecOiBonpBD8Wkw6
DyHZvgaA2Hd8DLIV97wdYE338AQbbC5plR7O38kjOTlOYl2GiU+dLV8GdMW5Th1tD2DqU/wjbUtB
7KlZMh1Rf/wDfH4JP4BD3tN78IOLGaX7J9rkwBRg7Oj+zFgyG7ylRQMpbK3b3eMa/2scCFbl1/za
RkqLWpU0kF6ET9rRcjwEOz0eD4scppwr5zY+4p2+vN46iKICT0WrN94hcWMtLU+Q/8i54ML38pxN
mkhWD92fCEt2Ap6AobwyQokIZ2VCCF5r1bg9PNLefyf3hQf3Ho+SABDoz3fXAZvhQ7xqzCF5WMUM
fK3qGSWlY+9xgnVjHA3n/dORuVLNd3YIkbj9DaeNy2kFV/SdxSuL3MhnY/HAGrG9sepmpRa5Fmib
UHPuLNBtQ4OHTtG5Zncupzb9EE2+t3/cKs+Mrq1yIkS4bLBhX+k6b0Su0QaUFPqYLfKy6li2rOgZ
QpEj6zrzdnFX9CGlLxVspczdK1yQxPU3rN//luGimdWdSR3MymNLfx9AWPYkxtYT/0ZTqYRr3zbW
6gQ+0tkRgCr9hbH6lysQXZG+krOsPkrl/e8KyIaQyCI0MVPDCrPlJQi5nJsATKdLZ0KZoohvSdxz
WwR4YACtdhkuSk16uoItwdRc42Y8ZZUYpd2CqSjMp/9bESjj9gEwEV7XfPCBRifeq0yBdpcZZgjG
HE1LbV0wE+1lkS0nHrPhg6jz276Uw4gNS6x8jIyHET6mJauOAqKD9lMsgnJxm+O/LKDPUTQakYR1
6Z3gh2mU8/SUjzqxUGMNIQWfUTFPD9NTaFdD07Q0vCXlQ7/Hd0bIhfvsnCJm4jlqSr4VOgTFwLKR
bqwmsUARGPBBBP6sjslsF6MRYHVm0+g9VlGMLVJrCZrtTZvkBONtRRJfOjXol/8S79LO1xcZK+h+
ApW37G8SLjT10k/3227K3gf6P01uimNudqlfkRfzZrtLrI/5ItbKhmwE7VbMwBg3HUQMFEM0p6Wy
LjxN/ZqmDGAgV+Qn7pnRQO02wHPM9hBN+eHe7nSBbEijMQL0wr9lbQ0MxlUhpnzEB7qW/pUJ11Ay
kaxfiw0ZXwL44dz6JFt7SAGg7GajsBDZA+GQCPPTXSuYetGhWGVdvf9dHMWtcWWghzRfkVLovtU1
Hpacv41csZxwFWdJFRcmkK2+N6clkVx574hxGs9+R0WVoE9+Gqy/SKemWfsFbZshXaZka1/RlgFV
xXtvjob/kDZBEGIArguCDwAvmUTdUgbsWL8OSiO0Vsq8+hi1aWwfg89WKfk7WUccp5hE5ZqhVB51
ihg8CyT3Rc4rCWmRPx71YJKJLwj4TteVotnJoqC4aDCa7E2dN596cXM7shinVj1bTB4o6hKk+uxK
+6j58UM1FhpcqxYS86iCBTWujLTyNKAbLC9ofEL9hvvbk5L/eob+jNgkK9xbDDPDip/7lY+h4EH9
T+nVRPYQrnU2YxZ8WA48DMCSCu2U09f7W4urxdJJLPQqPT3eCJgEFc1BwF8Yxhg3ZkAAlMedfVI+
/TEB/lxNQV0tlunJnrvcEmYX/IIj9Rx01gcu4Oj7J6SKw99E/LSExw5hTDyHzXOxGN1SJHFBvg1K
TpQ5P3TE349IREEB4CUp7HffKBDy9ouqd6m/2r6IJDhosGxPmI3ZHyBG+vuuPvmtC8z0ZYsgTgGz
ppklfXZU4fPwLVth0zemGFL+EGbsAVlU6kkpzXVPJoFevnrnisleOcXXvtQkb84TKhxDVXM/8zmE
7012mxfoJ8IYTDXLQZZ1VLPgk/jNANYXNxP7OJjcfHw168J21gmkJc69KbyNPmIO6dBPrgG57Kp8
CTco/3jWjMq2FPLXNwDf80u8LhoxWKi+FFL+fjEelXHGkYHtCI9NEpUTcHGPBA+VNsDDoz1kmlIX
uru8qNg8SJZJ+owtCefTLGE50Gz8FnKNkMQ5DCZs7BEsgK4X0aqugxwaKW/ysPri4WKeqZPGdpU8
4i0KQ5i66hGqx1K1EGBOT26N2E2BcoYSfGIrMqrfd7Wo2oVGGB3JUwmhOOC0KgEVZjUuaQQa4CAQ
e5aRrk5cAzorpCMc2TDTXT9POSV+e2815VeqWbuiZJAbeawomlcC2YFngFf9+PhvQph2euk8Rchx
X+Qn1Py6RDHP3r6dv0jOYdWtmj63oX7EAZ6qy4hjjMTF2lQ2jTJMK4fdqDC96VbWuZpg0B1JeXhl
D5ijk/7taKnmOUFY2YTqUNtoey/2WkDaUELoprOuqKdyvWqOq57FTei4+nEIuo/kCJzgP+KeJVAe
UT9GSbVibNxTDM6MCpPkdUq/C63gZ4P5mee7JwLVh2qjYphK7fbMIoVmVl6WzX8V9zpCHCRcHmqU
glutuNUCBf4Mb2xbRpbQrk7L3vamxC2ALCooW0z8+eyDgqoh7bnyAyV+n0P9Txcl1Xz5m6CKR+vu
Al6cPhJtmcyp5v5bpxV9xFlDQU3g0Am3+A7zq+cctWWPjJrE4GHMtgdun3bgT5f2BcT28X3OFFWN
D0TLvKgVk/HwvoYq3etJ+xQby0OQ8h8mJQn3bvlsUG6srX/Pwj3U92Bz6TW2+mbLPz3jy12e74iG
Y2O7vFOzYfKRGvijLb7QdBtQi5ZVIzMRJRSKqY6fg1vnVBPZ0hKRvvXkrK6foIitsFToXfO6y76v
/VSQmcxvNQlc8aob+l75F++A8fSXcHiVR5onF+GYut0PYFLYvNzRgtXM4FO9mP2blw2wsNF+VYg3
sWmZ3ZuAyxPmbaHMiafVUSJNYfDGduSCWBIOlRpvvIvSDyH7EdYeW9YLcL780I0S421E9jOJPlze
/OqnGQntPm1mT3oK7pdR1yHl/JQuTFqRCGGVQ74LUxFcGPfRNAw6kI7iXRyS0j4mBYfm36KjGo2S
CcaV4KyqO5/GqMiTTifrVnQC55PVoPp6AqZQEhlDGENT28XNFo2RjDfdW9oy2p4JAWk2vl4AVU4g
nPuMGY0uYBBC7jBTowqLh6sIUynGvJCvvSucPIbU1Nbj6akWB7pObM30Hp7f1k6SB+zCSfCDUEn0
/q1WmVk8VgD8QzWrw6BAefYZAh7K9o6EXLpVjN6XusLTVUcEN6ANvirAogd1rmm3iq/9UbjIQmTi
vIE9TrHMwb2dSDl908Ku0+wX6Al+54d2/s4s2HQokuI42Yy2cs1QDgmCOQmzIbVoFbKGS03ys7Zu
g2fYTAUnbIUp3rjomRNaYyma1ZKpkr747takFs0rvYImqPw+fI8YtPugya3xYPfW5Et/im1KMHZO
2uch9vTwRYoYP/zpRAVF5mvO42w8Vnv9CwYfQdFJ/2hA1R38nB0mnhPMzztP69H/YHed5IakRVyA
dypwSR8jznyrR+swQQxdWTN2/95pdmo2y6/b5uIESEGyIKYAMaq8H46A2ogrPgssiQ4WS/KPmUv6
A4CFWvPtXmQTQkR6cjI5Al4FBjy2UvzePo0pIQoSM1hLKKqumFEP9Fo6N6qGMJZwbsIOwpqEQ2C6
EjlbbCRMvEpkhFd2zSAJM9HFhY+vfBnHflSq1jWfiVg8sLRRHL6S1dcNSL4HYTE9Wf8Hp8VWEiZA
8bKbRp3yueIWNKCwmWpJ45V2l11DT9KXjKrVagV4hofsFQrLZJISE/qtBn8gMv8/Fmt3izOazeHb
Hk1kYuMrnv5PxN69FoNE8ypuILSSqN3P6qmab4HYFDH7Abip55gQCKfXAI++UkWnbC/hdMqzRPlU
zNqtT+rc91xPtEHHPOtYePvNtpqwtt71iVbyS+41Umkl08D6Wvg2mEkPFdJtGbXflsnjn065IOo0
BO2ghGkXoc4P244rnEjxpYkQaXcYatwnGtCClyAWMlrRtsTBGK8MrjQN9IfD2GarK1wlhmUd8GvW
mmSrVTt7f0Cg4C5NMTWfXFK1CBFw+g03o9dcVIDYLGQXcoHXGoIe6zAWX/fNeKOoCIlNb0/pwjKM
m3hwAuV1U0n6016njOGHPNbFqHMZMgop/iQJCK77CBSHrAZIVbfDgB54QXzYUGpM7mFrm84CRlc0
t6aC87GUQypLDXwu7NJv3+Z4no5XPiMUBKfrJ4/CwofVZK8WbGdhOAjW4ETLJjj8FhAnyeXxnZlk
wZJTPc/DAZEunbJ2HCMU8XEUuINlJb3YKQm432FaAJmG5ogNXQrKJj96ZoyY36o3lHxQkgl30tQV
kXEKKMqxKlKRMOEojV2B/CHaAE7WoHXhy08yX/noerD5cf/43XskxYrErhEYM/5M7MuYvrHAypfr
eVDfZMr78CBeX8BwKcm22kP0jSvTKmq+3lpZjRG5016LSr73acRpFGI7Eqn/cQS5nAoHEllPByZA
AUgpVAgv7B7rzKPofRjk8/pLU7k0ulPDxRIOMpLkeoNaQxB+kTGchu7s1uqp6U844DS7wCjCcrZV
NF90+vX62zo9Rk8pVnAt3f8WWD9IvBSE5X1Zau2dY85H10yYN1Vz2Fci1CJz7rjXFEhYpYzKxUJJ
qtAP2PauPZhATxs760u4fw1onBS4gR2WRWjV2S7yxfov27nP7XeuZyYD3sMcDvduNZGuwjECTQV7
PD4038B4NvDfhqYwRZwFuk2CfLMQ2lfp2RR8vLWBaFwoi5iW+Qhr+yLO2Rg+6KaN7MVgrh202g2p
7aHi788Ck1t7VPQev6yXU4Ou7gOzmp9VcBtOPp0pbKrkbHAV/HEazgWUu9PloOXSU0TmCeg4g2Fp
NBFN+6sQMzzkW8TegJpWxTU4FuA2p2aZRdyMEaZztuH7vBYYaqnU3cWW3y5G/h4cc9Fpax9lsXv8
rCOxcefZB3N0ImzDkLVwdGcllQEj0xWbsR2BjzSG42SRhho3+kDqYWPKdqKaGXfwQu0FNW8kbrOb
eyN2u3igM/HEkVNgw/4dyxlVI2Xc//yJ7lgqEDBWDyK6fiDNhgKR8q9IQi0AfdYZ4Rx5vLpcXQ2B
UWfIz4uBr+hfln3aF0jD2dEzAQP6WXvsxxSnuWQPj7xJiRfM1VbV0gTEoWaA5OZebJOfqm/Xt5LW
A3aBi8Q7gT991xjDTcoAmQ2B0iPrJJGqUY78mzSJ63K74MrF9MBgqoogb54iJkd3PrlwjCraZxVI
wapeEL7PXXcDFuxy0Vt3gr4C6/AJL0eThM5csdAWTiY9HAoATsSa8uL51Th84Ce3Q/fJ+/IwUZde
L1cAgwYg7PMAAUg/JjxQnyQXnXiMsEQMIMFn9YJx9GCym4dV5HdBooS2b6HJOdkEmMMw0zGF0FzB
Dl23RzYAWLvlN4qSfy7U3L29DXCW9eTwVA0snez1rgFHYlNVNVNuUtFBtr4WPvbTwo0x+An+k/vV
070IWX6V3sA49w4ZgN98OHIRdCIRSR1kTcnWl4x9nYNp0+40Bu0CKi8UHAfgm7eUbu4Q0k5UQYpC
g073aMjYEcIc0HBk9x2YrZkocQTuNQAMZahiqph+q9KgBWH6+GInvnbcWfhXXp9jxj9CpFpcGSoE
U7stcNh3YlmDJ+opw1Rj99K0Oo9Rg5Svc17CIJTU6AdahV3DL2I6Qsy3oDwEoPwslVT4pxMP7APs
2CWPht4Jvw82+REnIckgW1V+iKh1kNMO1WA6cZW5j0cdP/X6+MDtMCz+AoAseuzdxnO4UiOlSSsb
mhDnWEZSHWlKoj+VasreCZLCS0MGRpetHA3QeCPM+5WdwDANsg172nLG/59l8ksMRD++cka7/x4t
rQcokGqDXKlmUZqXeoH5UQLRs/eQ6ynf85uJcCkAK13z/VNVkvbIGCyztiOL4Y/hcpwNA/DePPa5
xdmcPAV90JOJt2kgt8ZMT+Lo+QyjH96cJa/xXZhWXQKtzP0/0O9SHcLZ4Azcv9WsG3ZAS+9EUze+
CDLkTVDxTFJbpNqHwLAElY/lgfjNSat8w4jH9KR/l2u54BcruIxwD9Qh+QUSV9jTDMmzhY41/uiB
FtsHdzDghAsy34gC8f79V4qe5hR6aFKobk8YelMYe/JxJjYyVOJ/MP9kN9AhHHzYnMMJSbVtgKhS
lzJWbgQbPumrLQK3Qgp5pOv4K3sCcjdgZSqPKjvFPV/cx3pfxjo6W+BP9y4CtFr0+BE/sl76dvHe
f0B4NFNiy06I4RbBE4U907P+WCC0tFf0NQ+L2xw1m8NUHXc+ifKwEw4QqVBAYcFflCA+9ElyZ5Z+
6+qppSbRYOfO9STelgTFyTqtj3wqpmGlhB0PKlVKnaH/T/SuHl370cDGCKs3cvEzTdsxf1BBfiMz
7RBaecqaRebrMi6gOmu6abQtC/XLV8RltFDDIGtaYQBP7L5aj0p2DDmYlRd9MewRCbqKa00bFED3
2SpbZzYTfcdbaMHUGWEbjlAiCeBLEw7VtA1Nrmy7lLu333rbm+zUByDezUZz6CIIjKnq6sUmBf3V
gIrdjSlIOrZGfM00QUpWDPRuTwTYb+8lPAyJ/9wBnsJLORJ0zxUiu5AuzzNq4OZf7lCIX4xToWQ9
amK3BPnLZ3Q0WZCm0eKRpbMg/XeW2q1F8yJGYz+TtVWde0WeF72MPtoK0NQcAxphcQdpL5RHvSnR
QitJMpFNIVbISauojQXh79ORztByhO6QHHCV2rtrHREa2t26W+ZBsM38o1QnazSCtAN6rJEklDwU
o7G9iMctqQ/q59cFEhv7bYQ/Gzqcj+XWCvSGsHJ6s/PCz6m0IR7vo9cHN1BBeFP9k43/TcBNAJJJ
yraRYdou/JswRazkifUfvrgai3UK52SfDju422yewZe08EeQhJqAG9x8scoLjKqwCMnGFl5j5MLs
GaXyCitAnpkt+44+3vXqm2UjK49JBz5Jkncsh8hB0WebN0iyE2zkC7dnPmSdWYyyYrJyWvdAVR+Z
JALMyHtNR6809QU7w5xrAUiKo65KSIiMVa6VJ+50edHEty9tEMgfPEBGOpYMw6GJxVGoxVYjakfZ
krsu717ZxZp1l6/IuAGEFFPosExb67aEPeCSnmqF+4/kQz8QkOMZl/SoUbfBTYnwQQm2RYL/0QOX
YgXeCY+42+JxiCNJ6FjzORcLF4dqhTlMmikd6mUcFEWScOIMA138szmDvIaip2oBmZIQhMXFIV4g
R0w9TW1vblQ/ql8IDbpg8t2iXV6QCgko/2onoMWjxhqcrDTW17GUBOZQ7uw5p0CfI7euK3MBMGoE
asyByA86FK1US/w+Qo46JF2QOwUzH5fd07Dqpp4PYIZObUsIY1V7pjcV8IXyhcuygfoHglP9+0Rt
XsPuCNRcs37ogvlIaGOV8+2AnFYtIcyZupGEoSnCPQuIguQcnWsiJ9L8rQN/Gg9xaFtXp8fcZnT3
8oGnOlO2P7/H0uynOhMNiQPGwtWqCrbHgsMeHxTF6f2eTO5snoPOeOSo8upUHUxXQG9p3Y1ybYUL
NNg1rZjexjYpyMzCGY724Yq8+CJi25VFHVjFom30G1pme0pGqzyYzh3JBSHydOMkI4FmJEN7/nQd
Lj/7C0uzzOtD+YFI5Vy2ayS8k9oS1Faa5Qqsa8h1WXjZTSo5+4WzLEe9poPzmCmJgsxWt09gE4S7
9z9FycYf1t2wRpXN2hjggimWFIK/omclANtlX9uVerbm5lcPxJHsdfkGDzmqU9IhbC39NkkgPlOf
CormKvBB4N0k/p6ghXE7DBNOuCarZINTNnLAJ/L4wIuG4vRixlyy+UNkJaF4eXuWcWx3fbKcVLyr
7KPHBqyFC9eAafFmR34JOYMiqdmCjxuJrzTr18W3OqcXPQ0Ww0OML0oxQegDCmay+fiQuA2/ZwCB
0GvBgRZyoGc50EKx+FaHZAUEYc932woriB55I+mn5NfdVnLIhh3kFOt/VRGMO7uSmswidtmKf1oD
S2wMTfl0aZg9B+1WeeKbf2rTH+fqMzjQ0gi8iOTBdd4h7FZucLWo9pkPJG7Nm11qaBPTnO0KvyVc
qgtO4mU8EIlKLKz53id3y8KeB0iq2zgmHrSwojTPyNvFm3HHYcmNG7adAn3+/6I1mxX5LhWcVFUr
GXlpYy80aOYlaD+3ucgNp4OwN3xYGzi+fDSiAVr+YK7UqqaBZku55pErWMDZob8YloS8Wlna7S5Y
GLO18AcUKau+0lbjj8gkz7iSxgHjVClf51pGZ3KiOKH9tShuFNzNfvFFYcI2xrWOquoLNtbBnJIy
lh6A4rn5+eMKbbltFnnAdvAPmJM4qXYLbiVYWXe+++wwEqrvmjtKayeMb2w/bVCYqELMxvKqat9b
Mz11A1FFelKoOEukWjMV+kljcH/r+4AIThg0/6gD4Gh89Ge5E5CwmbsqfZNQPEuSzT1QN3eQ/9kM
TbJCBivjCGGhDBoRpbjLP6TVI9mDv6J+g4NRDKxLGqpL6e/nqPMF3zgcV+UmUKCt7obMRy8OlqF/
OEOfCGVTbZ14RyfYkPUIO4FIblpB4dpitjlgh+qd+B6C/wjEGBpA9vNnOqB1k8JPTJ6YE0c3jKMg
RdKL9/c37RjSe23xxdpQD5cyii+rFO/vPAlWukRVl39ix31TceRuNEwBAUVFmY3EAPoPXSRGgb2Z
Ha5eruMJi9pyoN3Sl0w8rvm1WQAFc85DUDMWlU5ZF/3SbT4zlBol0++xQErpehIifTktgl+zErJC
0RwHCFqQCUXysQLTb6jc3KoQu8sA3NSm2hw4YK+M5Dd8S0lBi03y54xXGPWEFNyQKq12gjYY9m1n
BNkD2nuqpHCb8luQjOWTljtlcopB0FcFCpS/Wtva7yfwfxS7RezBr1QTW/u0zUs9yikstJxhTCkV
CApsNQkGhr+MTV7NRbz6rNIWtb7MEmAgtRyVv2J90JEU6CRW1C0fHv5N/Xm6djrVpe6016roWY4u
TdCENYxlo2vsDexRDLTXyy5ppF2+UGBQRP9JDswB1ckxRgXGB9ZZekkVcxsBEbSepiqVO6IfJKGL
sr2jUOQiW6amxh/9oExHXYdQnr2of7rP2/qwIn5H5ASc5j9zvmOjIZLFOYDP2CBY6uOGzOCv8utO
oZcGOafRABsLWbxfqAUaJfJkv+FbaSBdV9izn5ulr95hGW0AuC74Q9Kb/KE+bsM4L7loEfopKsjf
KbP2cRDWsNFuD1rtFVrf1bjk5/MoSlcl+zGC8wxhFBoImmT6LGl4q7TiyXIoCemq/HK9zH/i9rNC
K/L7DitDtXCDSci1KiEmLqWGMYqaQoued4JgcXXvvrLbxssu/W35iLrRnwbfInHX4NHzX3ymTpRv
Ffmr2GBl9RwEdvuwCk1O6kXkSbWg41fKoYLKDJ15HqjYzI82tKaNtPlzk4BPELGECTiEKpdwPp62
ei4nX8HYVMCdoh4crQI8HjWgnqg8FpwHBrPR/4tIsZ9gehAI+/nhaETN1QQvtbYSKv6F8fsbNBcv
nRNneM5UCLPQ52iXALgs9zuQbwswYybr0haKSjcJJACyJmcGp9KorAtW/4oWVX2Lm8yPOTxyjwCn
rJFM0rhd+6uPqEnt0LcvnYT8Dd80z3HNVEljpXqbT1ezlnAz6dn/0qao6YdUeuJeSaLCiOd0z4AR
ezFYkvp2IDeo8mUcgld80/FmILXnDmXPbQ3aU/NhYeMGJ9KGbZ+WH7PHfD6hubHWKUtUwibxc7Vb
FM8Sa6Jn1CVxcBF8HRqN7OkJq+iNP8zzEocu/Rhs2L4YD8TNr1Apja21FBwsXGMjeYr+ZL1BlyI2
3CeApyfNh6/TW/d/8eg1hbGrNikqWo44M24U/vtIKLCq6ZP4fi7EY9JT0KOfxM1ilofpmhnAUa77
TlYpvP0KFIyiQhqIdCargtcqrIrTKqk3bcgMXrgBWSXKB7qQJ8pDHGgfyjS2X6oWVWUiFSBOaI67
oSVM0/vFHRmHP7tglAX6iv3HFcFx3dtj1ec2TL4IuW6MZT0DgYzppim+yjneS4HRilElO02D2i6m
bPhFKYnVTymw51m1ZMzZvn3n2EQlolUmHzyfMz3JtHkzSa0ZzAaW7plT5Rsbgp0fJPEia8y5I1+Q
QGV7dVTm1olqEd8E1t0olAHSqDiPdY0z0tCEz91bsdjpwpc27aucP5FBvcIRevwWgtNogIOAI3oU
Lx75gkeBPf/VNP95ZD4DiMiVZyewiCtRgvdg2RILuYRn0+XkQvuLQNg0AaeiLm1sBwRkJdsE6iPy
d2sd0KN1eJT2QFXbepJ3bi9v9nuxwLtQUl9vwcp6s4mSNMpcgD9CC3dhxxie1FCF8LPCuJH2+HPU
JiaVlgUM2GsHXNnHkvoRql+HwTSaO59O7MC+eIDYaxPnvxmh4uIxWRziRAcnoGc91tlCS/Zi/iX0
RhFl18UtYJmBQZqNtgYdXw642q3ATUq4z3yti5mdNAcPfDpE65F64FR/0NyPnVn6S9OtFN6Z2iKu
UGUrKnhbLBAaM4U63TaRQ5UVeoqJosL7ciMmQrKAcoTMdDCUcQx1qnVx9Gk1ifGx8LOXAI2WeFkg
a2lW0CDwkude6YOpn2+KqUOOCplvia3lD6ToBGO2pbp97SqsZu8hxvDYMBwyhYNl6itvS6JR1lGo
k5/+2V/BPnKXD6WCL7QaT7Y0gyJ4+EVhdLRe0FAeBcAFPSEVLmOXy2pa8gaf2hkE1NZyX6Oikh8h
YUKd+86qsPpIfmkJLpgNipZY+BiCbcjsRIqRV/UZrfCCGEEilyJh/asrxt4iN94hD1snYcS0m68b
nO8HQ4GDRpfDA0fFe1MZA6J3aqftz49GNJpuqbrFGlAYEq6OWdqIosHCDjAIjD3fTwiSW+IOccnz
jCdsMN1Tl2Qp06WeufRjn2l6HlfgutbJU33ebLTGqxLUyiaQEsd5CQ86G2phcKTizUpVLT7PP+/O
Qey9stBFHjTvT5MFFXEUwVAkbcviktxcVH5mq5gJwu1XT/3l4U9Zbh6KrLO5vnRSbFsfxEIXn23v
NDwkakS2Mw2LddlhOkPbhEppCa0BCA4YhgvHcB59S3xZQ/KunA7ijyEsycURXQWbix0TodhTdAf8
fBwWhiaCBNEp/4QrJ6uoc3+TuqCKsrES+ZVk/pPn5cK0Valkdvh9PDgem0zGHrXzm6ieFl8nNc+W
Flz2UimVKvraSFxjWryf5x0nkOZ0xXJdUap9/XSSabbPeP8DhQGeaejwYy7ZNJP8wsFn6jIiEEcI
DVWNgiq16U4pu5xG5Vlfm9fb/YroejyyYuaxGZ/abmeCvXH9YFyjIby0CyRmxyMWKeQkkl0WaCVw
yAzYqqHraL3x2lXFUxYjU5XVGqTW1nixKOagBQ+lj4Wqex/HXGIDBFcUzsRlgNhkNNWHSiBdyddE
sY5c2EdNFCIhvCN0KW4U3wpNj69u7m04RM/7Xz7LNbBDvcKU71MSn0N39EylOYsrrTrZI81HuEj4
b+UrPKiF8ApCDKx4uR3jmSppMDfHEKeL7SJZdvXfyqXtYYAPzg2z7X1Miua9fQU3rGIDIpQIKpBB
HTcvxiKBmUBqMkgQjNc80X1wpKGrd5kv10dhYYiXiEoUNrNUEzjHDYKK1n2vCjh8bfNBTdKR6sm9
yF3owP4XCVwrO0UKnL0mW1M6vD/9vzJ52bXry/aS02Vgx2JnC3dqZJVUUcTsxxB7L8sCuC0P/0dY
sEHLW082IzetfWNG8SD5gvFquPUBEehEn/HQ+tQXhpUee9bMZ3jSkIZUsj1BYsSza4UOXBWTbdBV
3Ccb2qGx4gwNBuw93m0kRK+rVoe4ZHdeGSOYZ9JFj3pFN6/jSX23yAM2pB9WCxk1UynjMJT4Cnpv
dqyVbTqfm3JUv1SwFfP1RJhBak7QmGgkwMaSC4hvQMfeFeZ0EKYj1jZntobdbPnj/Tvad1ZGcxQ4
0ePGYMZ0PfNAZDarUCdH7W4hro6xKE7G7m/dAS+fmcaxb5BENPX6ShjLbvX5K1H45va2qROOQuMS
dlFE3T5q4dXVSUk/eC1CI5e25kQ37CXq0+Zk9BDVePzB3rd8uf2LV6j0zmburjY05+BYtWoLV4KV
OoM/YcwdL5lX+YilrnHG28TQU9lOGyofWiEYaw8YRqvXGMIdHANN+wXCGpniSy0xRNXIo0cT3Nl4
BE63mPeZo1WmN3lp3RXrPjnN+WEu4eLZ4gU1vKbOMs5HJdvPECbRF2H2sVm3+1vS4RpE98E2ouwj
gJzH2Pui4z8RWOREerup6F4LxIZP24U7r+iqqtl4CkEo1rYeX3oTNeccK/zi6dsiPQmY2op7JikK
QKwhFxVzInvnIBrR1xz83BgGCxyJJC5hZ2NGot45RIOCIHB0NpHQ8qqtktNWCeux4SARb+cw5eW2
S/QM07vPuurRBKeLNkdIo3hDrxgn77+kLPN90s8OTDZ2zMOgbV3k0aOjTBce8dFBHXbWryU6F56a
BAmKJf2tKx7Ymh9mViu+/OPw5vEfkf002lA1ODTZumvBjHes7uTDB+Dq5e6IQul0A/10EEdZjvv9
VdzO1BqPTlcvQWPTxJM6nTmBY7MbeNWvtR8AiczZvKr4bhnU7dSIa8BgGvcSDC1umSC+EKXVOHxO
HP3qdIGG4ftbrkZ0inVRNLYmXzS1a0OFkVNCwAr/VzzNv+2lbZHyEZ2ZHpqjZMhOO9cccAjBI/mS
SSzQEx/KJ4f1TfAJm0nJIX25j4zIns2mE3MddVkCjPSUzXacka0K5oOQcMclpTj7tFW5tFD2O4+M
wbGVZbucXLwx6ldBGpjjg6Ebu2+ihTjAi3hR16LAHXjrAUuTnBP5wP3WTtz9SCvorJo+I26VwdJz
z2vnNOscdawSk0R/Ls67/ZBBp5BRgUNGKw2xpJjtwvHiy0int6SZ3LOI5F3YV4bb39xt2+c9Spc6
nvgewazaHyAAZddVnIb2Wo3CFiJgOUuFvks2BrfNIz6N2JpmM41Fjc7gr91P3qLNykYHug/sRhY8
AEgB02yAn+3oTFk3n7WlkY2Q8jBp6F4BXr9SE1AbCVl80UoRjT2XB3+IXwG31TC0he5C2d/zz+ot
2kje8rqJSECNhNfX36W19jyh+VgmExMD250F5sEwlp0aHj+OI9MuzQPa1r9SOSuTq4+pV6y6IOAR
v7QCz8i/EZD5S+KUJwzQ6XZErm0S4Uu4ESInCw2fQ6YMCI4iDmLftN3qhZVbOuBYUUqzmtDof0fV
dzn4g21TF04nAkB1RSHKaT7O5F/UJXSNExLS5qXNTzmVpbdanghCxMiId4Z/PvBCsYG4Xp2qoaqA
j2l0GXU2eNLxPGcv0UK1c/ogx8dZheJwwI+4AloeOnXedSBeD4N7UE+ABpqAj3xGyOO0g7oWxAqV
z5qSGHL/fanhJlJjoarWhCovTCTm7ppF0U628Hvq1CBon5ATGmwx6B+lKXyXY1WX1fd1DjcUOLB7
PrfNW/x8GQXAZVsR7hl+MkUauD1tP+UqnJEFNdrjexns4RIAU0bWYkv6RWYQDKUHTlSqdXEHu5iQ
eGWKM1s6/Ti+VtNI32JidUXHkQZozJIQt6BtnOPOKg17A+Hw9gaTst/R51xVLoQ/mssi7wmfceff
VAEp55FFaUUfp0jU8eGI1cMdEwbc0J6EAfcPrj9noVJEUyZxj9CFOIE1LT8DAaM/fhnyJTpbCE56
1UraBM5ZtflzWe0ORqyyNkql8kE+lJ2uerHgOjslHQ8nf8b/tLaoeRyqZwwP/LXMsfHgjIEdhaY1
oUnV9IoUQOZZPVKXQYrs19zz+NJCMri/twZzaxRsRok8E10DSPFK8CdklXy9SG+Ow500UG9ynUBz
bHJ0ppr1aVt8g451hG+qdQ9TDckH5hFBMaYYRR12PWOJO0LCWVYElHQx21fMgzVwdH/kVOLdXXi0
SlcJi2yCqLjxGx2edsi2U0LLTc6ciuwkCZSjK7OBTqGG2RET5s0CmfQ8ZAwoFEEdcY1b17LNhlYV
qtDWSCdtc7FLLRFYRpXohkpMzt7Q1nloM7PX0g7MYgc5ik5zkgZif0PjCzUVN3BUhtMR1rS5J43Q
bNXDrPuB9kQCxgc/8mf+FzEzELqkS1jNRSW8hwPryvseFhh2V8nYcLZjURk0adxS9MwKF8ZjUc2U
w7EdN5qVQp+/FkbggCaJCavElp/ssqDfyx1rFsrQDVxPu5A5SsRgWiaojeju2lxZvbtPaDipgUYm
XtPPfUxmH2W/3UBeVNDjDdkbzzp54ucUTbobNTp2NY3rjoUO1ikhO3mVufLCf/eBj3GRNUhX4Dov
jbsMynyjobhjREq8IXZ+DGiJRJiZTS81l3napvD3S9eTaOMVqGKWgunOG3E3sPm5b6aOinyUFLXF
EmDNJy6AtRs0gL7xjq7Glxkx3OdonE1T8JN2xBr/Fe88x1NraVnlFfdP56Rno7oRrOAnF5ZhXjMo
IHgbXMe+1zfqmjcA0nbnRYvtBsCtWcXquQGuS89qQNUpxz/PWwL9Ohb58ZAtOQSnhIx/iJ0KQeeT
H5SqwA1UXsvMFaRdlzWbv8apjBmsTjlVuVR+0BDPocdEwBc6Z0Uwb2RDkDf2+znGB+lX50aZ+LHa
IQz7ooAPFRdjHomZ3EzVcAouHvlMToncUeF7ol8Tf3vFq3ufLh8seHu4cOlzSAY3gOZVlpqrO+9K
AhvC4DWBuf3RdxqmPGKM6vdViz3NlsytnEutQp1o+BUDKBRzGzQTYRZxBYuKpZF2WaldWpUuduU2
PUOGGYqvAzFNQT71TYWVJD/DykDRNfBBhDXSyzs9Yh8uQ2eqaMNcFCZEIhctYmYekF9X4lRb0W91
BMblepUnd8TWHm2+guVhb4SHKSoBHsj5GByddx1oBZ4m6Nyy4H4cOZSaT1DkExbnFHbSG/8aY6Ao
NJQJ7PKU/gbN4iiPNb3qlB0s7H5P38uONvCRSSNcj+Zsg3UYNGCJxrOO+n9ZABzWndSuRiRRCkBC
Ka1AO14+nFr4LQ2kyTavV0+q2o2TT/dZxsRAgqNFpA/2NKRH6b+uOgXdhAmeV3Bau19R1TA6IAQQ
STwCt16H4OZwH1RcNAIYG9iqDPHVzoK4Tai7lI+mlyj2JDOTHBzw6+A+qMaFOJiQWm8ASy42tCQD
CE39/h3IB3L0g6UhBO97DtJ/TJp3hj1vl1LOKcg4+ojZhy1YSisxbPSUYokYHGnS2bgVNPeLfkFr
T1bl9/UOgEEjDFXmvpVSjrKIaDyVGL/X7uzJJAesNyz2F9fW4TRQNMTPxNPQ5ysidEvQR2CnBFhU
Ua6GFtw+wSFZsY10u+66E8IfEloqKGv4mVqBGyu1uyMQG0dpM3v34qfoMMAfE6Mk7QlPyDD2MxlB
SZyqowSG6wnzwCzk0hT5pZxcfLnJCroVM/5y4JpCp8s+sAnMIxekgw+B6pCRpKvOz13iJ+nuB3SD
eC0cyUWaJ1HAQLIoKgcPkVIeJ7CS0FXXBsNHJawDUa/x0LVonLKbY3HM83RWzgX4G7HKlMmJeD3D
5smJ//lr8ap1mfqx/6+PL87kCEJxRZpyo5KgsnZhQaFA08DOT5xjWlPxrO7PFUf0e6qut3EcQemk
H1/uCgZvzzSq7n6vuUOSRoastmSWVFTCPebhModU5w6wLw5eUn5MXKfD1LGRluvB3Nnyt0c+h0Gk
0F0aMbd80RTzkhV7XRtjNl5Xfg+4EM1xLSX8wURnHNhTm+ihknRqVgCr5z0ThT4DN/saiJCklx+D
K3r4vWm1BYj3WBEMaQ4lzSBKiYOFZFMgeGJRHz0f49k1jj5Ki5RfzgiIoy81p721t8lYod8zUdZN
d8RqF08gIKJgDHPa6H222HsE0L11SDpPwRvsyftshHv/K6/w7/IGvGia8gNIoli5r26XdeFJe7RC
itluHN9Eg9mXE0dIP6PF6+ehm2FBHy+FmVe7asZBjEk6MRR3v5X7SIAEXmhsJ0OCB812j/cFD4jX
CSRuvQhsqlUHljkN5NBdRovoiHONfD0amp72bJd6HDK150/vYiXPctLR/RrhVJ1vS4zo/gR84c7Q
PoePNTFucfwo+JF0eSkaNoYfQTUwSNSk7MA6ZVjy+a90npGDHjbfeTs0auHrKN6hY61/+jInsk1z
s9d5AtNTIvUqCVvAEBemQ+/78DwXtIdBq9iVbI+8eeqfQr5SFAqP/baPxfTtz812MrBplJLkGda2
s8Cci4NHeKq8xWc9+FsC+fnEBw+jyq/AkOkCR4VJxHH/ZvuBPS8ZQW0x40i4MFM4h5FxXM7kMRuT
zNd0KcyJcG67LqmK47uZ1HxoV5xogXqd4+HW1O0CzRa+DHN72/JNbGjTMgaTGzB16OcZoFivQGjU
9F3O/a0c4aLqWuA0uJlDTgnoskQJSaMS4CX0fJaOS7SxSqwc4no3ItB8VHA1DaUgdHimuh1AY+pu
o8WwEH9kcu21j1LYnq8REsVgrgUvJBIWvZf79rdspiUybOxJU6hLSOl0kz8ZSBi7z+8P0ktO3ARg
ydkOddRnMgGvCknalXWNaqawxV7aEa2Lt/ehxUJzbvVfGFJJE+V+vM+U1v85SqFjwjMsbC6LqTfb
wyC5nlg3B++GY9w1bNrrNClCONfhJogpU87pG9jGA7ZyJwKZOXYs+Szney7EeY6Vfabg/Ue67XNr
3ELVPh4hOGxnhglm0pBm1Nl1cVzrDIUqCNxcJroc66sE1NPUy98extuhuY234yawpYmi7Ji6oMwX
EVLPK+mArM/00STmEsw7K5HffIK1G9/RBa4VSqUj8HPIutsdX4LkMVfzWiiP/mMQEtZBvzKOqEwm
eI2Ke1Vprsn9B+Y4PDdeiYjz0iGL0wkGlZv3H6c/xRptUZU6McHYy7SiVk779hiVbMZf2vFjHFkF
1CkkbOyLhTxcSwBHZW4WINmrgDXTdDlytrL+ULomzg4uDYxMMhFtoiEOpYI9R4A0B1BSyqebrJ48
E7KlQ2MdRIHC27T8Dk4/QdrffBDgh9zNVa+09CX5fLm1EWS0+DqbZQrT2txfjpM9A59zMKqt/87t
vjmR3NEEgz2cMD4v+jgD73MxjykIbF0ehaNBrfmNl15O3cN8Svf5l8ALjEZOcz4g+0WcUj+KodHd
LMWMsxId8EpAap965Z4C2ng6KN7cJ8/89TpAfHoVZ6w3k3HWKRk++7/r+l1zh3IvMyZlj+kig5tK
dv6lFoG8qXWarXGN/dK0AN66yFM6Zlp0hW1VXV0xyiYA3mRoSUfvoV2TyMzYF3J7fsjWLg8dvgIz
H/uI8xSZm3LbUwr4JRIkbgCCxvkR8suZkM2z+7ekal8l8wvL5AH2GVvTzJuPpqV66gkOjgAkXv/O
H9sG8YpLo64llulWiKxPnBDEBlYqr+puXdpC1cM2JHA9yHiABE7Ye4F3SG9GXdBIzAhMwpsA3zav
hkwXf54tsOJsT4Qts2TRVHxkR8LZqZiI3kV8fpGzH5ImxMtjUAnWUZnPPrB9EFQmwO3+JWDw3l3V
LVkoMdeSUHKfEEs0yPP2dOJ3CwbOs+6MNeQU/7EfW0jPgX+I9IKnc5KgbIMN5c9g97fcex+sZT7d
8zCEil/nUdMZz1VOxEOSuX/GzzXL3HrOfO+2AhiGKN9vWuPcjTid/ZT+C9VZbxIc7ZVF+aemGWSo
znef58frTRxJX6TPaot8krW87nhmGqhLfD35WUahGj1bMERpJdzbhdM+yCQSPKUBZiRI40LEGzNR
uMQgpOJk3DXkbLlLUJeseXK2qlKMWtTTGqfLs0vWHi8IrrsGNLt/b9zezKO6mgg1Rwts0QnBuHAG
OZWOcNRn08ImygAV3/8yhgYTd3paerMduE4q3fd8pAffI3S6poZOo/sTqwrr8BrcG32+G4CCyT2f
il+48qHJ8e0NYkz1zUayWUemTrs3b95Lbd1rvImNt8gO6L9EoSQkTJXOfGGoYQdDoRAlrNE/nWUX
hvrERLrXbZdOuEqoYJIkzJOUW9DYsuF2lMbvCBchyZENRBsoSs3rZsM7b+Fs9JvIE0MZayMwF6Rm
Z3epMxacki1TH/aGQBrDdmzccBfoMRafQa+v+z1fQgKDF2im6ZayTc0sbRzyy6PDAOj1Lvy5ZZTU
jS+Ohuu97MaB3bwQ0Jv7JoydrkAKoa1iLqDSrWfIylf1tQLeP/t4sg5vh4jU+v/OhkZtqwSViWqm
jrFCJ7o/fBcL53nUndF+NbvCSHKwhmx2Tqq43QkrTYhLFUhDaQyl2liaZhdCMb/usHtXZR72vDoh
lE+gJRbIKhT3Lm3gELgmkmd91I28XVvTuQHZkyTmVQc6VrKQinYq0P/5G1ZkEl1motUUJEPPrgym
iofqQOhjtBIxuoc2w0r+vCK2a5uG5Qta4CzPL8WZCDzYLgUD/MgFrBcvHF6Gh0vAwgJ03T6WW/tT
t2Wg1jDSeSJQNmwWVH4nlPlBmRpS9bZ+HT6x3gvdnhzwQ67AbzgryLGePlJFWCu6EKl5lt1KgZCK
r2pfWXS8iFgDmXjqKa3OCZNf6YS6reF9QKCvkq8q3XtP0wP+a7ohHjdEm1LKKWt9uyeH/5npxWfg
4XohKRydElVKECusCtEQm0S9orP2LFS580wmusSVFIrUHvHxEkge6VCt2eCXD9raxQdEwlKTyVDg
2B0uHJNHhZCBogVR2iu7xlQ3LnnSLA1N8qCjnBsHNn7K4uXXIAECrkvrygbhWBy27+8NpiY3Udry
B26+m0CQ3r5IjNe33icQib2OWpf2uWvbdZZJ3mvSimSKzDpXTsLCHOhBfMJ31wR8/LsIWMZVFViu
2s+ueKAqttiB7SiMLJQ1RC6n5AYEyPpX/iwvkfD/6gT10QiB/N5O6Pq0dmIlSKZ3yAr6kcK5u/tb
ptdpVe8cCBpP19MxRouL+0RBqsU7eTPPg+fcSeRavw6C6KRJsRIgo2b94ShCJTcwVTX8xLX4aUeF
avpDitGAiEuaMppnbGAH5S+zFs+J2o4voB8zBzmbUTKjEy4R6onapgeJ1jHXvZ5PgpyNL8l6fRJJ
vLvIYaRA3EtleOSheYgCHToX3HGX1hsijGXZJD2q4NhhMK45tkYron3xFFG8PJRFZFBBYQReU/a5
nIsBc2NAqApiopP0Qy17oDMKExcOkma7WnAW45hLKP1nAZtxS3TrP4ntJ3XDSXwS4nFEwO0+xnBv
flBiDpjUC12zD/c2qufOWOCNp+C09IlRpvd+7Ik0/T9zNuwTM23FpcEMDi0Vy2FrgPSPx6Yh1MBj
FmMXG2L5wVqiagoFnddQR7UksZmmBxe3nVKwG91zay4tZlXoMuOpEnAddXUq9ZDDPQvMwLB9Y15E
Oln7VRo9DtMzD0gcT9UekIIdd9rzHvW37yukILxCkaAIKIzJs2g1a/DeOVOgRxKSYa1NhG6wzUlC
uvgAZYGiLfFjS3Qc/rS7nshNwPGLWWg6ba17C2JB2ViFrkhhKIVLShSadLCRpx3C6bS/B55ecoAX
XKW/vu/JhCmBZnMpt+8/Ixp0+iqRZuA7/Ae4eAjQkeUhiBIUxbjsRogwgluqZ7JNrminEpd9aX8G
j6V20q2v3gW8G4zLr7v5Xvn4l8fplB8RXLVgF+JcpRh33EApcaa7h0EdztrHtIXJITzsEKbPXwPi
w+h5bHbZotipL6i/6kinJgwCezO+JuLgblLgxdSBYZiEf3SAzsAtowERbku08GvLdDhmg3kRi3he
amSMJSFOZ3iddhCn4YH+1PUEw+jcnOt2EjWTCTv2wkI9BtAebz3D7Mt3Q9xSVMsrJOvGsSFwOtqR
r90QAbWxN6qmlRbhgDcuAwLajTygnhOUAs8CIWZ4KMswn6/9PGCqPGl/Pue+dCbxEPjz+kEiT4sV
NOOH5CVbROGrPU1Cx/BRjGWqdPIhfGAv9DX6czksR+kqx1fnAR2jYQB5qVDKHN14kRdANvBOguP+
Fs83fGsQaRZW8Q9nUwVFbtlAEDH5fpIhLB6sYpfqy7QG6i0ZDJk3E4HJunT3YFxT4Ts1d6kZRvDH
4BpOkkDAQ0AH7p/wJK2BctoIakIO5q6u4WoVPNDjVF5NtHlC7ou/LmWLCgKQqkBs4ZPudXenah5M
6UUZWBhG/bqt/2T0khe6WqS9fc+zxnrlf2vu2Nqg+1JCtqh8ozxNfnieEezRWx0BwU0BXoNo+ffz
S+lgWMlss2bYc1zdn3rIIFvPmyFTMOxmOefcpbntKZD1RLGUQ+hLGr172/9EAc66gE1Wie+Vehnd
wkrLh6PZsoA8yhmfrLbcDKWUl4rIV2CMdalxceWCj+Xaq1q41my92umi3h24vKXQNdPbEjVzSY73
IPh7aXICnR/8ot/JqilVcBNPLwDysBjo40S4iK/KZQ8sa/N8skKZvHEDCVJjUUbawhqkU5m6JTs5
NxNJ0xp7mtpwCNLp+JT6iADGQ4LG+3FRr9TckdzwGpnrlii5JizoClsLnx4VGs7vdjcAkXnn+Vva
yT5yNSagWxh80tMxziwUGidGDpAiwP/aeT7PNk35TKunJm2owKFuyob2q0vZ2zYD3Gx4qcYyPIu8
VioH8Yp2y+/EjTPLdgiT3r8hDzcq2Qe8fTmj0twWUeaSbRIDERYktAZ3wGFJAXKZFddNh211rGkW
m8UPKWEvqcU6jKdxjmMViZ6l5M1S+Y9EBhgstXOJGCqwfxhNBlWXdMrn2Pv6+8zx4WyosRtsAqHL
fLrkTZGkZAPTItiLsQk9R6NDBmQTgLoV7yuWli7xS8YluMa0mGLAd8ruR7ztca1MUZsFioED3TGV
/RytwSSaEmDyBJZrD6Qk0psW85V8EMMqf2Pa9gfsAlu4yWYI3vFewF2M/fUcMe33WNS4eP3MjkDw
7N+Ac9YhRbojMvs7eZ7Tlnnbu3/3J68uBCsA3oept2Ywz/nS/kozrM/VrmW0YKeL0SUSnNdJWdYd
6tkMxOpzly5uhHEje9lWZ/nrwCIUGrvmQzg34m8Dq4Ki77RJ7g1ifnBXWlV5HoGg0TYCZM8oN7n5
jqQ9BIupBtBQMvU4qo/KhcTN/IGYag6po5fLxHgMVSOE+O4C3+lA9OS+t3MqrODDcr3MJxcsw5RT
zH3ozpVjY83ZRJh1a9N60/x01UkoDicTtz4nk/EJ8+NJx3JkloNMpX5EEtNldYs1vrhCid2Ty6Wu
GXBrevaP1QLfCcWoKNDMSxsqLZnQS/ikG+JOgtOJJHeE6OZ50HvP+cKeXBS11VPN0OnDg5IQ3CJF
ln+CFm8mXnRDRMhGgNHj5qTcW29s2XWNzZhjfFFJzKmVY9Rgrregn91dEupbA+um1U5FmVFzYwrd
6zQ5dBYewnNC8l2tyIf5FC8tPcdmwo8KVgn2T9k77k32InFHZZWheX+5kT0OeiojA2AA4PU++6Kp
OweIuPMrY2GL6RLMzlhjLTP1AzSPmVvMvXIaEEFFzRwnhpv2bIxQq7u73rtI+M0VXDvJtPWbnDdI
orEy7+hvnYlovA+pl8GEOvx4dlaxWh9boRVFC/5/098JpvhOPNFwC1+WIXjXyLAQVY6NcPtpXHDI
eQxdxb/jydMlF5k/JQv8CI1oYF5O/d31DdDgu4onmLE8R6ehPkWO1E0gMqJDVS/QakJH/CAN9FdC
880P+mESSbUQDtQBDRVAgspQ5vMYROgbyhpUTPlNF8lu4nA3ncQbEwYFmz6Uwp/Tj4FQzmakI+VA
rU1i//jCwO0eYEMjvfol0BuhK0/A+9mkkJJZW1xQrFGf8DH9ZbxwAQ9pbG/eNIBdwfXyo2fcQT0j
EqSmMvqjuCdG08mYCd1TX3IbQqE+UzbtQIp8ZiFr81TxLhTHSG1IWjR2lz7yT6rvnJv6T7tWTozK
tNJQSzN8JlkV70OfGlWer09bEjnc8sDb55yCrZ17OMEm09yLCvqwVPEsxu7gX86BsJXn3Ig6hGPw
u79TvxX3xeEaOqGo9DkTrekIBnxLE5B66+9fxlnBBbtpbrUCR6n/Ki2hXW9O95HcsckdfLgVZ7gs
W2VAwabB1ozrB5xKm+1IOS+61mytz08+ZNLgbfnPyKwj1dXhRt3OhX5GcMMJMToKiHmtm5V859m6
Kzrom+yPxPC+5B9id37GLRi7+CBi4bZmKTeFK/3ty/93Ff0Nr3ooY6cRUuSvHEhwfzN7HX9vDyeZ
nHEHPtsjSqEh44lvefaI3hgY4hbfyVG8ojCnWW1rLfB05Ou9pnc1Cy6inUXcvNGxId7ilKcdIlmy
J6ydzGDhXkrWTU7Ph9tzXlSMoXXuMVksdJzmWkMmY2mwVL/lhbOOC9qAB6RBX/Q5UWJYtDYEKE6i
j6KdVhS5YNnTZvuMuSbr3W99Dm8UBhVe/K2Y8wiEobrOIW6Im6BRF2dUg/XrlfBmOIQBvj/vPx33
4UmwroYivhgII/CFYaFo3EJ6Pbt57IBFrrVN+SRaK0lnRnLHuMvYEqn5WysQ3ZRL5pb1wgLJeWWY
m/bt8UIke3xxYlbr7HOy3KV5qdrf+GnvWaCCr5pcuG3ZKRBnt5h0va0OlI2osveii3EY1Gzf9ih8
5NrrhrveE4KoMFzaLE3BUld01icDoM91bCwcVwIAKGaK3Rw1NDKa/Fts+nrElMrS1AiticsFSugU
7U0iMtyxDfxhZKupNkngOzZnPMVYg8s1I0mjnhxvRJGnebXHqAwZasuh2NmkVwuRAOlBvkBT2aIn
Vb/gBn70BF8ID07wQNU/uwBBGxE8+T4DB6y73xQn17fOo/6f/ZYHOofF8C6t4YJCWpJiaKh1dD3g
fho7tPY8R81A+ZilSvGPOcsWfG4zXhnyUeHAcmGjhPPPClf7uw0z9oJiPnU/N4Xs3tXY5hSYb2Gc
4RsV289PcmzHmaUl5N3H2H/jDAfSOI/OdrmQbavxDXVbgZUPFqba5hHUlp3ZxaUiByw6Y0ALg0pc
Y61SGob/0bIlJDspT9vgQV+AICgguslgdTFNoOqRXxVkWzLWrCSoF3KU4e2OVXkrTVQnJME20Nl0
BFPYxpLROe6GgdUv4dXFx5C7FBE6szriP6ipF8YnQPboN2qDf5NwZekBe2nf82Ra7VUNWV393TgD
4clIQlOfGjbWnz67Qpkp0yCu33HHYseIBa60i37WCxxHjqbY37AOfsZ6jpnpz+tUk6J/f6Iqtp91
1ayAETjO9Wf6RJuTRRdxcHljnHVKUFPdItNMKJZjLXAYYL5egOJtDCAX1IEYmlvwq2sTjtsLJ6qQ
eTNEFdP8DRLN0Gvu7zDP1fzfckCfI5cNhYk9gSQLMoXZIsRN847VkK/wpge+7kT1CF8K1pdc2Akp
Vdf6nBgiJ8FMqrSlrN2vDjUfkdtHNFZViRpffpwAv5xmZRtq38S8VTfHjJ+9G9p8erwYwlFlvLw/
+xyLjYNofMAil2foio/QBB4ktOx29VR3LoCOB9bCnmIj9j+SB83pjcviJj3YLg2HbdK4ROONd4+6
X1ApX6tzpCWu3P2fhlbdGetqjDEXBdgop2rQmrDUxhnr9F5nU2TA50s3zZBYVsynbCJ8rMcYr+xy
l5ny9TYXOjrRu4hx94JHk+iRAzT771IJftm7WVviyrZiZNObm4EifCPc0COV3eD8zpIZep2ihKgv
0wXJTZ5vJkTtIm+2gsJzYu7t8a8Nz4wJKps5PKpm1sH0Qo4u1CX7QL1WcQ4YPqKRqxQlucvpX0FU
j5IHaTfuuZlQp/+VlSH9vV5ye8D/hZEp7kcpGN17LiMjGYJabhMQZFAcy0NHPfQgxqbA7evoqzFF
L11TE7h2S+ExBaL362/TyByJ6CSbo7O+VhOZ5QpAZcW5EbHsB2mfslFQliUtBs5y4OKaqfA5wE5b
/gWCAB7gDbu1+tKewK4seeUtSjRdfFeSe8KxlkiM/qYxa+LiXdop6bNL73GixWfHQIkipXTtYODS
y+juLwNbIcBLMYeRCQC1cFGsmyKn8871lFVjc/9xph4nMyRxxwT2krnzCyB/VSzAHwCXYGbeU1Qp
AJWMOAnJrsBx6FzT8tnrUrjJFq9rmppnelDR7d6Ttge0qQl7yZXZppMSUVEueW1D58yM1wnEcpUi
eipwaFPF4m09Pc8pBdLAU9mGzv/BBlAmSjXY/32az/xxAIHxCOcsUhMWKfWFPR74el578zWhPg01
D2cacPZAhVXg64Sgry8LFb0ZD+isOe7TGGgio2UvK4XZBe6+3om45tJSlnJiWqLxHDp9qdMzcNRv
5ygtC+ta5HszAHsWlbsr29yVqVCa5chvuN3tlqcanHWNt4B0isRxY5cbgQDvimoaOTukiTWi62vT
fttuhV/6Y4+VRbDFJkie8AILSFVwhlJuBc98RmGhOy6wu8K9feddPUVZWo/Rv7nyzVCyqGBPRYj1
mTiaUwnC2ZzDWSFfy+CIPt+Z2rTcGNkAiPkc3hIXytu2pQoelp3RVGjdrbyT+BUF1zsJajXRdqAL
uhXCkdp23GQr8x43awYdrF8NAPHf0NuBJhVwy7tI8aFzrkv/SrrL2LRJWr0Bk8S1B+wTFOhrIQ2j
SzxtTe8mw764/1tg3tzWR/ErS4tdlHGIDwnfEHrnIRqdajzW439PwyHbuGrfuwEcnIDENXKccS7a
YwgZ880iD4+V4M3yKxfo34FB8taqc3Sy+r4UM96/OqI5aWwfoVLB1x4HsN6rPUQWcRcBIvYvn0Yl
LhWTHNNhb9+MG5uISDrOFtJStIIdeDztjBugYpD4tQFR/G7yRD3MmOytvtoQ+jMNjHgaArbOg2xn
ZJCNyMIHUeeTrswSTfqD5ISBifyAEY6Zmy2nS7kFmhnmx2mvJgLX33dfOcjDfFLUCfRQQ350jXko
poEq9Ly3XrHbr+3U156QF8Jn2w1V5kgp+iJ7FHE0wBGjmJZ98aDz0zjhHKqJPzCf/K+dFGRvgAcl
sHPSnGFOl7hGPTi81MseQipQ/yJi8/4MYQ49vCQ7lEyzJpMmlknl1ykCfpNeJMhe8IAtWYRWn1YS
rXVOzYznqsbct3VrVxbAO6ywuE2K1dBNdkknx020G/Idi6o+hhMLiy6rEFyae4lOczdagxnR9/6X
7THSz0eoBYSxuvQXkkcR+y94UOYV11ihVB3pVH5h9AFbVuPJdzW3rLEq6UOSPLqnKSo5JxqKdNcr
PtRZhG+4jlaufX5E+hnK12bW2+d3mWVCqieF7QP+DyRhoJU4efp+zEZ4vImPOrJMvQ34cG8UAQRn
/PfScgSxTvHGi+P8T1DmaSvnXTnlB0b193JDD1p/EXsaZOl8pSgN1ZczPCwhlowMVId8+L9MMvUF
yKh6/WDjUD/lomQCBia+NuuNcDZoPZcXRkixO9QKaZb9xWaspO8uoA+feU+jawmOfhWmQxUlVtcm
j6V0pYPqO0UuHGK55Y4MsTquH+ulSsj5fGz2Tw82j3PsbN96HwXEKbx4QcQf7FS4znu3BjAGDBzL
CvBEDHzV5ai6T33z8JX/JDSqk7lMk9xqBa7zgYBj6pARepzqzUO+KNYAPsKO+qhC5NdWDDzBswKt
04O4vn6UoZsIx1kByJ8szSjn9EsduChz1Oc/dPJT2NwhODmb7WP2N3HNCzO14GicTELKk550Dlr5
E20cb2u/VZWhFNTWCmNgJPxEfcmKmH9NjfhCjnteYF9owO1MN2J8oAKqrNglmP1csAD4dj4Kjt1B
DUzfjxuxNHKPbiQFVnDChtFPQL8+cIJsbqp5/Qofp92L36z13BEmgogkRy2pZysXIJK1U7XybN8B
8kN3B08tOJvZEnl/twqPeRYHAmOaYlDWv5Rb1hR/QYwAwpzGfUIcwWIcE3PB7HvfdNr/iUixTo2B
29jPiEPMIWuZB6yAE7KgbvTrwYXOPmKmxhAFOAZuGLM4JeuO7OGW+4XJi2V8roYpXGAtRHdbz7NC
zlpeSbeWG+b9ZPIOT1K/FMXpfTDmsdnZCZ61u1larBzIDdBW7aufqH3ImmX/HvwEEScBf7jVSSdo
5ayqcb04xmIsqKcAVWHznvgpdPNgGhX3INxNDOkpOPfb3i1tTYXjpAOwnAyz2FChE3+z/OxJXxly
Yx3Ig0I3IhYgRuanLea4JTIZi8+SI7K9tLSHGPY244kfZ4y7kcMuDFWItkYHd7ywHV2AD0bEIHBw
QOeCRcFMqXYP/Qeb5hmeA7d0P8XYvpZAp+DNx+Jeuzs43Br2BRGXGumMRGipkbRf6gHLcqPehV2H
NsmFaFBrUkUD/SYhiRzHu28JmcTFZF0+tL+IbW61BoZMnBOYIYobHKUMvj4+drVjdstebNkrkNBC
Ssjx3WMajQiJTXdHnIXFTlRldlEi78lSYzNyx4QQDpAinUYK0V3w3VWzyvxnh3KDv4YqjeKoqOfK
zCVPXkXK/Lf2k6LbTwhH+3Xv2EQFMwi2c5VOWu8dEDhHB46F0iSVkCH9lfHXalDAwWJzsh+puyDa
Fo+LgMBoRwACQDoXiGSA1W283gOIkPE/Nxnh8lLTO9bX8LjDWeMRIHwXcngHyvfYzQoUE5MXsSmR
JFQC+5Evxobwbtk/iI4wFHDLNQhLfmhzFgvq86wgmguPbNvJ+N1rNyPST1tbb9Nz2K7SsDfESKzj
DbgKjIVPKp+kF/Jq45kBQSgt8fXq6csp658VFJqsbTGa3x481hM8WkYPMXny7q6+GWK7on+vCxcu
dbPyyyNTG0hz15xbs5mX1a/q7u2Db6KkUSNBWV8zwooNc609fo2lm1VgmtyR7OO/E9wbbdsyxn8i
QejtLThQ1EA1uJZxD5GYjOCh7MWzd2Zs4APZQbxw7NkZpCEgNM9Vv2UHyvrLNGap8FYbZ8ZMPKm4
MN8dLEMM2+IOdnchPOxJqD/3lOfD1VTtUpDwQmy4YUTas+LPnuaKtGMFbnpWZ/Dm2jLTq/9VetRJ
ahoTjj4X9A4cfCDqoAGQGDCkaE4fBIvri3wnRfCkcUFMj3JmRApXXMuSQHDs1i9vXM7VdFNn1nAz
NhIGAbRMZ7Wj5TBHG2jy/BdVYbWZuRAX9Ab9QRuA6WKckVb/uElEM6gEzPjk7KIno9gjw5eWX/KW
XggKA8in8BFr2BvgKHZLN16DV9HIaKkwmPZr6vFfqVnShG9rliqTTMJ3k1uVARmpjMvlqYfcFIR9
kc3FzC61aFHF3RRLcyRJMpHzDfIgibTds/zGuR8FAs1kogarhoiRahlL2NAcXifqCu+zW0GtAT2h
bxOFTSvXLndA69ttyoXtAv4E+zMCZ+2HNBG03sTKsAYVN4V0LjTVPhzSwqRfB0IbCm0ijDl0nbXj
HWbcCETltt1vLN07UVizZtg4GPmZc+0eeRiq8lOfNrMYIn0pt6w6AZD21byVgYOCYXNyiD2/f8Wv
flxlJNi8fFv/mQXDqVpsry3hbdHCNQEOMwORDezy+l8Z7bCmANpJeDev4Zfv2yqKjq5rOaL6ERrH
a/UuRiItLSQdxqEiQ7ZRTS8So08SyEGNNWH3c6a/1jy+2z5C5IEf9y6puxuNR9GcR46QSKicvkQK
tUyc2+8+/ycdFG5GPW+qXYZdocKU1tGZL0QZIseBFhlckOOR2hv1unCDu/+zpgNVIQslrKR/kzSU
sHygMqIdNodNRgcrdPdvxMQkZjJlj1eIS+bU+6hYhNeK82Flh+vEO2lWJsFQrjeEBKXXink19EYT
hQaprNRnUGY867J1oMuQ2YrNUSyRc9SBxjvzG9wOlVdA8VY937wHRUiLgkA4KsWD0/P9O8RjOwcJ
BwkLTPVwnzVpTfm9oK3eAAUAk3fKoz4N8rjnSQbD7fvtEOhZ4wwUov9z+g8KW5p+QNcxctB2efL0
PebLxmBWLqB8LcUHOjE5AHV2Pv8UumPwUzVxBP/12fgwIDMr2PgrGzdSUCr9KG0GpTIAlodQC3Yi
+27aFH0dLA+4yDqp+mpKFMT2XV1AgkXvD6hLVoAmSwpTM3P59MDJ8WvL4c91gnsTEQ6pu8sppcv8
PvFsaOkHrvYdHXCR+6aznqfrrMzwLDGTLhidkqSMg1+QT7rQyJ5SiBP3ApTCRRsPW3PQ62NkLKga
QKYylUBJUB7h7c1frS3Jwjk+XoY/ATWECYxY6jd2Md7Dp8zwBj4I3Trocr/2NY0Fe7XsPRNsnrwP
NwKaDZ2fmtw1jNWyFQRyr9WcQzNzqEdJnmu7zZSJK3q0gkvVU77WYk91NuKf/3BPQWnjw3YJlsuV
cXGKNzajpDtcmRvXW6lLULengtEkGitFEE74kHT/4BcT1cTAp8HimR8L0m+Hxxylr7CYA2hh2YA5
INTcgYb7KbfY9SPKtEOpBcZ9nJ4nvWpF3Ne6pS2eNdNFCMgkXUAQHtSyLHH0vezabWgjd+E8ykf+
pYVRTEeC2wPEr0Rf4At445akz7A7Zro5/41lATTn0Dn8w0tXSccsprlOaPnWDc/s20Bpuv7BR28q
tXR+clHBisOwEEGJhUY3llwBGneiJSlFKdaaWweIbYJrUvC0mN9uIEgZj5wC8dqx6gSam+sDU/BH
zAkVL/MyuyHZrXoMjF6vMK8fDWi903UutD7Rjqz47smSOatnKNr7aZk8MlhEjBVHgfXNRdHYSOJu
T99hyqffXHqdtRj4bt/2/VfJI6YB0HJtIW+txmAFfcAz3JJ1DbdxDlCWHLpwL03XBwXhhS7yoXsB
82KRC829jDMJ0DGrtbjH11bUhjKBwvQYoy5x68aJ3nF3u81ldFy9W36kBTqLD5Ha1htzsMIpRKVH
3IomtiT4J4NKc933nwXJ+tBkXMfo7VaW8okUq2uN07tMhaLeJtxKMitwqQRID8FGp7GsHF+GaaBJ
TVtYIt1v6B8RiNd7SR2YpHykMjE/oRrCMLSZ+k7BJ/jx1UWiC2Wb0eS3W4xOoPs3h5UhlJn4pQWD
+DcBUOjHPI8eVlytjHbjGcctkvUrM6pqU5sqryxRgfveBZ9L6IlakytmukpZDZsczivjlVZK/Pz8
O/bm+kWpXjAEK/A2tV4mbniUShvuO7c31CEAxsXdJBYb1wQ77dR2ATIUuCHBbmywSW5UwMTIqTlb
iH1gHDTa4shAb9M8KtJwd6NTwZdbn5n2jlcwaM0k+KTkOMuHuLL2OyEuOVhsvDuERItXgcYxZFi9
+68dgIXrvWF28i95+qwySura8Mqi/0XdszHSVIASUOEtLVy9ZLchQbqGYD53rQIt/6RYlIPMVqK1
GAAGa9bbARFwgE2V+MrgoZnHEkA3s5ySji9Zpk2P06UlArej9BvQ/isJMcCu7BvtuXo50oNUPNXE
y7KXep1x08skJY5huBKfVDrGVH/SCMhc+MRXtSLUXase83XHbZcr8LZI1DaHV22fSp5zrvltqIwn
zy7l0L5wwP2uVlWdyrPmqMKQL1FmBFmCTMju0Pcu7W818HcMLIsaXKksKLZDSlO8UCabaL7inIcA
2rnekkILRzK9u3CCN7H37Ob3Lo627HRe4GCUGe9xLS8kwuCjNwQDyl61WcnFmrC5tOuAanDjMK/b
bHgjODz0T73Akf2nKbhRkODlu+wbJMh7Ab4FOesMwfRYcs3N9pAhrG7TuZVFfxvTG4E0rBpbLQjk
bmMbmEXMdQyY5bMmorCHPOi+AwGz382fmNjnjoQcpQgwngx8Txc7eTJRyLLmWrlrDLZ8MKpERJcg
3a2fD9PlyGTN4W9CpXA8PiOGgg+KqTls9PpYe5LCRG/hqJWpjCW7ov32QX38nwkx1EObWuhurc7f
M8cRQjTc06kkm5IJwA4UoiELIvtgz+M2cQ5C18n05W0qoB/9Jh4xo90IS6jcLj8zHgVVRoClIsUM
b5/1t5HuVrSX1aefJ1HupqyKqctLBWqo80zGT37DYUv1xe+uP1pwGJx44bXdXRfZAdpaDJXAjzhU
KnvZ5YzUgbK15HPRc4137tamPKyrj2nhLudsNEcJR8oA+fC8O/jFbxwvFEeSZ4QciyTlUZIy5eyT
jLmNMZ+1HY+6anKlMPW2f4s8cR+yUxQG//HqnZShSDPJKVdndescv2VnJtvg1Sp5nyjEW+ESaokd
vXmo1W4UqFBdaTDP6E8NLF01mf05U4tdWsWw/uWQV5zgOn64z8+uPb4oDeC7c/FbFjw+lzsb5yRg
xw2mgFNFJGHZO/lq2c8h1d37rmu35zNrBmRXZsv3oJDbVW8MrtuAelwKEDtgV5n8ol3nkAIWxvFM
2FHN9XHENfV8RWx2Lh2Q1IJVHOmigSYngJeTfLSJIRbiOb1RBqLZXWx/CutKzSVECNp75KF9sB4F
hc4HcBxPGqN742QDNhLjUDHl4vYVZK4MCSEQYn/ajWevWU8k8Ca66aKIwo5aQk+LKGDGPkiqeOP/
eQchTUjNltzanJCZFzUr3x5TaPpuI+MpYARRoTC6z1kmYajOfCp+H+fMo523+s4zOoEFCztuqfA9
tZP24iv8/ezsLk7gLuOC556GcEI9Qzt+JXCeZiu7QwZnvdoL9q2vNeukK2UyQ+TAmxlw4Vc+EkTb
Mj7kVtLwV4JWGmRvPxzHWZwjmZhCuTA9RMbxTksoTRi/ukhskiBkk48NoFPjtmLDvShT2PFl/2XR
GwO+7rMA73lwsYLQ2cP+LwusIhn9Cya+2uKfUP4zI4HgRs3ONuuR9y2CO9A3q68i+nvOlIlDGE5b
EaOdSREVhVrXmaIv+SclKu1yJbqHR8Unf3aOIWyDXcDv83xkn/Vd6vYeddIUq4RgC8h0yIS7jEmD
S/WPXJu1vlj/5tzPW1svUghfjJunt2ualXPAbHCHj0kXhRThsEXnpjfc+wG6zZh78v7P65KsOnku
aSWnlZrfHlQOKHZ0wFSOcs+1lb2Q9MC/09IdZ7f3sIixvDgvIKrQWjrTUGwRPDg0eCWX44ps5LkD
0H+CMTzX842UtnsOUZy62HRfogI9G4oWPF96nimSxT23gbQkn8D1OGN0SuOvElpUTPBeErR2vbhT
g3EYUdXcZ1X4FgJ/Qi4XhTBItEWiDYE43RnjKb4z7h1gNX6QqGLN3JVy/KZw/igtWhveQXtz9cfV
2WCf8Luv0W+YqAt2i0ITseTcvG7NaQgTTboUPG6yrjmktIAG7FhY392yVQhgqr5QmZp6UW8JTtbe
jxNOgKtneo4g2ibSDBBNERF8UC/38aEp4/O+caBuwutYGgLm5xAlNi2ToOP8KE354KqEdyE0iM7V
y7aU+KQvbpGyV8pZSNc1CLH8eYzzYT/fI49BKafVWorek5vH5Ma3L+pigi3Ptrn1KJGWtYw61n8j
eKRvV9l39Lnl3otTmncLOQc1PSkcnKQft9LeE/XtZub9+7YvaOhyIlPl9rtLLtLThSnLyTJqt1xb
Nvcp0A9yuYZP9aeE03Oqp/+jNMqnO7wah/rSLYjwsoQ/ul3MikiMEYSyftBUoImIZA+Ilu5/LuY/
iC0ACLUpzUfq6FSNQMjiwlCuut6X1kHH57d8uVh1s/SjvekKxLZphKTJTLj+yQZvAk0GsnBRhe5o
u7p+cMOPbp/ytEmOhKaUz2SoWCb7Ynu0NARFi12rjhVdBc4ZOgmIELEboC9m8wiprEhWbwATP6di
c4ZIm2vt/L89x+EroYooUVzbLOAuMH3f5aUAZPt1i/PSQmOAg4Xe7PobxzpG8B1xafBUPzjyinqe
VhoANXp71YmbggEZJWXwK3ntH1VBZ93RHEOoqozoCwzE2nKDmEzmBVm6LsGa6alL+qk/ysUv5E6D
USe3KFQjl0yjEO5btKyGtw55foQ7UTqB6cIzk28F3yKAU+Fs6EcXqQgiolNuxaoeqvPcRLrGfzg+
Ds645EFZWw5/laU/vDcJweGshW+Vt9uXYzHebDsNQnvyOY1OKsQiOEYsq6ZC6+QaNt1+rZwNlfiZ
tpt9Op8Z8GSFXLzoN9T/rPBKpOb4oFF9A6S7yupaTD6HBWpKBSHQgOk9ku16RUvV6sw53DecCORn
jEMET5FLxx7nAr8Bdm02tfUl+/XKz1zW9xgxPC15DsBliwfbx4KdIznlX9JtvZCZAI9fnVxtNfie
dwL2F3XE8iaAAIIFxky4NbJfsbEyGtNHkg3yX9d0pOdoUoTyV81Y6+V73aWvrv6A+sdvRLabpE9w
Kqoav1TG1Q8SKFbHv4/e2i3e+T64oiCfPr0/mG0zKlWg3zdalzJFhm6qT8Lo4izt+BVsCxReMliL
plWvK62pPpSSAXvQk81clIL4H3eRSTruYtykss22M9TkFrmg8RPHFP6jS0jCpBdqq5xZp9XzpnRH
nEx1z0S1ja+47L++XQGTeBS31veg3IqRN+/mv/7av3gAYprX1EdY4BclDLBirDQNpioXOg8/gObi
NBlHjoSTRhIJ1nbcHXW8b50Mpcjp3IegnKMAPaSDGNrSUnwnIM2Ta+ZrMqpJv+hOGh7wX2e6F36k
f29EqMPQ5iFF/T6/vkrS+uZMp/lQTOtm2VeWGh67SrFZpih1DwV6Dk78sSXMzobAYTqE4S3BDg+6
EZ32ziFn7k6s+a2Db2M2sObjVpOgwDb+UycWfIWw1kSsGcafEB63SZuBpQJg6ZuzO/ju0mhpK1k6
2VPV3pQxJ9642n7Sai6QX1YiQcV/HVhKm20+cQY92Lu6jRCLzUFe3bDucSVk8PMvB+JzGt3nHaeo
qhNpQZQLmffl39wobw97XdXngmy4Gadj08raWGMJj1eamcrCHgzjSJqJiT4KRgeOXyMw6PP2L8yV
ZjP8sgeCxUHs0oRUD0sQ8W/h5gU9yi2osI6M5soHEx4tCtbFQNK8g7avvw9hirMo/46Sqczy73Kw
4Y27/c2oaE8rlzqxV/ZwMCb/ciNe3la0CcQ+bxs9+5F2fTBSremzn6oCC5dElLbqk9t+LoEc03dO
ubM2vSzLxsFxpPI+KBiDQqKtS8fgVu9jAr6eSMbZl4d15iR+go7n3yKE+/omcirfbL3kKu+IQx0V
QV5l1kJTzF0EmKQWOzoC5X4o7Lz/C7wXxhUWRcUrJN2vnrw2UflduryjgyD0VKCQX04aaPfh4jVf
8HDz17GwSTOXkzj5T1sPKCxonV7RxRC1dWbbI1I2coe4K2jZ8XHyKZtRVXam8VmnnenvzTaNYNtB
WAM0nf1gEu36KtzrsmY/PoiczANcVAVu/7ra4uyeoqp0C3umnXW0pY617eV6kt9e2BXxgk6s3pnP
zkkeeLeAALmmEcIslMye00FasQkyRK6ZqINqIy94H/5lPgu9125dx3HBMMV39p42w7FLBejRnOYU
a82ZKEa/iQH7yvNzN82B+rNAt0GjXFgb268ENyMPCROC/wBzfDPW1yUmr72fxT/unKlQWwCK/SVC
C0N+LCkzgbYakjc37p9WuniME6JGAFhnjuclHcyzmFHDauanuJbh3I37vckVCkpx1PcFuNZp0dfo
ulJLvHH6jOEEfzpnJhfKYPrPL1Jw5XEnBl93Hotz+MWOkuNhqx26s7jiU/B/ZWzI1R7qWAHhU9zG
VBg+ieowLAZI9QcMDif7drOBo2EZXK28G1eAe+Ldp6LS5qj4dXcT7BHvvQ/hJqsQx5dQRPHYlah/
zDcG404GcaR+jAb5YGCqzDW4gyPd+hS9sck5Cxm5fQ1UctZF/V+xdwr2SZbbISzre27ZHqQxfIjR
54LNwfl3VlCWG8T4PBbZOkxxRqMF3x/sQhD3+5Qo7kWqVNGexvKJExbmhl91cyJ4FIJynggcoCpe
NQHccpKkZVX3+dpxzEPemc1argfhbzcDErYGYz1J+6j4znyjFy6RUSNpP3+i9P5AtHQd0/Y0CwgK
mR56OhVdUrLtXgDJm7xvClPOwAhLkfBXyKHtDTNZf49Y6wbs0BnLfGwjRHy/0dr6DNoCZi7V2BBP
34gGH7gTMDDzJXk9L/g5W8VGh9fMtgAM/dh8UcBrv+fj4HOrnuU/rSx97JKYcDU+A9WI1AuxuYIq
H+o5jamQiKeeSAKzhD5vUwIQc3P7gOqRVFfhT/n7lAD0gVpLXVkyGm9e2MgTFRiVNeOXnOvPuoTe
xJzizP0LcivgxYDU/1hRZ+TC7K4KeWSom6p7lf++TeDZ7F2v+nuDexBf8m1DbyEh9VuStTGP2oyR
dImIJNhm8ZJwyXesfSqJaW0y+qM8QzM82O6Fu7i8QKsNqF3mywNW0Dnzq/I5aLjlVpTOlbDNuJt8
BrXaApBqCtGakx6hbR+vMQjcIuSvl9cKFHua9a9zjuY83XeQpn7ssS4iI39ERG6xmt1JisVos/IV
MUv/gULN8u/AJl57t6W117W+EXAYIKAnGFS/9gRH7LoHPaaOniRb1DvIjdG5kXCLxVo7GwJ9cqiz
2SJIOKvwWI6rvSLi7FI/JiAKEOlVOkr2w/WhahDh1DnGd6ue3J/dJIpxwY7U1m2jXs9h0TBdRxMV
KObYSDVh0JhmkHax6jRDw4Vkh5P9WSoZIuvR4G5r4VGxliSnJmenEyeyC4G8avre7SY1NTYTvFW5
dP2xfkMpBxRFXxapz+1aMWkTy3EpRbnKIQucMLIfhwm7kRenzKtRWxywg747xdsd050ZanEUkg10
KC5Q6xQSg//rd4O15zuvfKQ4w5+djrsiLkXLoifNV32/XaI6pMJWeUK6cVy+o0ZV6P/lm3sP16cn
f2KcOIzrwntHgYGtDxKebCLaGILtuMunvIl7S1yFig9KlS+wnlq+D/aHl94OT06onaXYMrHvhI6F
keKHmHkeOK7xp6Z7BUK2aA5cJbepLxUjWznFhCrdZ6TtShhMSAJx733XbMetLCHbFhCmABzbkmCF
6dKLuQjYtq/Jorc6u4UgoQSDOLFVkwHTzolD5x8evSvtNBlThaPvNtN04XGYl2KZmH3xE1X3sdOo
oRAa3anivXrP779Xz2O4roDAbWY9bqhIYjUq15Fssuhz3LWOy/93lZi3ciqNFcFW+k55zaNaKxAs
BaRxDcAyhiqLKOptogJ+Zzhen5Xzc71vNYSC7HgtntsRW8fQUaiFEnssE6VxOIoiQiISdojph+nk
jQrgPiQvBRPwUBKVaPl7tS26VYQWzOOcowgo+JHdZpypcRlXC67h6zKGOAMNTS22yLmSqDB/h7OR
8XuQ2ljLgCrAFAjKLHz7PeAuF4t2GueFySuAesUPD6WeIItLTJawRxr0zQldsviX50nWezPHv8sq
0p+BYXrnbipuVT54DIEv5yXf+giFI4vhQEtG2RZkiHHULZ5ibk6OOpoDZeDhwk9YMuUPeSUIwWO1
cmkq/gTa9xay+k0XFujmrvEl+1CwCJ/8Ok7TwLUVkSCKkzz2kB/h53lLtWGs8Fc3YFJjCisJoiDu
A8o5m/n93iEEe/Og0nxLFk353c0QFWrL1uHZr+MdrFgFcCdlrpkBRv3g0SnCGPSt21eJbAY3a/9P
VPKNCJz7wVzFWrwLzEPX+Ej8jYu6dRsQUK1PKE6mJWeu90kqYsPAiJfZJf70NQ+0TAyqCPz7GlJs
la7hEjdXcKHOz4rOU439ruCs4Q99s+9Al1DnJhRCCto0CtFdE2ddyKdaa4H9nGZkcZZAtAx0CK4X
kULhb8+NiT5F7HXFtykD9jaDb2rjA6h0QCJtpQDNg1jzGpIM44GkF9MzELmpH9LSGoDahN3ez7AU
HS5K4qRfd9y1/MrZ/wRupwci5A7rGGF37Sghc3xI62L0sBwBmtOd3JOOSHuzY36cBRd2Qe/bwIcE
rF1fiNdyATXxQWHCsr6YwTgucmnmggfH3SvFvecZpV58Jk42MAHkRjqYdZ6ZATlhhLFefa1XJEZ+
QEge867ZvDUarHdAO2+TVC1F/L/3mlWaTzUe8CrViQ3bcenFVHW1AlaryadM2RpWIv/HfdiGl5VY
V3tL0exMLi478BmbjrsUTaFoWPJaZeMObJG8DcZt6hIeTDhXIRIIxgxBMBwIYox7gXxgX6yK6YZt
H3auVqnaIlAsFR3USBinHT+OnV6RI30MJv9o5a3Er7eVJUg/bglS86CNnK6Zte02mz9AbxHJA3Kw
wHqTOGr9ZwTTmeTxl682LMzjDpEtu+5edyawNlemrgZS626g3qq80EiL5ez5kugpP9rCMz1EhsNu
5C6iBqsZ+LQxJHR9FPajomOR0lWP5AnzCpq4IFWPHOljLzggRZzVUnNPX1MBRmU14ytulnCqWYCw
TsbQ8iOMTaltgZHazf+6HkyTSAp0hSpm9eDjY7yvZQxiDT60IK0nEcYfilTp/sqwwct7OA1auxoo
es9lin2d0Q3JOQ6BYEyZC6gOiV3SWppWgezrbD1yY/gJfINBDj7b5rxTQcX6BXvUrGpY0Kg48KxP
0d1ufKOK40Dkl4rzvWkJ6gPRHMX306fDLfNOwLQ6AP8z0+pBIjhmjlj2qf5SfRWGYQHQnuYiG7Hx
cgNiX4iscHBTzTJ2N95lG0deYACJjxPwGjOGlTTr+fdgdQCn4nNsCyZZ37cFqS5QCk3+YbQgmCCa
Mqgm413kwJvENwFh0lkOVJ+SQ2A8MWXT++cB4P8FknDajSmOCRdYe99Q8UnCKhQ9+ZDRPrFucU6l
ii3zZzqlxk7+5m85bsZj95OXYu8KIwz6/RrOFmAMGFTJlxScs3mE7EDeK0xmZdeduNC3chI+yFN9
VyHiBiFMhtwgs5h8KBVt3ztOb6xl+iN9l8Pl5d6R0XgeZ2uvmoppQVorTOC3TVyCTWVjCWvbqnT6
dd4WZv6aF/dPePPxiJ8hL3YfE1+czVwflzAX5zmeG2t3/E0C6qjgxMBwI3nO7QwPsnqHMwcGxsWv
pklWN706HLrCIcr4UTQMVUQNvIb8W/i7RKJKol9Exh9FXjGDIf/+dobL+mRbJNTD5+ef05tH4Oc2
Yh6+cvUU27y8wbcGOeVwPKNznAByxZBfL+sIhY5kXroaGoiKbnrglvVPArVs0YVG3Yyz3rpU8r0W
kHDMQwe7qKg2e79DFz3Ui5+dWb31P8o0My5Q5tB0u8w+yguk5lbuP8Qwffw2REAXFn9x9xvQcvNN
02LmJpVAj/7ST+oOoRSrax7z+Q7Ry12BvR3PfSo7X7CiOR8DED3Yg8ZFiRMlCUCm82AcZcBneMdW
wsp3PFKa5mlGb7i1X9r/xULO/u+clLlTKOYP2DuVcb4t0gqjP5EkqhqY1xjRBO9mNp1cl4zvkG4p
kSy6YlO+D0nbb8pdOR9iEiwL+OBn2xS+CyJP2//8z8dOlMFRZ7fKYvrKXYOqZl9ntOVkelFVlGdA
vGNFRgmKmTw8m4LFykFZz/wPpx4zUH8qTJKliIuMEMQiKn7H4PERyc7oDvDFGMjbSyjAYb4lZCNv
m8mh6e6DmxbTwqOwevG+RNZDr14AW+f45zTiEVgwIioOJfdsCLTou1ARSg6okRhrNLIEi5OjVpxy
lkOl9EDmyXYS/TafozE4d81ylFYA9GurxDRcJ0VTo2SoognP9TVeTenexg1/eyF/bb6n6z8PHiwI
1EHtQXjNb5LLg8DtmDvvVN+IkgfnYKYelyFAXTP2VD5q1S82C5pp/h22iX/Xzt8LJEDsGuuMpH5F
qgyvRFAJUPRYLyD8BZ3zOSeVVmKySiV5CGEf4QdTPDf4bcFm1igGCWLHmEUNQiuctZTTt/I2XCko
aTYJ1VMTbqFZ6A0HVwCA6GegN0DfHahcIka0JKNuSNvsKDzNrAQsudw7e3KpnvWoUIkYTRkBToJx
Rfc/F2OoGvPwqnVOyYwbkX0rO3LZE0PGgJCwOIIjSa3tGX/m9zfENZ15sr92FiH+R87zKW+pW10V
U0371VxAL9oiXoq0YO7m6UbqPqqLNve5UtLZJWuUIADypKhxK+W7d/tmSQdpU4+Nm/WtG7svJ4vJ
HLAH92oAHk09998YlUrerHkkz7/7d1Ojg5nCRbe2CP5RMl5unoAJPkVrS3pQN9JNFa3VkqHvj58U
BqSfQt4HN3XMYYjf7jXXMYbVM23CfueYRozG/lb8K+keNps2HaKIkinEXas+XLSeMN5vjBus7355
X6xgGTCyyiuMpiaLAIiNT3xjqnv7WL5pg5gNoqX6DJ09t3bxnkYv8upZlBtzAV8hdWz9JSuU0ViJ
7PQPdaGa1TL2P+m/AizgJukWpfmlqTxL2p4iv9fbdCxwfdzD5KJIM77PZFa+yDx08p+S4u6FB6Z9
7sffodY5Dx7D64fTOj2uCWap7m//ePnR0wUP9HGDDID8B4DJE2Ccx0JLdvCBOyZ7ettyV6vfBjZa
ErI4zIAz4zZyS3FiycTyrOM6uDuCl4CA7zNLFf3+EWDsEWls1jC80O0IKRpMe8zeiyq20iXqF05j
StboLWgSA8Dgn6QfeSM4I3NpltYlp9vgP2O6nleDk1k1Jtka6gn7itJ4dYR6tWcYZXPmKbuH4sY6
wNzy4IUiqzi8Dd6V79hWZJ03LNjIsum3XmZGPzBVuGbKHYrpo7k4JVqbwc0Iwyx2YRE8R2fe2NP1
78ng7ZPI8b4lUYtCfuKGVhyH2zw8ZhHhcvWUBgNEH6IHttat9cd48Y8HARsXcVwKGQqHRQFq1gel
D+RlQIthYEPln33sn8FreaunrB5py6ffzPN2do0Y7lXOKKHl0iu2x33iK7j+b35MQdCr7JJ1eH1h
8iWmA8KTuLg04Gj+7hfmdzj3Paud3b75dZVV9ohJfMw6MNejFROY1iO6GuoMTyhJFrQDV0WBCR/z
X7EIp2EZeosFoGr3nmtKO8jDrh9puQtTZ/9f41GAyWDyKHTspi2j2RHU80Kt46xflKb3RJInYc2w
fJvnu0kWvFT0iL0yUst3A7pzbIGoSo2iafQjETvTfxv7m9WiRLzH5xnkhT6/K+oGcORb+cygIU+6
sC93dvXEpKSrR7udbiYDMCOcb9gIMce0sjv1G9tqAIlkucsV0pCaSwPTL1+MdFC0ITboxVy1U/Wu
Rhi0jfeK+jOc2SIvWJ0mDRZDJ/TXm11yuyovFqW9OHxtyF684JlcEnAndXgg21MlR0y3VsUU0XOU
N0I3i+DbWW0hcjMrAZeyRl/WeKPzJp7/4/NN7AetyVdGlf8r4fuAr+e8i/1+4hzJ1i/yJ+2w7gD7
kOhUAzUW2tH4MW0DBWRNUp0fzFCOzg0B/KFPewihjMWbdhiCYA1h7RuDe+fkueoJWCX1Zy7uT7UW
kDAkJgzfVFWFpJLeVoxSE04DGMA4MiiZcBivLmxqAA9a0w7PU0BDFaiUNWxs1ZfM5DY5OCObR+Vw
vBzO2B3dkpAnI+GsFQiT1VM6Dp7LF1X0s9dbuYEYNlA2qmEyQW6+0ZZIusF37jBFKHJULx+BdivA
ZHoui0S9vSMZcBQ0JNzysH3mVVYtNFBOtDw5DmUuRu1RNskk0k0BRbhDWtvFE32LA2WvXXPJyl5f
L/HoOXOiaSJcGC+u4lDyaq4fXzFwFnWGVGsargiIsM+9DzTmo1Hw9rQYTfzRzfX05aKqOgqUrpFg
m+QnSZKmqTfGNs7JNqr+l9Z63NxY2XfbWqcmNVd08dFZiI24gHdqm5u/1R3JfnVmc6kkpPRQsYCK
kEjCvQijIzkIRF/nP0d+8drbzTimefQUHVIZTYA2upY2uS49XiqTdehbL6SQaT6Wor2u3YyCZcvY
kJeQjbDHj9ZhU20KvNPw7WXZJEbzH3lmGD2ZNraXn7y1wQwXg8OIvpQckQSNcRyj7fxpP7KmOX1h
LGaDxPJ7Pwp+NumC3fysHVXu3XxQSjjLrOTmiB7OxIBWi6gdGwiwCuzk+9NZw7jv+RSAm6sgvzVj
fJoO+F+hpJ7NW4eGjVivl6tsD3AHOJhVsbF4GZIqp3biQireNa8iWSRUSrg9dm4sYRj5vjz6Cixx
n5GBO0fcHlAKjDtOYxXnonTT8HDty8LUcYxT2u4epWugwRljawr77czsCm+3UkFZnXwhmciu2Tvd
wL+Oa9ksDQFbg4WKVegE25Cmjfe77O4xh/JOpcAqP0QVDUb1/lIcziw2077xf2jA1zsUSy2efg4l
ExQ4t4t1TdUZ7oRzY12vZpp1uASynM1qw38AP6czv0l7BCPcm8cZRupBLOqmbUqqkGFEAY1b9aXg
5p1QQde6J50TKAi31wedR4vDuKbjFw9Q7cuQfnsNHdeYvYoKXAPL8cln+WUjzl/+I87dCjZaxb7S
Z4ImQNpYyDpFVWSC7eR0wsvaaISsMv85x1Xp2yTtNagyfL9VXYzYM5L/9E59mjr5VaVIvufmY7Si
gtfjhlylEhbeiqSieFZ5R3//JK8rTp2sc5IplrA69Dy/0GkYMWZlewUyLSkB8U89xEWk1M6WFlj8
taayH2xqRyH3Pppxpc9Gr70oF23DSwalNatpO4OMbBAFo0wcD8hjWOsBrz/0T+5X6002w1nAouw3
SZf+NmS9O/ydIcADzW398uJhQ/HahEj4pSHI4xfwc/qRcAfS6rDYc7JOWDONjUIU6ZmzODwlKqtT
oA7uULfP/Gx1EwPKAK+7D/4p7s1rmobJ4AbXxji9Mj7ZCrju99eItHWMKDzr3rJmJm5Y/y4EOpBU
4iwYmS2wFflN+0M+d9W9VXkLOEW3O3fyuBwRQdhpL8TbWobSNZmJIbvAi6DH2T1ImtG+eZTS7t3Z
VSnf/h2PDUnGMjWf/S7ycsy3M2VxxwHaj0jBFPXM7gBCB/HY4P3SFC/tUtjnNvc/5DRXd7oOwWWY
vRusDx6en3rnaYVjr3jOis1+2oQ/P2rCsjPXADqJmnNrgHDvQq/J4L+9FSVmoR1Z6uAO1YEpMq1K
k0zm2iD67KINCD6rrKDer3Zg1vqEZP6XLu+1BtvWHeu+rSTc335R1d7VkLRGiN+PS3+r5CYP5PsK
sElPrmoyzt0iJSaxajDXhCuQffq6c3MegVwuCyqz7TU+kmsF/ie6cTx3CgnSF4P0ff43y8V6V4KF
anNiw6Of+s6B1C9JGoljm5Z6IW6FI10TkRJ9nwR1MJZJG9oFeP8bFBPxzHm61/XtJPABUU2w7Hjx
s6pT+pDf+6HhWp2tEJtB5pcam9T3UShOF2BbRaVQf2ZWW/usUdCoW8/A10g2y/JgIWUDdpjc9gMP
XJiCCSbEQIx43zNthsamapiWnot08Y4LvbniJ4rF7KJOtqaIPpxgtU4oZ/rPo9jIvbQfTbt2jFAK
oI2ogVCCMJRGGhR3RKc/f/VWbBPK68hBQTBB9+hieWsnRPYMDU++ldGpQl48Jghglwkpcs85Lvt5
gecObjvLYOXNJwT4/OulAr30Sd3PVTKOGLYngk5SbcnVJeQgS98yYNjDBrbVhzAXSmD4yYElxMLI
M03haHWdJVdqV6hR21lTudHXma/ltD86n4YsMEvjAuypJssOo7jHddH8HKzsV3F+f65vonkJWDqN
aqZ2zVTSkqTNJ+pJRT+Oq3SIjPh729YVjrCSrFJAAnYz7/p/yZkqhFzNFrWzBT9sjwKqXUHpG1ll
KRvl4yRABbVAtcq0aWtDIRLbBCan4B1jbe+PTsNsJiCRhfNIWlMd8Hsl14hMuFeYCsErvKJM9dkW
p29rrdFjj2GmCGSacvMxLccxoM4ITeTxErvD1IQqYp+Wwo6HuCBDBwQOU6WMNTtpLAq2y+ule3u9
j7sOLWrnkUYskoiUuWXnSHzqP5OhSrR1MbtheDk3AYUQER/s8WQ+R5ZQd6AQ9AhIN7za3a0Ecdhq
BikQB5jwgcpbb7qqK40g08ch7g9n8yE23Pxe02GDflcapx+a8gl6VhYBiYjyU4BltwJ4g2KFJn46
SgR52SXaozLQcXYQ1MYO5NEnjjBsRRoIg6j6W7Ewi5n/GuuxkDvIF83j7FpZP4JJoVzh2U2+ti9L
Y/3hmW979V3i+jgKBdJAv1DRN+EaulvDxnamTFS6AjAfLehpoOBZPxoi4znXNRU29BaRgz8qWRI9
mDSNJD/3aFxjAmx+ae2dcdlCxiDC5cda6bpwfjid7at9wYtzTD07hVzbn9vbu6LCixbtBVdNHE7i
XtM+zlJ7kQP+0fmtsHIyMEpS5u90a7ox32WiWOG/cmYdTDQIVm/8Tgf9NM+gIMyBpJ+S1uC/pV8L
MHXqgVQJSNZMFvnMv/EwnGMUgId7zr84dMsEfxICduwl9zI01G320yznxAsXh6cSEx0Te5ywK22t
QI/EFgRuoN6D4V1lgOMZ2avIs3CJQBsPaIk2oFAk9sOpmJfTBlKlByAa2UdnBQzS4Q+NAGOFjGkR
V3hMdmIBagy8T34hyRqleoAr1JxTEv9BDr35bTdwYcvTobcCPRmdfjn3PVKhsG4LcRXlZrZxo3e+
Vo4pqKQnCWhQLrXwxaKGPgDLdLclOgN9dbJFkri3zyvBm4o1EUbHtP4vq/AY2dKb5xY0lTzvqiCx
4WGAFQJd3AkhFNbhc+QzvJxYzPwRFCH50dvKIYdlARFdxix5NsT24L65gYipwuBOALeHYEOlZIV8
DHgoqz6lL7lI6fLQmthGtfIma0v5TOlnKkVTqf3rDupmpYWgH7iZaqJgAB55vu/nB7zUyxafL2sp
yu+0shZC7suoL6CeuH0Lc7AI17J+vU5PkpLs8N/n+0zmSFta+4QCRhVtz0O67sU0YSXq5PbB8YyC
rL8DWMFhxkWKicIlLOiREDqO89JKJgr86P0MJx24131yiL54em7PaBYmnSN1kQ+WROkFvmsoF8me
uDrp4Em0GOzhZ2WU+IsVYPV2QLaFW7eh+J7/lIuNDIKn1iXXIXfoyvImklIiiCLjcQQhUSFHh8g8
XD4QF+/+aGa8ofcDmpX313ZVObo8msuVTiupWlE2YVjqf+NuQRWx9vpjBkGmEfwBVB9jMu/lqcR1
eif9kQYo9pvYJTqsW/C5hz5mjEJ6aHQ7yechVdq4gtvzU4wR13PMmFgnQ+rbyMM1KIXQzWZprPZX
3cLtac66tjGXAa/GhPDyj1XLoW6QbbVlANjZ/doP9gIiV4alB4SjSDWqFXA/gKAHx0vB02Ylr8md
oF3/gsJD3Ncrr1cZ2T4jVVMGPqKzrq50XTft9pY1cPhHWvYdc7OgiDZo1mCfTK8QSpcCcDptHR0Y
lr92RvwP9L637bAfGJJsGriQbjEuzsvAER0YxcTMg7vUFnSvL/hkjzNX2PH9UEwJg6GuWCx97npE
bOMeAfgeMLljBQCmXouzflmv9IGzHSspKNIRludmrqikiCD+qEvy3Qq7wSNWw5yPzBnFG1B7PRoU
NwM2Qrpvj9H45mEqXi5SYjvVdwuqrnkUboiMKrs3JuXyFVQVzOO5j+xgTdoPsrF4tLlIjsGjka94
OSTUfA5P77s8ba4Y1CSbsF69SQoGZn+vQJTv+hyzHWvKktu35NYDCItb97cgvNEDzVgjVNudImzd
fK4ZF37y7dT4MWGpnPgA5FaRvegmn4Xi4n0f2ARwF/Vwqpqu7LADbE9JEf+1ETyC+QiXt+s4D5ir
7FgGPnPvbjhRIWJEJzAGJaLvpFfe9QXJdnkUpGfn2ilGt3LpTCN2DAoCHPZKQuoownYIIQLJwHUs
Lq73hswD8Ub49I3nv/hQ0Y3mcYMfqeHhHdQe9/knNzu+8LrKiVkCl/tfI5BNFVKXGnWR2l6xTJwu
slAoIiAaoQh5IWu0RMUDb+FHpETgf5YWxRE2nbK25H/50O/QdFzLQhITG6Az620GnT9pPXIm7B9O
Cipr+HNRluF6kiX6xxHLSe/+NYR28uivaYRhbG2ELOkGRp2Ll3lCWqEQ6EsZxefeFc+wneJxB0dP
Ml+a6E/Okgpl8tPE/2f1csFYyAKXyXuXfgmOxfK4kAudBKp7yV/Q3bXuxduU2wvCNoi+uracxgVc
WriZM+uq/oe/42OqHbK7uHrdeDns1iK+stv8Fn9Wkv2cI364ynTJ8G0O1orvIp+OdA5uQgX6MlVf
SuvQ64XnW0s77eJf65RbcqSzBRAksm4hEA1p+CSmYsFKIS9jwyyp9Ng3xmDL+Mj0E6Si5en2ZtQg
WFjH0lgVtXEqUQ3oE3kSOBgBzOpE94G/Sha554Utpn4y4CO/eFhWtOxcd0c2jfVE+s8aN29Kjb9A
EbQvGLV6b3htGH7vWfExsitZuBCaAShHIdmPpChF9J5rHl9O70jbf//BrqTVMxKIorSYE3tLXCVC
/fD8aP4tENxz9a4OJH6W1omVvPDpHBlRL3fn5OlX69nDuneFViERt1ViUyThf2evYXpni3BvoF5/
pDB/kQOncze9uAH8/WowPve4GlSmjjTcPtMm1M0WOzqZdA+cMksuA0EJ+ybQQTLvCJOdNs+if+gy
/dAZaOLNrr5WFSRG6huA+HknRLA1MPPyxuwW5KIwGcKtAEhoOHfANuJpSeyag0reuGZP2sUUIC5j
82oGbJiP3CwtglVHA2GYHJvUUPwi1Ou/Q3Q/E2rYKkTaK7C5SDkEhfDGV2XnqPxEiuTwiXUHNZNI
fip/lYgpkAHXBx3kSiJd7KS+XbMDXxc+V87ISDcn/GPIftCxrjfzapTO0VgJ/Vk3j+ulHFnsMBqR
iIfgCoVs7H4SPRU15rfLKg9lGgJ05s1J6D18xXLqFNpm3HwXcr/vb7uqpjrFABytGZ+0GQAUwVCH
bJTavCFQSjR8+2SRuKvutEf3/uIei+9bopGYEB9mNyesMI3zkGZoYtcZ/QKTV8bq//1L8iXWv75R
/KTjAIDXeYaYzOsCUQIrdgHo8a79J9LaW5FoImWhFyE71S+Ius899E8n+lFQNGFTz2SAooOh3GPj
WgFPc9L2Ct+GZxO3TlkVBYcuu8o2pgvKeLLAIlgqn2zLqpkoC98zo0fxVSTfGdbhxIqppf1yZiST
1/ukOkJJyOAqkkdbxok0SvdryvmChBhOXgHdzNw13aF2QATbn4BgZ20R2iUCqMRhWM9uq/C29VnP
lyr/be8joWv1f/p7GZvaIMJwT26AO1yqrztudhWMYRVsrmejUFoh93eHcZRd/i7OLVMuWGzHmb71
cWuScJq2zR1AHmiXJj+7CsOnT4lDSNWBXJ4rYS8FzNbPm/w9YsSQ6aEX29cCf5loMgzV9yH4jt5/
mzteFxRW8sZPNIH5kFHjKuvfMgnWKbgRK7+SLb2a98mqm4TrbxWg/dVREsblK8RuJveGEHN7YSbc
oGlhIpd4+QRxQszfyZlinwl3e8raezm+YRRAr8pqmh5zFTaNuHzo/0ZRz5POvGJsbyXTtwcK5yPo
GCRQvAc6ctuk3b3AAUeEQuaDQIqwm7oJEGbrr+OiSNmmq5rOasn97TYPYr8A8mkGZ54b3hVVYLDr
S6RDWusJoGL1Rf5hvrgiK7Nk2LoKEo1QF1SwMSb/AYd1en6daI3iBmztd545yk+KZMPPi//zqzfA
tYkqxnY+dM3918htCcvzIYja5WaRhqWpjphFAtFJoW4tsxp2yLD947GaMWCPiddLabetzFe+W68J
SKVda3YqyglSuGPFPffiqs9VngUeTv7W7zMK9Ad3pNxF5OAUXid9cQA8AtppZEputjkdOV4d0GU5
BjghLKaN5c1Kp8y++RYZ6ADnG/w0bAThEp4/pMHpDYECgkNfDJK1SFAqFkOu3zvVvKacqPirGfsf
1llrx0i5qs+bZ7RCgY0TgH5OuVv1ED1fZj2jsB8xT5iKI8GfG3HV0D8RibXcy/yCHZRZhiQNjeaI
SdQzVqh5u1SXeDHreNBPM+PCLXb4eJ1UoMqX8ZuvmUVJznhoG3AeraRWUk+22EO0cOkbtZyT7yRC
jz+IpT9xtydQXGj4/TrI9CcYdVAP/i9TfzxbK3qMSJ4QGDYj17Bjn7P8r1lvP4N83/YbBie/NG0n
Jz9nuPt0zmUiyaRi04ss9B/BwUH8xIjl4JG1I9kap7NUEnmL4cHO5hQo5zRWTdwmyPcjZhiJqGHc
OYt5tepmkU4B4bgAbylHs6zESV7yByG5vaWRiF03il8z83ifywEYGpsnHl9hg10fw/hChYCmyrGu
DvpTGI8DFqmJpqJ9kBzXPRogldZD8XZgvBu5NSZd2pwTHCMdT8i7rEnb/1QKhaGzlcZv6vEk9S0+
tbq8HETnBT8rShfNBcrkvPyS+euaE5fzUeBB0rj/bAv1LjE8H++up0If3tJcWet/tRdCGRiyRCCk
EHTXDalKPRrG51wdf8NQpSGCe1zfKgEd+stz/KLMOnKyr85aatcoSzY9PQttcXSCPfxMK/30/Hsy
D/Yq9CI4oEWTdJ6tFSiB+2Vt9HRl/0g64z7C3+9NZYA1J5u4RpYFabeYNhqeKlNnCyLlJNA0dhV4
F92aOFlwv/suB7fcddIhquYKUmKELXfRtiDu3NOieXqFQZexMi+ztjhqZk+Ea3NBoYFSmX9Esi8K
HenskxpE8CHSdbFwc6W+g6guYyLmJjlWicZkpkgy5p1+V803eM2BubShrwS8j4yYI+jLaAPcnYmV
lKTne6OEvg6492C8zl09prqdw09juJ6yd7YcwlowaJiv/yvKI2s2UIYOYOesQocdc7bbIfWiEqW8
lZP5+VgFcRhhGqV1SBVtuSR24MgWE+KIq2SYyhAqCA00y0kHFf5SZmR98rwQe6E5RTQQwn/WwYDa
3R1Xkmjp0lk1qNm0j4GHFQB0R3O/YSUg+BEBP0LDKy/pc8El31yBF+klODugBiuS+WdenzZlRfyl
ZZXuxIPTF35nipdOdQ44M+xN/xgJ0wwsVFRIBPqVKXFCXt9SGTcYvYNaHwXCnlC7Xbqb7e92Yt3s
KNYCFCTGs3u9lw+ROlHL5wf0Wi78zFRDy2IinRnevrHoLTotCcZtVVya3H6AknESKddAzC/+HM5r
eNRE2nmQHoqK/h8XPshz8Hp2vJKLoZin4I5hnGDL20sbkFgvVrIIRO5XSmYo0P194c6qHVMdMYTq
RYSnJnHvHDOY7INNQs61TLBLIkug0uSgHxmfBZV2+EIbFF1tqJiLmlJg0S4Oam1AVLLYVv/vpMMd
rj+VAoe1CKiPI9CaaVbQtQy4yUOJQlAxMy8Av41g3ivJHd6v/Xegc8YdwRlcpOtaTMGEhuh7vbq0
5vW/B3dW2d8GrNIyvtUgtTzktyTDbfWDUMov+JBDqVnMb3eIt35SAeIRGiSGmxa8QrxhkiyGXQeB
QrKUs8T6zNOPBrT87T14NAGbb+idUSIRBjono9z0uJxiQHmouKWiEKFPfAaxnykSM5Jefdu+Ta01
dO3yd0n7y+kcyVReJKGN0iOxmL9RlB5a5E30mYWbuYVE8kQ64gddPwQJPLs3xG1cc6LyyvAy+m3z
ClrPKF3RDUAA9FmGdlHfcUITrIC9bT6NVp+/C6hmbqru3v+a2CpjQM4yvp9maImxGJHkFFTFPda8
PRVyNoDLXBjavVKpB5RJ+sxMxD6b/2d9FC65VaHFrsMdKbtsl6BOaIHBOMMwyk5Dc4QtjdUCddVo
UVo4tXfD4cKyJaIA3f8PtBBLZFsgimhvF+9JcTZl3BWmSszmA0+eRaZvIfgnUs9z3xaIymsbsGYd
QtkmcuayV27zuVzBaqFVSHfwJWTK99E/xCoywQh//ze0L/X+YQ3o6nQnuQy9aXk/dT83ybfQjYHV
BdH8ZZZr9LIfmNw+jFwP/a92P/X2gDvYcQVAKblRa1v6xMqdK0UeBaF66p7R0kl6bleuagQB15ij
7nbBgpFcCIgZeF5TBJ+zHaDblDsXVYnEUD5KsojXqgQT1HLbNnfm3SMUOQ9rzZ15M8Ve9GEYz1wE
gDWZsTlx4EQtMX+kFUft30aIQYuyAa/V3HIGd5n6tpW8wiqCvSHcSJ9MbyYnxDajU9glCS2Zsp0L
2asuGqwuYnYlqMsy8dXlC8TYwBZfHkVlSXVp7+GuvrMPotVRxUMKzedGznRCmKwcL2QH7q1gfTlk
C8mBrBSL76ioQ2FTlUcqktcPEVeakp8QyLr+tzcltLmTLu5uKl5lr2awFquYrJpYIkBJ4YbjiSHR
TBsoXdDtS6xT01RdrzC5ZK79CpGo/qA1GwbGhAsUv84QzGoLIcUjNZq0GpELT6YSCJoJX+oeLVRI
YmtQKLtqoeXgtqNTDKYM/j9A8Jc0jDgl2iPV+ryeNsV4vUIhHf6c5LVtq+kGG9W+piZO+c9UseOS
x+AqTx3+Q0hgaKcr533dl87OAzgRqxSFq7u2xxNKzZSOG+9H5E1LhphWi0otCMKRry07Uu/pXNC+
5eajXfiqU2yUIGCGSNjd7D/GwzbXOCNAS3HSX450csEiRjmT0CGVssMytgHmH/6RvTF00EvJR9hm
HSb3pX4E7YJ4t5wUeuUE5jUe/5d9YChdDH4zuAWKtOFTCnFAZlMF7MkqKb0WUnSg6lJQTFoQ1e2O
ryfIvIWI+fmV910M4tlvQT4bYjjeUEAeOJ4wvJHVxByloT0iLlXvSDh6BUVVeN6CVjL02tlL3uwa
q/4kPhdkfMeGpvNxMriwM7K8rVqP+VUJs2zZclW2t2IauDSgtCJfmPCZzfv0ynrxH3FxcEQUsbKg
6NguJQylJA8g0u1zykg693CF7hBJ6slHaqf/0Dkb9kHNmdjdXYlUgOD3jego/f1EppREVCGz4Vt2
dWNoistfXALcr76fH0bb3pVziWHXH+VlRwGS7YctzIfZ4UQXJl9pF/kcI8PzER5qq8G7tJudp8ei
DqnKJopKx6ORg6teLI6OK6SZCa+M+QhqFX/tcBcBMS2gVkmoHQhwzehYhXdT/oBjzQVOjrHQvIaS
l5awnrYE8Gtm7d9PZ3r5Ea6wRmfEc5IHcb6h94yB2XFd7nCC5xldkzE0fPqBi/T0FybsJGLGBb1O
4AUcMxv8tBatF6BHgpal6DCwdHzbT7PZXAEaDIiyA5ggQhaQXsEz8chldmbL0xk1jAqabun8SMTn
CTk6XBH32LBtzb+vDu9oVKQXa4Oi6kvqUwuxOK750yg4/qUZxrTVgUF8qVt3GGxq4Ko/ipCMfRVY
MgQa4zLwdFddr+KfEqOGA+PqJbhi3OlBx0CVLRsryACAwrLpDjlY/CsqPHvTc0FZm18cvUhbFctq
IeH2kBtZgVPF3jmEPyEMKNA6A0nV8EncyTHBscrKD177u0o7hewGbYH9CCN0f4axabaqcZmCq2vT
dFoiMvGmvFnsPGoeO22/w0Z/uRNIqADrwQDKsnJU74mNeI1NXe76pxQlKF5IBplvixyJ4O1n279I
grjXcPVejVQwgxWoZ6DIou5CAPIJFGCZrJbuqWN0EUCfyKKcYNnJc/Ai2JHtht8vg0L5CmDO4rR8
+EpCywbrqtvh7pIhyWuJC8Ylu4MMCMjjh0Fh/n2g2zYpG+CTcPevIgB9DQOzwrSMHpNjtg/+Ut3x
VTFT3sWqjevTY0mrZQqHX/WCm9vJ0E/LcXjoNz8jXrU6xJVP84z67vE+s/jU2gn088ME44ElYtud
vHxUnSK/mmCUwftUdSvcKj08O7EE4RazFO7YkZnpfYgeQNArUYHMJgT2mJfFNwqNCjUPzLpFlmzM
Hz8qRwf7W1PUYayJE764ulRRRLT48q14VuYJf4cT4bAHy1/l60NXdb2egFuMqUKOEvJF2ykiVTdl
ZvPSSTn84iMoEUNaFzAsO6LM8afeqS6rhV9VTvYO9Igvy/RbJZVANNxQL+Az0x6jaNMB4J+VO9fg
aiIeVZ2unM8dW7UvH4lMVxPN5YLznLMwMxEUSOMmAO/aFiGi1LUtA915jqOSdgDR2AagCjk01tqJ
UkN9lECPQwLEFK6m4QL963IzCdApM2NwIb0jcWn3NoE95emSGiegCTqmi/+hYwadxKos8gyMMePE
vCxtwDz9s6SHY06TQL//f3VKle9wamSvjqMK6dm4UCUQoCLImRMRgSZi0NS6WSji52mToZ02+9Xl
B/QTEk0ZYT0vPlc7Ykwk1cQ8HolMDe0N649tCLIhD28Lcerm1xqej7HcFTfuDemAr2K2znGxUs0/
HuV/c8nwxfDb7lF/pV2/5scS4m3iKUySnb0gPDtZNHXgFOn90aoRA+ASj4w+N67rz1kJ98Klof12
W7yVfnoVUWlDfAldfg4mottsQ3dV7eANsNaqWCENTsUri8TvvD/7gPWftx4cxgYseetoHUNSA92t
hyI6kPzk8vDsFG69+eHcc76YZscLqjXkeOo9Kn39DpcX7yedTvXr4dDU90ALjG6u/pOXy1/B3zA9
koPnVJMHxQFXTw0BvZ9HBtc0OJeomOdw96F+ze3w4Aw6xmWb47MWCjAeIkeGArEdf8/wt+l+WCH5
FE6toj++YheD6wHl+9Q6b5JKlvGPbSeiLQLnr3mf5gIInZ/ErLa5OUfBBjKtuIfvOt92IxUsKaqj
IO3XqLBjLlkaS7fCxmsluTXmkllOwRoKqqDaJeAnunw3FyqBqL7yiZy3RkxrxivuTfOsXALjowKE
R6GKp1hmYqJjK7gjMXvtX2k22YryJq2zPfVSRhZBoXHJaLsp5zn/sNrChxJrMrCs8cE9Ls38Q3MT
+EqPfudVoQRzmSVUKxUOOtYJKv2B0IEhf2hDuBEBPIg2AwnqDdwNG6Tz4f6CAuwIfIzrKdV0j+lj
MN22RXxviQsoc98piljbBDkOSr2pGWB1vG7sZSP/Jyv68JnZ4e+T0/LD/GLWON1La+Kp/Enl/yOP
P11+Zry5Hio87MZS+Gstnpn5DuLxkBtijY4fPQXjgtLMnwK3gnxZxCmmvDECTZsh2+YVbPps6GyH
LpEWbMgQ1LDXNBl0XdbLjkhaH+M+jETiIWNn6STtNg0+ZosywXx/ygzvRkmYISG1B9Pss4cCUtrk
ZPyEnHvxWPOfeNs4T4zQBZ3U6OvlY3of9oeMkj1gPWAl+O3UdC+2q0DxN4Sm1nXTsryqtd9IfnzJ
HRd/O3RcIryvGTUZPfqZKCfmPqWR1sKbE/y14tQATJY0TkvV70GW6wE+U3qWV4xizU/AWyfrAO/H
lRsewdVJkEGjJWyngdpgV0mJAH+LKgxybZ6Kp5kFEMdN29RSYjlaYLsSYQp0fappJmUzPIw2tMgf
+QLbPlq9XyQqkKL54T+zM9ylQSzO7sK4O5g9mkj7mg9JTdMd1Yu0BAulgVG1MvWP4HOvob4THs4Y
EoBqF7vFlZQ/efilufCFMD/9V7RkCDqtdegV1uPpFHKuyoZeMUYws3Ax1mF86kuJJ6zmQWCW3mZM
MEIRdGnJOFiQgHG5PFeUwdue5QyKrjXn5vrcVulNbt8y8841gvF26/Hc4J7KoFkbZfL9plB0AvMd
CO3mUQOb8eK7RVEJEziZcxtg7b2lMhLNuZSGm8sZQQhXecW35fPGh+NC7Dn/v7GdreaStJP+D0ny
RROR6v7A+hGsa08HZOgm4WGxRdtxmXIIqGcnVi13NwfIuNMff1xjrJaftXwZG1vqojTkOdO+d6RL
Wvarh6FPnd3VF5bwhsJKQYirUPxIrnK5sviNNlZVuu6Unq4wfYwYrfbfyu9vSqqvgxBxw3rFu6HG
qcLVttTNbYj5coa50gvjxFsNO8aWKreJ1/YqBLAN3RcF60hUR2UE7VfN6FyQCDHAAAx8aOhMcMP8
WXRdYrejCQO7/DpAJr1kRWWHHgIiigh0ZzDf5XYmYujalX+BEV82tN/HAiZ3F76AhF6gAMDRYEev
r5GdwjPrxo0AQys1ThtzBm/gt1Ct70Myw1TyfdCfw7L09asIjTVy1+IKuX04oRsnRMOeTXyREuCD
LSzvs82C7wX2vAv0iR6CQ3stJtgh6oTCKR509urGxI+yHvV9ikN00EEH0xzpBTF+bnH1GkS7Wa2B
JhiXHQAeLRkhTQjkZx31stpyQ/zmoHYWmU/88uNCUvBBFDWVbn4p2HCpAbcSbvxFa5waeiZq2qWh
OKPokD4xAFGD6EMgBLRPCf9GIuMS0IR7oex11JEsfgtJXGhO9vTQPO34Klsg0hEqLngefCq9Wcpz
Lnp4298ItKFldMIIaDPdGerOeDA46jXa5fIXuaMe2iqXbzIKkKG95F5WV7+Zu8wVmm6asb/arC9J
sSiA333L7kRuUWfzj501jld9auraQyXH1SseEEjXbK2WKgk7oSw2nyDNHqdK+JKH96URA/LFpqZy
VRA3f7n7lM2ICVmSioEOuXVGoWAgbgKP/59IA85u15JRK9jMSpnixiDPTMGxQ/p1LD+nKULcqDVP
on95YyE5BqVs2yUq9mSjlzcoJ1IUc2ATevfUBo7P9pbaPWhFrxjwZr5AcgDfHlnqzkaeJjAhgWfB
9nIDNrzdqFRjSAVwZ0x9Y64X8wu2Pvauy2JBHjIPr/1LlB0+X+E534L9uUQabpI4YdPeUs8W9/qU
8lrYel+I/IA3fU5ZxMOaisOq1aRcoaOJ/4QAH0Kcv4OkhoOR3bzVyeRDr6IfJa5XvWLnI3MylKs3
s1MuHv0LZqwBcZCAc+11UCeCWlgnY9ffHbsx1rq9ASMkkB+sg99zoOuPtgviE7bNiMob/vrVIvkW
xq2wjh4pEl9aFGh5N+7+0f0CFgEi9mX1c+BcnXw1VRD7kp5zh5Z0fo4sCrW4tkhrfSm1XHgaJydU
38xcihd0pbHJzz27n3mH5dIk5mWojtibD+Zu5Svh1UiwUL3sVRDpCx+S1/mgMyZyX5K6cKPieNYx
liCzIHjDnpDRa6xmx0raohUZLZT0rcXuGBLRdEiwR/4riU/k+mrdz/pyol10wSZYvHee+MDuKuWz
YDDSuWY49YGqTnNABW7aXb7M6j367rUG9QJfPpwwEqBIj0fRZb/p5MTbla3JcIQnd8i8osPBO8Yj
OGivFzDafFrbC8iIfLjOFDpZLo7ALWQZj5r4MZF678MZJgH+dpegfAi18yx9abap4apbC36JoFYU
k6IGdp4iycvd3CkhpgnIlMQ1SkULfTld6MA3jnzq1RwBBtroi/TqrQ4N1/twUgW/sL/nVqe7Sj7G
vCEwJ/Pi8IYhQREGh/T1w0Uw7m1OBeZ+kgAhbtPQsuQt/89Y54UXDKxF3ma27m7U7HX5d8UWGVSt
Tby8qL7iDry1QTth7f3R+shruzu7zpLihGsT+cSXJuS7f1NuEbZGCmvyo11dgDPkAYXlrLwpPdte
sgfbLAAD8vrcxvZAl1FOxC4LVsc9lskFx+fE1hgtwPZJDvXkNHYE9/bk49B73k50SO7EYsTXy8zY
qecgBFzFFDX70Y0FnDUGWonBhX/hSTilqfN3hznUnGUmf3t0Z3U1wV5w5cXqde8IgcA/e3ktBUoI
pLInANp53+c+AkU+bsAQ1FMm61MmaJyJfca5WU6PIJKpjYypdZEVXpd8cMPqgH5dRtTMlXTA/NtD
TX/BbnHdVDGRXi/ENolLyCPAfxLFhsu6itGLT8Q7ZDCHYm+TGQO2IyRjOKD9XVnCQ47UnY9OIZrj
YzqIWTUiT2Obvh8mUqPauy2V84TBwQR4sb6R2igwlHZhfQw9MY1RaOWB3aRgLoRK+gPWLsNlW6xB
ALvdKUXwanqvl7Ux6TFXJ0009xnhgh5GyUgxzNBFe60BXRlOqFCrO6f8vO0mTK9cuYD/N44IVyfm
Lp4ZsQfML+tDsxyJ5aFjKmWCloizaxcjGQLbIaQLgeBdhOQ2hlRxSpgEPfaySoekfGcfGhHtwQ7M
dzxOt5OgPWgZr7sl1ELZ+F6YgIMPuX6qL5sUfooQZQsT1KpCh+AjuDfh4ZSqNFS2b24wP1E9cgIm
dqQgMCjslYFhxpU5BnAHzVID++12lmb+afvfiADURjTwQQ1FspdaJ/jBtUGFOmyUiN3jMYT+geU9
l11zAqAcsRgivQIe4tyfWuZV+HaXBiQb1UAuGm3Tr8X4HJiWsdlT9fzPUnrHW960D+Q8irC1j5qe
RRXXxZGjDT0ZQX2UaocsqXFs/oo01lPnQnT2yoh/N7C2LBjP7ARcHYEaktSXLbhaQQN18gBRMtDv
NI+IitnywWJuJWkm8AxvCaaxK/TNpXjRW0rlr5m7Asr8zdSntF0AXf8ZuxfvZvhD+AmveZsO9Rzm
SFM2RCHLVYs/ISTfjjZN8vm+nktCXEu1CyMTUKUGGpnofOghpMHvcFxvYe75G9zjNyxpxbUeVl2d
wHpAYM74w0sa8lMqxnGJEy2WsgjGwkXGWwezyruUTJQ+zOW1ln/hJ+VX+oFIXavylhnIJ18KPzFB
KWJAtDHNeYlfswEDhGufnbBe3eIUkGzIq0RsxFVJFai0O+muI0S1Px9twKR9UCZIo7D9dmO0Ieb3
YNiQvo24B/u89csA15APvlYU1cjHiNra74ZcEEzLAEwpX/buUzBkrsPua5AcHc+gFZsJ7Ta+hl61
XacXki87KrfkCg+BUhnuevITa0cb73IMm/zl4p3Ok0oxVazDeosE02sC1vzy6Nvqb7cBUKGSzZuT
KXIKt5L1zDjl6EJSgJ0HAPrDvl8E5RncNSTZX1c1Xhq7NduRuod5FFfA2nelpTvrvVwCZI7i023U
XahDn3ffSc8qOUJKETk8AMmc43hkk2h+KO4FtM5FbMI3QXL6zCuyx3fiek09lH3KD0Ff+rDXkiqf
qS3MrhPqiluFX3l10zgsMcxrn74qcCTxqvJBLHEeEGhXcVXlRDbeLri7sRxqen0Dx2cZsyDaPCpS
PKXHCbOqCwBadprlSF+yH+uEW0Sg3Jy6ZqKCYZhPfs0NrYXC4YFXQQS9RcXX87tAkOP61TMAPYK5
KZI+Eu/U77QKdbAZxh0l8kw6ynlPLeDWEkO2xRIoFuquWkaDUxhRU1697Jc8TtJK0sE1ZGkEtEPL
EB0SPrbZCMERUPREyMfLiOO/JJUnG3v+ozytr/bMGAmgoylV4I4UoQUB4GBp7w0PT+LvxpXfeKSU
6eJy82S3Yh1NQbbFL4ewAOb+CLSmexzLylotTB9EylPnSpk8XLECmG1Jet+ALfYJWpuvVtn8J3Qv
X8m397nNOxTTgmybcHngSLFE4dHnvmRSJCjM2BlAW4Jwa59Kvlqg4UUGPoxFgxrgGfrlQ69H3sOj
unkey71NVT4uNN8VK/YjaNZx6ndR8x8MAnJFHbttUhvxdwSZWGjDAtkaMawWrJpvi7+Ud0hPpUIk
QMvnYVuUOptGn1w+aY7B7Dqi7gkzpL7CNHP+zU13YmCAGMCZSYnLjUj1UzfeRrQ5aYJ8f/xd43p5
8si4XsRa8Gh9X7U1lA8dOhVuZqsAsTuKKiXEYrLID9lIofsLMlEGSCH8afoEEVAZU/UVLF833ak2
ZNhlNTsVY5QGJ8co194nv14UqWpNFZ1KEP3l942HtwtsM5w0oazc4YUvxsOZ61cFYgjC2MKvfmvT
cxN7d22H+khiUbBu6UjB2bm8qvQOjx8L/GuD4ZEECoGOH8/QioVoIXCGJPkVkpEddvpW1GEMp0S0
P7kHqV5HGts6YzmZiShejOWFlhnfJAokNkiJGnWt+OIlJd3OYjdcWICKK+qPFVPrsYBQsY0GJ35W
S6VunlPr7fp6xsvvDOXgb+nx9tvGRKCTXtg7IivZJjNNWNUHtT5caCo7RdvbGc7leOKvZn2SlgtR
N/LvSWpOX9WZqir+8+fQxj2R3NRpOxJlnCT0szHvLcOhS1Bceo2OODSmUzdmM/f1WrTT/1rEbd+t
iCU6yZAOT53sVtjMG6+MQCDIYfvdqBCLgJ/j2HSpqAGrI5B0YfMxrK13UYpxX/cCTg0mzHpsFTUs
VIxvYL+AvBZY6Hi6WD5lb/vI9lWS+H6N+0qQaw6U+BOjeBdjbX5ZqFMCRu6tRuQTWKa/sjwc3z4/
OPk7gpFF7bP5whqOB0KjF40QiwvHES1wgfMqMhvgygKMyF5Hthtr5sEVrbJNbjY10UGyCvNYrPEq
DpwKb+C5ZWXUiCisVnXvkaN39GqLe2le998NI79eNXaPEAj6Ze3c2MojATz7tamJ0i+0Kvoybb5c
3tZMe+WTafTbPfwmol8y0J7JS3FMR5R2rvKT3twbVqxWUC2Mp4wrTye0rVTmuMuz50OGcz+360l7
b7sJyKt4G9d21gbhbAi97QIpUcg/RfA0q15fjF8dCAl4L9ZKuVBagSdQTQ1eWogGtxDHuqXES0Qg
OCuHA5bNbpfMvMhMoN9In8BVh+h1iJh0DUla3BZljiXX1DKQj3DDufCIyHc3GG9f4qKN2NytotbE
K6UtGXjmiHzd719KNmJNgXleiGlZDOWsDs0FISyJBe6/ZvbJWWbnuo4QlUbogHIYvNABKbQ53Lth
bEhP974a88wyao8OtJHLj/IrOS43YPfRmnC0GL5M0lI2bgCHqQJATJ0gqBCWgbCVTKp+D2g7L9Vf
SLT9ncEXnpMl2xjGLCA0+8poEPMPjjDhH4VSMieqmAGKUaO6pCOhoxm+I3AMX/RaFK4f0U0lsF9v
+ALtuMbuQWDhXmOuJw3SYu2NaYX9gF9Nk6lzVx0VRamohBY7MVrJslpeIuSaynbsAZW6iRHl97Pa
UtiNGRyqAPZLMLr1vnO8xQy2G/essaqn9UOFlS6kpT8Z8mDYISGt3C1cBjaQyDv7ltPj7gLAzG1g
sKWNIfABXGs5lVknqBaJ4VcRcls3wF/iQQNsofCummPCNTEy1hE6IIe6kRcb26mq+HwwmFqliZDq
vRChtnkhFr/2hnpfClhkicK5S894lyta2BTt3WwfBv1I3zmV8gkKgiky3oPBvevKuRrDfu0lftNH
NA0e3IiqLkBIN8yGXzgnDszYWa5u4x0Ppv7cRqyklv2NqY03SKGJ3hjxsJsRREfbJKnwquF92hET
T1liuieOtSas5YaSo05y4ZR3TOTKGQg98EGdaZo7RBGDxFwJx+7Y73KmOr547OqMZlEDvkXFVF/V
It/AkWt8g/eo1m9cgMEDp+or2e7TqZrlX7/KVPFhb3KbDWCsO5iOpUgf5paOg4Jbj+02WdzUIW/v
55DPVRwHUwMGzpsFlffEGDHGLrpCiU0+6Ip94+ls089qgSui2a4vFPAj6gt2Znq0ys9rC+JG/xMN
sppXS2WtmJDauSHY9J7yHgzxdoddY3bVXQ+RK/9s3eaOTmwLmCkZ52IaOJVlPSI1imfymLymWVYJ
WOHfIrJ8pdoQkNiarrbckBI+2Q7qmjdbKyuRoLuUPElFFzPhhyjTmbCf+AbF6nDEEdk/PuC6JfeE
QVp3YBwPM9lHOnj3QW5nlSYbS9XJ75HGF41bRr5I9EhszIu/0WcLpi/LWiMQWSfR7CZKYl9VC/WC
nqqZcb5vUnMF/p34x+LSv3Yp2eFG0MYzF9FygAHVYy46kx9vFjDmumbWQI9IOuetZR7uaVvPauzY
iF1Mq/sJjn+c73Z5LkZ3zClgSNWCf7WlAfjbK0jt/NmiEDs7znwXXc7a+Gl2PVwa5NjajThHK5CT
wNE6jHM9a68XXuDMIaIrMQqW/83Y69XXnSuk7FANAsraj+smtynJr56qUEdNJk4bP/ax0KGWtG73
4yOdGaJeOjFHbMea/QNjT/nKOcFpFLtpMFiGfpGXqWF8deoVR+60MslDKTR2Zt/lH8Do7lO9Rlu7
KCmMldolovUCzHLZPLm8F08EBwn5CL9Oy8YpVewDtXMjmGPGdlVKsUcYdxvAifkypKY3O9LdpmfP
NJ63QbbO4swphxND/LQ71wuA75TEPjD+mr+d77KfpJmuJpUSot8ULZXifWKx2ZhF8r09Thn/oNVY
9r9OOSk9DZ65mX+/OWDknUcjmnr/qa3b8fSJuUdKL7dGtJfC7tRZqajY/+fB3ETX092SAgo6+JOl
ZoD8CzZU6OINBOz7AUqgQG8XqFtmHnkTV73KAJlNCX/tc2tMmfPSH4rEcXa7ApGhyYoUwNxZ6yw6
0g8bbLca16rftaB/wh4D4VtwFxAKPjMSp/G+K/0hF0cIdLXq8ikB9OgWlVjK5aei2V71OIDJJ+aU
w8iqaiB2BW64gmpQz/CjCpzWd1tRyJiBBo5Md95WKGwLhnzgEOyVurLRJ5NiY0fp2UkFCKp1bLVy
QVf0krI5kG4dYC7MW1cYo961w2wChMG4JS3nBxeSAejpRQerOOqfBVBd3SZftPtOCGlGijRzgf1a
JgTQdD20/AzGkMRbZ195oOYwzWG3ofsChCbEgzTTbhNjGjf/FCcd4ZmVs1BPG3UfwqiVj2Z5A9m5
mEy9v30odxzb0xSQdsEnrYtcgBE9EEQRr5SKy3VOvtKhbUqjKF5GMT5iAhjbdzE2NebIonWoNXGs
3H24vIInY7G3cg5GQhY7zotqZDMt/erHEFmWONFhZExD3NDzvPDWJMN5gwKawqX+Vt2UWpNMcV2T
5ZmNKRnkzD4vyCbJNNnQk6kEAZoBBJZyGvD9KrOrxV7uNfPzkYf5QIwST6C1gxjCZSajJOvUCVTZ
e+yUt0B6EBhLDgXqRuNJP7NU43D9RhpURQQXiLHoupj71EiXBwpjPoCYCT0X8Xnqqwy/UoTVjvbp
d3QFnLzU512IOhR63XAtxVFX56DzhKd50O0MdMjQ85iwGJecdzXfVzKxH38DDy+xxKIcadBZTsi9
rgjVaPPIWPUi773wpMK7cvoOqTunQcr5redWSi59Vpl4DRSSvy2I8g/SdRM5LuEGvjErkQGn0r9l
x6aJRgwla60MlLppo5PRjg1qmGb1PQUtFF45eEXoF0TM/bn0wWOMrneNjkXyoY0GU/vqk5hy5T3C
gyoM68cHqzJsDAuM/tAOpLSMIp/hwtiQ+rKJUBh54rh7MKS4YaMvZSN76/dJx6JJIFl28J1xLkRl
jaKOhN/DS107vU82nNfL8b6WINWMGQqyYI6BfhIVLPCNhk8T+oUGebfkPwoq0z2cfhiDZK+u9sft
rQ4B5bQbkMSKcw5i6xUqbCKPLskzpuWnxarAz9N7m71hhVfCenbTULUv8mp9qfDzPk7RR/BIIPKL
t/IX25kFP0AM/NgGO/Qw8eAW8xxnQwEP+NhtfkEoJr0Hn/DRxqeoBn8haWqDkkNMpig2CqITJclv
lr2G1DoY3EO3M2DjsORs6N73LPGD2dWjYXAeuCMKqzrausJDzuTmG+gBCwSY02q0J/DV4LaW2kNN
9YV1JuEv3F+nbnd6rd1GdFmMK+rDcU2nCUbBgR7U9QnWTeuRiyoHWw6ac6DpwBEOtpu5dYbCPV+h
a1+IA1EyvJ1og0DC5d7YBNMG6S36PmNIO/MFDfyJr7oKeOXEfBCf/40tabDTb823vVzijiPpKhOK
iLQjcLuG6gqmBO/t8GLt/WqDHfD+94Q2b/KitNShjjxb2vYPl5bjBOx9wtCL1rnNq11u/F2w+Ura
pyojqHXg00NMwEB4zUzQg0lKYsZSH3x7APUdl4Pe1zAfBbK7HGAlNUVuUYr+x2kY7PdY7y7b0aB0
m0TL+A3gJIJmfGjzJ8mnXaJsiWd4nrnGF+dVGiCfTpsMOg6aupa4rZG1nj9r7h9WhPy4B052V64l
Nws0Ql/lq2fZ1sKPMTT9seeuWQIA40uPne2pmLDHiCXA0iXhRpBhwb5DC+YOQyYQ1OCc/mrAHvYj
szHP2QgI8J7y3h4tFzH4cKkjzYthvoa6Uinpv5/D5xoWuXJ1jeQI0Top7bTS3RWNi7C/kNs1Pr77
4EjBh2dSF8GPKKbKXQ6t4AdNnqZvE4S9yDh2I3ZQ9knhMTcoCO2lWHOw4QKoER+SSf3JNlwjnpQ5
62/rdfMEJGpOYVtOxrgv4ePmNHwRxL0gfIixEuS1IrfAdh6fgYhhHIIYzRVJ35w0+wHWBkDsLOjJ
kCswLpdFR6biwfxtMlP2KHZLljRjq/HjUzy1jNCYyEEoT8OvXk9px0vQ9iZ0eChRoLmOZbgRkwqz
scxKoZ34EYKRtwLZIpKrTJEqFd3ODlMYEKf8ih6N9Rc2ORnaSw+OHp+mwU29+DxE80Izv33tdRhP
30J3vigjYpRqlPcsF5z7jlEatVsRq6sd5PxK/o/TpqftTDAsuQDDUv5j4kyk2r9JgLOYBS/yKxpG
49RPCDLH7AJpfKUrcVkNYWVhWKgIFP/WXQHpqhdK1q1VjMPxyv5d7GS6d5xUaWxmsKAJ0Mtzb0MI
bYjOHf3VyTe/Pm3CnkpypJguC/+iqBFcX3Y7aHuVfsUrLq39fv/YfRsSwu6RaITFX1h8C0w9ZZXx
Ylx4CYiPL4LDt8rz0jSDY3eh+DvABMQe2Aw/gFruaJUtHM4VYIxw4OWRpUHmSRIyXNadqQVLM0xF
y91iPqWXykgvjcnXaa85Jxq6IivqdVipCCvTLFIJfzBu4SFXNaXrbNIF3fN7h83ptMHDobJQQ8Mf
dQsyo8b05YubMWtKvVC8izt1FnkUza/PADK9NBtgK/00ZOCRxrdcZXr/HJ30trgqmknVXGa39P8K
t9CppB0VSno3bWazhMSEgm7+VyLQrD2+9/U82ICtpjue/U4R2prtj9lLPhA0DcmPvXjRnTWrgso5
ZigIdwAO93Srj3x1PETA1V3Qk210UFnu2RHjffJTT9DcL65zOoWouJSIdmUFNz0zFSKL303ps5Zh
rkZP11e3SAf8KnQOVETpqRAyVCo+d/u7cZSAewqgVo0d7Y6Jh6lZKOMldcJTaWBreXk1c/qAY1xx
8s/amG+N8QgPjTrffXuL3XdHZWuea0rfVUCSNTzXYzgLjlGfwN3t5Ks0Wmh9BiIBPh36WE4qqZ4m
1LSUuJYrJC3+tg0W5wbndoO64P6bWpEI9w7wD1w2VIi3wvqBu0TMRGCJhlfkXFc+WhEr/r0jEX9m
bocv5BUt/4CXgebQvRci8xQHJTKK3Ihio4q5ncL8c/cHhowD8v3pkiA7XR9L3IoGIBOmbmvom0RC
l44aCkWasX3p044Gb2bLpc6J7kKRhnM8HLFI9FHqgTUZTFGMl/1Byuvm77nHU5U2s9K8S4omzKvw
DToxF+yUckAS0JJINFKgZ8k03CHOWdbQ30k0Lyh+fMAqBzdrrOU3XH+/Y8rq3WVsY3XSspm2kv6l
9jd/5NkaHMja/BVn/CPY0qBHLGePnFcTzX/0ErwYCDrlMwTa0/2DcSujYvad6NNbu31RUpdB393/
FqydhCUa/NRHSgWOuidIuU67C+fh2kk4rco+qy87TnxY8dfNRE8oz4MvUR+cVgexnVtYX1SL6z5Z
Erkk2sInSJGVr+rAtyXq667H1jsYehLeFjYSok1EQAVf91seWr+DSKum6pbknCIkbbbA8Z8ZfMOK
WngauT1hzA/7X3pbpGS+I9Rsza6+6d93GN0krEI7sOsVZDuE6hHwlfE/XIHOBz5hBClYMwB/L4zs
jbUoo9E55BKRxwyEsgXhB9NzIlfGMx/NSZ09egplvr2ndxBdMIlv0P7Qt6C+ksPtTeo6R4ugTm3E
NfiZYc6mp+2pY7G8I2lM1CU5q818CUk0dZTge5MQC70GbPug5Wca14KNTeOL6RGllTXcp1xGvjlj
cbzMdy+hKLLCezOSzIHCN+8LEqOlkg+Tyq3sTL6g9HcixZU4NnisLJzUEE7ta1VllNerY7UOOyek
hmaNeL4qbl1YLUVzRC+oFL3XZB0va1o5Rj+8/BNXP5CPjY1YP0waFaYP1hQz1qoLTpUJVZCF1k/c
fJ0hN9Ko9j0I9GCeM+bJwOX6KbbpHatZS9dha3v7Ask1Xc6XPw0IggnUHWpwJnWU6aFUm6IpYlSl
Z+24PsomSU3ZOs5PaCYnB3+qss91/8H2y8oCCzNRKeW73PdNpDhXqMRzGqsjNKCMv/rnO8yINV2q
sNfKHwm8azZNi43IB3bWY9mjDUE0/5uMQaWN6pVUdW6fV0YYUQ/kglMClSwNW7SMroD9E61fQnjf
KtiOxVtyb2rra9scZAKvcuRD8wbGxs0iYdionCRmSJAwISVhTjixCXZKvMOfo9pahS9mH6mULai8
YeA/iyJwpXdUEkYkrmO50L6TwdKJ3inxjb8GhTY2ZGcTbq2AsrgTDwPV83kysQpHord0UIG40G7a
DcoCrXIGOKbj0eIcphTgM9gh0lF0j7CQHfv9BYjNERtXfFVtJ1fgFiLCctyXvV8OrQfD6te9EoWB
FqtDfJxIPGi+Qhm56wxOHASWw5JV2b825hEwbMfj0+qRu+06pnBtpfgyUFpOF8zpQ3mHI8yfSATI
oq+l+BT727UFIh2Kr17NKBj7zWFHfEOYZYzDJRoey8p3fuXFoawCTxrSL6gr+6MCIxBUPzfFU8Zg
cJbZK8EQY0FQjbN1SOQXEFJszJPwgFKNqf8NTCcJYLQ+bKAkcS6rdz2AuTloVDB5oZljTAsPYBib
WRRylsrimfuQovF41hBRAGFkZCY/iWgxRsAbXzB/+L0wGiQzRqMDmVFRiyqQOHW2T249zYKr+7tb
YiS56Ybf9TfczbYBRbHw7m4QNtukYXxFf25e8o730iDJVGZU6mk2S2UrwKU8WIfvBTrBsF5YRf7L
ZplbJxbcvxkUsA75+vj5/0lT0xQ8/vbyCkPSbPBIx1okMkBy2veLGjWOE4v50UU6LM2UjSLEVDm4
oHfBcN8U6zmdUhLl41TwRpwmFgTthuHmAxvBlh2Qr0iZqyM10DAD2QYNznKF1nkrxNaNTETqicNm
jhrLEmR8JIy+ZpZiAkralRq7l6P4bz4FRh0zN7rOtf5z22xxJRW/QERTvLjGysCkZUEDEkcIvUmB
K3Vb0zZew5N3+C09v8domUF24FQZjnfruR+HEy1yb/eH/tUAwoq8EybJPHns+hYrsQ62mB5Ke4QS
FaARIxUh+4T2JHKkTaUgQzTMU53BpGB9l3yaqc+cjM5RAmhLBdVD2u+GdyySg7r+nGMd+Drfym+V
spP85jmOhhQ6Tk4V/U+nilJB3sQNAQYQ0vf0qUCWr29P37Jheg8eYDJctqxxS8IbAkTG2o4MjCwv
MNptHvbqWoAC7AV14/tldLT22+QHmCWINr5FUDVcTRjnTrFjkJLVMSrOqnQE6f6cG+0JmHHZAKR0
v3RO0aFND4fo6fjd8ekKL0JgmZY6SdSxrg7etdwFsYn5UAT154UUSvwSSeNANGmWXSZvCvhhDe7H
GttRW9n59MnVEBi+cWp4xaXaa0aDvwRu6WFGb25QDM8LdxOpN+FxS1wbXUJdjq7rJso3aZheaydQ
9pdmmcy4ZS7AZrh/KG0DtgKrt2wSO4tbJB+aMlOOlGAL+9u6Rwp/FiGRbhztuNAFsTECkX0LVOpI
QV3f8npqnFLN+EWiSZ52G7GLNaPtHWHp9J4HkdehRrDva1W/vlkdDvEAFHxhtzYoUkVgqpxe72Tp
yTqc947Jn73qYpHa7C1LRdqZ7AX/X8DmCmCDAwwJ9yXvQXkhN2OBtq+7dtF/HuLFIgT1nrsyovJg
EqRSfRAcdoXlaP0Hf4ez7o2xXLvtOo/7JZmZFrgy4j+IBPsZJDkEb0xgz0bhVtrHuLjPIoI9tXIU
MNBDPs2oiMCX73tMbTkOcGUsSKT+E3bXAA4OXftAcqEjYeIYmbLxfqMie6IbQ8txKK8dB18FV78m
SgcZyfsWdE90rpCrlo/wDrQMz/Y8suQLXd6Fei67HFpPKvTRmz4SgJmIq3ZfvFnSwWwrwbllwL5D
aHm+EG2WH27szdf3lsVwDHr9rvJcXKlclxrhAEqQj0X7x3mt2FuosFwXUqm6weDa2c4gIxWRPmD0
E4JzrCm6EfTSrY42HvYs2U+l+5SS8M65ftQl6GITUiaisdvYaIu6hwljYW48ddTTSGKlpsyz5F/y
7TIGmlNEX1pgTRi5o2K6QoAxOA0FZU6yPWsMAmdxnPJaTokwpkDDD5xB1pDifh54vVR/N8VIgDbC
bf76435dEp5YBlBR2xrPbqWk1oTwrvQDqWrTJDTkoAs6NyFD/4usNlfnUd36zA4RXbRvKX5ym+Dx
+sCmKfHIZX15uNPMYvQZIzjQTUSIPyvPd+JgeVXegLd7aLiRprJYttFNla4W5pyy5hqsJkTOVJpb
qW0tFA0dN+8KUho2Hk9UVM/pG7DfKR1GGkkwr/OV+DsP9q6b/4LaU7e1JA/xXLSog3LKkK4+KoU7
+jWjVYpqIiRFGXz66M8EB4GBD+9gCI0+BGHnnQH73PrNOXuT2a5ZSwfrknpvoWeuOF0Fh2yKyg/5
N0Ang3tbGoF1ZlpVcVmkgRmykV5tRAdz37IROH3J4d6FYo6zyWIhqcjWJtq7946RKxu77+gdN+os
f13sxGFwaPGyJEjPE3NE9A4nMDDAz3NKVIl+iiuW0TuoEGmfz8eFcoqp3yCDzLoKBvt65js66y9r
rP500EOhO1BdVv/7DZRHMwBPpHQM5lQNLaqBFMtMUI3bFl7db3v1A5K/LarNoL8IHWWAD/9Ec4vT
3TlPUU2jTNBMR+IP05bl0NccKwv6oVBEWN8d3d3XekH0RigiCggVvBnjcKAyneYbnEAIFhvw/KWX
kx85wgqaMHMHgDrz7zESJoRm8NLuD5BY+KWIoFbh8NmysELfJMGxAUX8cJC/5Qy40EJHGpnoZYil
JwEFqrFeyFAQt/rjbjDX+4ddUWEog/RPp2lxZVqfC+W5QRBVH3jvVMuDHXdq0ZR8Q5Jl6O8f+cEh
yUxX8ZFFzS5m7+iznmadS+fLeqA6dN7AofX7PGF+7dg6EqXqEoSElB6kbuTpMHw6gqiYkOLcIwtQ
3pZ+gVWOquWdSijTilU57lSEjCMRwW3aki4cMDebh92qa0E0fXEbE+h5hxneVbOwOtBEbS22QEQF
deqYVaAq7dYJXvn6tpIFxgTbK1MppEhvADDxO5r2WHmcpMS/wX/HOsKJWFsr/TLhsUhrMYSi3AvK
QWZ24SjquVsJ1wcWFPa3xdLE3fNsEsPAjGa7HdeSY5E5ZOgbKLU0yB9ea4goiK9n0aOC7/yPKEBk
OZtzHbLa7C6qAkzI5WGXsVqpP3N9Ejn7ZisyANnE3bcGNnqKxsxvQ3VyNyjAAtLOVzYcQmE07RRh
tsIkH4x4rfIE+fOfhL57EF7PuqyZwDA6XQbK2pgM4KTpnMSIeyrU0jSOfzwmj0vimCkNeCDiS7t5
+dtW1+LqYdnw1dYb5WAHJgHaodrZoCh8Fy6BBSAhvXags8KUCxQwE261Ly7c5OdVKIbM/ruO9p7X
807dlZmNXLT/e9f2kleZcIkykaLIiW3dNzg6+YSF9W9wQBtgqxZMtPDHpMGhQ9gEw4oGJLmdFD/A
jQ1ePQvo4mE/7NEqNb44ZCyRzrfu5W5DCcba5IewN5dia09MBVAc6NPGuZ6phIIVqhkY9yW/8K8P
RaLx1LxjsppovJMESVXOJBU/S8APh7hVAiB2PVKbCKQYp7CcT67BgWH6nqfTCZDxOXy2vkS2L57c
tDm7Ny98yoH42BxTYmHFIZq93K4v5gD0gY+Ekxk1yC7jUmdYi0ltViWO8WkurrQd/kSsCXUhjkC8
0GloLnhQWuA0lp62QURE4UBhcHuqF2UAN6E77pZcEK32cJr3+lM+x+eKKtdRMaa9yNZTV1ZgAFi4
k+9hOLaLf388Y1nSmQr12f3B9o80ONgvtziAMjrEXrf31q6CPKnA0Bo3Zn7Q/M6uZS06wXO9lUnY
EiEkJ/oriqeIfYQ3AxjyiX4z9l2tjFtMpwZi2yt8WfaNhfogPwWiQWpLuQHaJOUJY9Yc/xsRNEKK
9bG4wyf6DSrLNuQ/oRaXAlR1uhXES2uD3tX0BUN1LgKGrIq8kX0QXKQSS+3Utc8D38Hfbi0P6eip
rXFR3YuU7CXe9r7V6ysh+9b70gY74NTyiUDLxHuTvxO4/n5KUfLAn7UTwAClXhLZXqaIJb92jiw0
kgIutfwAN1d972xBqAsVQWx0lCKvodKZXhk/IcERvI6oy6XyTfCs5/fPad06qySpSye6ehUSEkkp
EXxyu/Bl8lguOI7l49/Qp9Y2M2TN60stAB5egX94+aZX6ccvpBxUoRVf78U0pSsl6kd9fAYdP3yC
TMq6U0pkgwXidJvqeQ1oclu/50VvFlCrNWWeXEnRRM1uSF4s0dio8g6M7vd195Ptl5uGH67hxto3
8su/wfRnmUBjtQFXzExgG9Hi+DKo8p6T0P+i7urLrZT4xptqnVWkOSZYg/5UEQObjyXN/kNVMYzZ
oRd/wkjRYXD9YvbVdmNAjVkDi3xJx2qzeBYSVyItUh1KqfyEHyIw7+2I8NISceriubIRowdkVqs2
XfdYXVKGY7AbwZALczERj/+VvV2xABk0LPnJq1iO6x8nQGWl1b8l2bddnUd3a8VkZxzW5VaIAGcs
GFkHYY/ohleKx+OGlGW6UYarHP1avNeVkJSdcSl5b1YMXejA4SCXUA4ZBQihtbkUxEIv6HaPiZxQ
DXhhL5nrR5IFtz8lyMAwkXBWT1VWB/cXvVq1OaGQ9i3JJFuuAw70ZcG2hp0mNL8WdynH6pJzLMWq
n67Ntd3DzLSH27cxxE1olG2v0GHDK51w2NiwHziBIHjP/ZvlTCACbRKMDpdHyhgi0d3MMA1rN5RW
uDEiWSId4fynZ2QAcCaST8DRXmInAZA2sGICyKEYFMj/YTVJmy6qEXL2/FOexbi3wNQ9qrLzciDO
N9x0jlFcPKpgZEzS+X+E/3K/bu1VnedRsAsDtSOcvgpZ9/k0Nyx0UUSiOjB39pBxsT+FWqBWlJPH
jx7SObXmBDOT+qKV2/ip6t24v0EEmItHqZ9DMhK5z98wFcNwkxV8UiBrocgMTiRdaiy47sno3NwA
/0LK9DwbkFntlAcbZTCafwTbqwfctIjo3G2mB1Q8LoSRU78VaUxbzxqTE4rOoHASP8hWjBhfyLiP
4WWWlXQsRERW79SZtT3aZfXUqMTcukL0RXLb5i0jNqTCGAN2+cNehYprrOyZk70Wu7B1JMzbLWf2
FAEs+HyW7adnfNYRmeqB0CY6nLKgfLdnghK59R9urkiumcO0JqfyuKwK/2XHdINoFwXuZlabNYE+
rlxlzSeijObktxIjDTda/M2yqSqyyoFDNSRGqwQ1rvX+cuZhqN9wmL5mTWC9r1z+8+k8DpiesX5c
wK1e8AeHe+fKViuaHAGjoMiaxg9XYb/hb53fUEC6bI5AVK8v4IA12YIzBCmI1/10EunY4lVZ4yjc
ZqaaeFF6B9tCat+jbcS7zol/etcoqTeufFchQbjzY3uypylrOf0q0cy6A3Xkzh1ivTB5nEQZ5wkm
HzXudSjbz9+yHmGBu7+hPKt5OjkfgNiM2nvZ9uvbuDtygAHLa4nEMbSZqQ0nze+0fB4k7ZgbUzmw
KGb6LrZeBLMMBJd6Nd/ay9E65jEHAKreP+K78XqFRG439C+TyuTDrofZqaQDrpHl4sTRRYf9G1O/
joLjPKo57iEpRKHEtK/HiXhguuY19FaNYEDO8SE+tw1xPb1e3ySOVQNw8XthqmKLAwKY3AsGfwYH
FI3KmnGZ3yQnDm2zIYhC35+t04qDdEldhiMlOWEug/2su+HlQVZAEsu7bPa5lrrCuRUiVkR1ktY6
d3auifCd8o9+xksYmS+radUBj7mCD9B7BqA7UJrolPIHBnZbTtD7/utf6qwYpN9FM0g4Mo4b+0L6
8BR2P6lyrE8Fq1rUwKwY8RwM6Z7MHcFCesII4PV++fdqUJoeYXo1adaSiA/W6RAmOr4Dk3bxBTTK
UQw7liqKVv2RBN65RctFCYQ2XhXlV3WqNcirVy0Vxtsi0+Aje9gf9f5BMSS5+FMr8N4/9QkTtVQY
ecqJj8LuPMP3z3BTgXriQxvddG4a0GbeHJnQVIL3Psr18NoTHnX21Ke5+WboHBE0BuEfBWI6B6Sh
ZrEUTRWm6SpYExQEyRXW6HuECSYMHgR/ozIP+Xrf/Jldy214cyxe5jsLk8qpRhKFVBs0NzVST2+J
TGRVMaGj+IuW1iclIsyzr956ESq2Xcw1nvxVfosuds04tx8f5I7aLtP60HsbdsNGKtFima7fiFtD
Bn0XcO37qpgi94Esb7h26bcdzKe1+Wj7+48NzRU+vH6Fblck4jt7DV5uqu0RI3cVz8hgy3VsmfMC
HlUWiJjD+iECWlzp1ia7OQcROnJyrfjGap3W02dYch+21DQw7f+fNUrogsGv1C6po+qwBaQcAInf
tgJ2fdXncqin3ENTaQO6tOzrQpoFb2zZ+Qi7M7mstrstx6aSBrynSPNSOx+dbptwWwK/BYtMle6E
TvlNlcZYmbEGJtXUoI6VGNPJtmlzj4xcjVjcJPWbFWLzAEmoiGcExJjLOPQilAb1aapRcn9+JyYt
0wOBWKnWQVlgQTJbpfoz8KPDdCojNSOP7vTElng4Y+lVg+5OJ7WY9zn1HMg+mbc71+OEk9GnLpYc
cZvoKZlr2aWipQXbJZrFQN8+1o9phe3vzda7ncKT7dGik7heGjVHALG3OW5RVw2t7FiKOeOq4fq4
yIblhdDn3ZsRat2fx2jl8KrwWdKJ4RX0CYJzSp/wck37QbEOtB0UwRFxpRmLoTO8rSM5E/M4ZMLF
mtuF0r1e5XFVio6gvsGlhOUGFUDB5pb1CHs6fKCQyY7+KEf8YvnVoGEHCNmobsxOwtcvLxr1JHAK
qXzXrGQbjFb2up3nQj484l5gagyJ+vVhF/cpIfJqlrLb4XuGV3kBfmRaM+e/Aj8UxKwR2lc1bbN3
0/x8IrbAMYLR6pcJ0J0zfATEuBrU1Cb+fEtKZPqJJynFCzUeQrhu6XHZ0URv3vOhUM4DDHc3Jhec
IyoQnFHF+V28dnWFXHL6MhhKts5ilOg2t9XeHofHkUZs62hDnnh57FKLPd//kab/48cdgLLBoOh2
aQN0FJebdig4UCTjKgissGW15n2zlfEWwa+ziyC09DkOM7sJd8Hi5y+/6StCazYSXBgGp97cGYO4
pGYi9I3MVL2hvyfXnk7PogCZ4jecJYUQdMwRotAMVp4tnckASW+PVavVdRu9mKi78q9iYHmoW9MP
h6oL5J+k8Hhbyrm0rL2BxxZzM6muZ+XVox5ku+Yyj4NMGjIx7XUUJIqGd4l/PfoCspBbYyysVHbG
mukORyypW6v9xs8jvB0Qw8gxszSC24/goM+T4N9qFxX4Yj00TxDbUKbzCKXs36gAFh/fDJLFDnvp
ZoNWMn8fehnd1oPl94luK5YAb+m5f5U8eHNuOrcwdgLsKo3HmkJAlZhhoxievGKNiOIv75Y1phDb
SXDY2V+oVjPI5OwBIQUy+x4MK3Ly2MNZNRvyQTn6tXwmHkQ70tGqb9Qsm3yIVvvq4tH2fUdJIib2
pyyUMigCTp3NBXSsqWtPMhsCIQEKN5POciKvEYfuJQBfuWUBSyWxrYuButOlJxfzSSIsMb7zuT3/
ka8nBixHtd3Hkq/XeMA5NFUw0nxvepYzL6J11dlyYBAzwW4m+fTZbYeoSTXkyJay0KwIdQRBOguu
VwRbTmwehitD7r9W7l9ks2+fwRxMZdXr1fOfG9vwsAiN5cpQYC/ziR3rqS1yoWa6Dtlq+gNd1Ech
25aBfndDlNBH3U8fB1A9gJTlgLHR6gmPQDH08uiJk1feb0A7ARGu+FkKfPqwakaLxaGFwCo7I6bR
/DIR+6v5n7cVFjm4StDV+XTm7ZAnU7UAtIgMN0gNsPqWkvcDeGCbs42jp8Xscj5PkCvKoJAeSQ2J
afKpV3n9IyIozSqVNOdBtVAi59L8QVPPwayiapUv3svlE3fGa/Z8bvXVDfkoHfT9sA+6oN8QdZbc
4OBxdAyHXxYiIvfKeAWovoGfeeQ28tRwDUQFGw6NuHhP14bcQm4zgQZ8EGuhE/auD/Iok39t/eZJ
Cb6EMoirsYn5dMyg1zOKMVqJQHcfHY+XalcfyUc2Jr+abh9SxiAWUFDzQdoXofKm8EA4JVumAS7A
rIGtabwF2D+PayJXl0+Nx5ud84BDbrdlk4q5ta2eVIePeHbzP/ELst10k5GERE261qFeb92U4ii1
7jBJg8MFaUZhqPbCJ9WBtprwXMuCuSied3LwafSQ1xSjncVq7rjaQqOrmv5qocPbm2SFOpWFMtpz
8sr/Bm+U70CntvofDH1ijUGK6Yu48BudEPzjBOUsTvwCR1Nr4Vj+F9L0USEoerqfGSqWgdQ3FL5x
zSEi6ZSqOuTpNPIf5URUaea9ReRTePheqqWPbyukmYQxzNcqFdLt5dMHC4kk7wj7x/HUqcmQ30y9
zzJVn2I4uc9zyuNdmnm17q91jQC9+Le79SupM/0vgzvmfhfEaLHbAEfrvD5sEY8/+V+jgKlOEqpx
KqFwYkfTZjCxMO4XHtwEyjIC2/g45aq5+wJoblfCZNuLuX5TNvXN3yoJjQQdS0bWrpHSs7XWuILf
FaRE5C2yDY73zbN/w6u/i6fdg6wcnrl8SJArkt6zI+hW1v6HZP7WcNSco2hFNN0z8iNlQJhZX8bD
aTFU1T7am8h2LRnIaurXmq+ksPdlaklJ9mZFDLmsNkQ1UKawhvpULun5dc1Vxrhhbt5rRJkWvcFx
x8T6ODGB6H3pjJaADMD96AJrrWF11P5h6Pa44kjr8GpYS4PNwU4XEb6EsnkNGveHX0WydH/2k7Dc
03evuoZZTDg+WnAHnMYmFXcHIhvYOfd20YMYTCU8sBbu3HHrmqXxN6NO1+KtgsDrHfbewW8LhEa0
sfTXTbkelu4hLOmxnKl3XgfmYdUzDURqPXZBYGC4G1OFkCPQ/Y8igsMqjs/FjM6ZeWwfV7RSDuCj
DZXL3qxawMKYWdcYqoQJ+c9Rj9/sBu5F2q2DbiLGtndp+UTtKbArSxAuLuem1rTeDof66kbmWBdB
Og4CcVrndhDWG6q+NLT0IZ4KTrwHPjnI1DSg6rzv8aTF0Txrq1iHn5RmyFivBzyRvrgiaoNNz+vn
AD5hc71vKYyxJKGSmrlgQ6QRU2Qcv66F5khaVEY0xSBcoVmDzCfMEhv/Pe74zUcUS8AD0KyN0dmQ
SbF9AEeF28ElpBuxZXLCpRhX5PSdtKoNpuDk2f+UzjzgK8vo38mkfBn5p/JMeDq9K0VZCIQAMnMZ
6b6o5RqKO5d+PQx9rzNDdO5JR8faTIqLi7FEKKRsUUbFUEVhd37MQVJJ6cHNZvyAxcn2YwPYDAhH
KnYiSlBxKCwNYExXYggRTqJPvmKja05KaQVeknd1T58x0sqWyIoINu57v0NOk/ZBeUo2Q/8VhceA
3T5IRj5NqQ8KQka09MBrvZADDXA1hJeBGUC/PqdQQkDKj2KuM0Euf7+h6Zg2fBIY0hvf5uDMUN19
wjJ2Y+AE5Vj2Q1qD7/zZDxXNz+9wuec4ADS9j3hTVDxzmigphW9i5zYJq5zkkZhtplAxrPDfTV3o
ENQZinzGWjmPAiJ2o+7rAmnrxYyO+qWBMliZETOus1KyHQJR9aGX1u0KZzpxLiKsh4gt3mVQzati
kbi4/g/NO9E3nm5COmz1Y4UUzM9P5OOnj+22gcitLevYLfERFBDizto0ZQ76Xee1mNPh77NtvyAe
HqF19rP0eFACeHhCh5EgvJsweIiA/boimzsxN88CGIAiw+JXd33t1KT8exjKo+bzgcZp7WxA19qB
sH7qzAum6j6lsq0ns/67cmsT3ZgtmU4E0vwhLCO+zbmPiBvZBu4jNy+VbdhFnmn0C1MWVi6Q9qnk
i2qMzTz0yTb1BViYJrDKI1lykN/ekMRsRIMuD8wSzqPoWspCeBQhjtNuU5s2ARlfrW/lDeakLnDA
uj7ZyLqaE+ak2Ud7qADR9pccqw63+rVzPuH7PoracyUDYaY1PXOLdtydCGtlCNcu+xGi4g3MhbAt
j/uUe+4RRrVpjs1DYSmd1SUvfZ68yFJzxUIlnmh+eFW8dGkbdHbqqhBAjbdI13IGNxbP+ZIr22KD
EyCY4zRA41brD99cdWm3WuE5CEHfc42niC53Wu0l1VWx/2mBieEqTMZ7c9GKf8XX8mQ1lOdWWhyX
pgG+cwkA7qEIIhlhOj4wiZG47u6jwHwfqhZY/vQmR2JWfVkc2DMo/Nt0JJThlCIETxbnWKrlZokp
ToYlgsX91/LoUFzTi4F/kxNfRnFnoUR+GFuEKx+nQOYkYu1wkQQ+wF7SHhwxnIfVBCTvPwPV3cfS
JfTwNz+93CtcuqL9mKwosP5NtzpbjBqBMiNiuSJbS1YKrLvDcheVnLvAE4eSGvcFIB/2iyk15p3M
lDhBoG9g8oyTO+ehAVDyjvuQx7yT2oUR0PTynLuHZrfaKwCNmtjje8etqDraDKd+gk5+mBZRwrxl
ORgAtux5DAXhl8k1yyatgSJERUNO5IN1PKIz/MFmXUXlbaDj24Iv16C/P/p4mGQQNAnLR4psRdxf
gPuiseckLqoJ6w3Ks/GfDpbRqb476XS1KLwBAKKmGuv1/6WwQtf+6ZFkiXbkG/0g/z2ijQ3fY08z
1Yo6xNnj0tvJdCEYJfWBVbmO/aBwbkH5g6Ee3z52LsSnSXR/kyiLT6hyXJU/QLHEGuhQkH1WO9N4
/yiyT+KBBiIsMVbShpHTq0qddcBUNwWWs3gklGyBIrHcOTEhQy+fBCTiGkbqBt8cGlhs+ipgwmiu
QOIqcVdFn44GHsOl9AZeOyhTUCF3eU85TVpRbyailIj5mKyIdB6/YWzQHyegnH5FK18FWrpF16Jt
IuDdty7XhTWAtnc3pV3qgh5j5JK8T7bCTVL6Lc/HmyugTPYy3P6auusxzQ0Xvpnz9tMhEXu/8vy5
QbpVx1/hFop3QrycpSwW529ZGNYhZ5wsAYYBz7FGKgz4raYZm9JlyF85kunTa8iRXTtNs2XbAS7V
GYvttcR+TYfECMVG7GShVytT7nrqfBttRpJEzq06UDBnPYwFLoJVH/QPrvgEH9/2MFNUQEw0tKXq
upLWmzXktzD5ZsbbFwcpy3wRIYEHmKbHJQmcYSsMCOX5znsDqnV2iX+rGdIzn9IkPvGQJQ47R+ST
DP9TV6WT2PCwcvuLndQr2Oo+jjJpGlh9X+Hg2+KADHP9IPnCDgqrTjlqXQv8lkAfljJotpvFL3p7
kuHP8kiRr77BxUIm23y8Wlr678mI+H/KITvpcWozGRoggUCbNtYUTioj6n0CxHjDELhrYI7v8MLL
JXlAAB5TwpWp/k6bmMWmsNzRzRd3kOw0ObKtx/sPoZSFEfSOGMZHG53/S4gqI+0IK/RZ8w0eEyUm
k3xMo5YB5XHvg3ClAwRJ5Hor3s/rs4aCnTOQMkc0cJdSi0vZEdCtb7oY7PKr6hLT4qqmTo9W/mwe
3scj17LihpTHdpoemQ+RSk+0bp1xwI1VrOaCZtO9VlWX/BwZkAR7X4oG0ypPOGWN+rR+702a6r29
hJxzc/ozM8EzFrMKF5NFl7vQ5NHpxWMU0Vi3MW7jP0ZsDavWfyDPZE2idP/GM1ccoxqbd5/+mb9C
hLsKeyew5NRauzLfpgv5YjNAvvJxBjo6cX8lnLeB+AhnZr4Nx5lO23pB4mYpXUWOm+/zB+/FyNBy
88ic2q7Gk83Ck81dtrfiG/0DinDhZFVnXOr4KePBehQVxZvDLC4rcjks/DmVYZf9KkZzOoGAnf/j
HZioJ7kOA+k9G7vlxLf1Krtp/HkC8K2HqjJfllwTCnF10AmVzTiMZ9zckqxaFu7gPIv8LaVxwQWr
xtHo4UbTEFZiIwenwqoosjSJLBVpQa/6DuK1HTzo17zRPCStfQUAPLf1P+mFftNRm1P6GOnTOEIN
x+XuUdRH8eiZYQoi24CKpA/1dBRal/UJqH2UXv9B/xfAYdyDLUlcI+0eYcyDyoa+3et9MovZaGW1
BPZCnksvWb6DkksNJMl56Vv+O41xbfrbaJPcuoyS1UJdMRd5nMcTbeTgwZgRfFsda7szwuAwarjq
2s2/PtcdN9X+cZ3OQsH2LI4vfVynCnEMYYnWKj6jJTEe1lyod86nJM4M9bFWvyIwl7P9kSq9vmcK
32emPPksMVr8U3lOYuY1d0+HWNmWK4kk/EPOPJy0Kq6O1U7Uzmj7d9PqCngjtNQBihA8y4m9XeYA
d5nSAmPbYoyF7a0C9VB3R/27ft94+QYjyJZI0lUHarWhT3tkzBJHWhbudutOiXb+Wtfld6cssasY
gsWHL7zZEa+5EjWGQLw+Ob2FAGyge/LxJakhQyt3j4hpAM1P/fT9BYGTIQFiq+uO80iZRL+Efcvv
zEDKnISUKhR7bp/hhm4f8hcW0WZQj7+o7gpgGe5jDxgHivT/VsOp2XkR8WXhKrsGS6lvHCvGQjUp
kWNcpiLCSfmpeggZHo0i0a29eM7Om65KSGQ7mnhAE7HzyeksrrUL3o0/zP0xUMtxrrGXhBAokqme
Rj9u/PogAL3DibD2ezukGf+PeOAMWTAKAe3DPlQcFayTl5MIFrLfeZsGn15TWPcHYitzbCEzytPW
9Uj+xafUv9pRHxWcsVXlVMR8IU9fgWxcF+qhFy48BX/oosjzXcGm3fZocinTc1PoGEgejI0FJD2e
uXadlWALhhEDcs3MxXbjJ9DfXRCWtWq+ZMY/qg2qb327Wd7qaxOfjl6u3VzSjM1aCQwsA3ASwNP5
RDE9yxWGMFZAhcrzrJNkCcUkduoCjnlS/AzfiYO4+j5oIEFxuscSjXZYqRSvzqVwRRolXkVtd725
/4jzm2gOSMLiFzXg9m0gqOTXk+IXrOeSEsH9Peu0z6I2FInUB3W5N/FGp7hrQt1oNaywYhkMEydp
GhcgnolA1BekVTpntpTEvc91vUY0a9pVr2ZGHaqD1VXBSO9bxywR6LlOfCl2RH8OWxGrI+E4+S8X
Nz7+uZw6fiUbJbKNQvyBv0JavGJo+84eTPBnH7p/nDy7b6BWxdtwQFkNa6/cyCusXXPjMrmfZxk0
HqzhSEhirL3Kr9sr6w4GasP9AV8jTNcjFP+UV74WWE0syMFSvjiFwiZ1/B/RLhDP6WzyVcwrHCVF
6RwqDtx/OYxDsCd8GLWyCaO113k3O0iXQbinxj0p3x5m8Edq4Q69CXmBzgBp+PgEnVSoUPG1EpXO
IWlHMGO4HC9avAs/lUHZUFOG+T/GZy+uxBqzC8VM444xoJV96tL/yb7qobzUXJ547YKl5hGh5LJm
ZXiBd3MpB+yGQk+DF8R/Ket+dP1Of38rL68uIhIU3kPeXLIR2YUHZpVf3Wobu0iczuJQBsfi3ERH
F4mNFIddGwLbhDnbTqDWviX0+vxNRW33OtKt560FmOjYcteJnhzJHOfgMNlbkfS3RP6QrehSi2uT
aLiQIG6KFcV0osK3bcaEAL6/otdxzm6VBKryI+yUSiVh7vMQ8M54NoU5rRi3safFjQeUwCKqJ43I
VgsIxcv6KxUcIh8SGL4yGEPLXOT3LHOsHh4EnmcTY4tgShJLy6JWsNfmJzpqEgf6OAZlc/Pe7JVk
H4IVVFze7nNtvFp3J0MTvxB4oBzQEI7MukIRMW+/NtaQmgMIA5Ooi8hmKFGnO8hYhlp7dGBmfqDL
bdGMRpCU2AQsklSyfLKyeMxslqNwjCWYoUYiYUtQKNvhp4OWkLaOMyH1XMRmSWwy6/puVMHkH31j
kDd3mByIiTW+Ap2AMIPTz/TN/aDLLC93Dtxi1n5K8NZuIPwI6mWendEcMQrefAFwKFFKC8sAZZtd
jEBTMLnULuC0O/u4wXro0OWHx++FaN8upmuLsEKBQsYj48S41OyBaIhME5A3YFQFG5vRjYuR7BRM
0875skpnu2TUfBR8Jy2+kVCpJLRT3qXaWdN5LaF2Q3ia/yRshLv7/N2bFDGQ9tU7RBEXZjEFq86j
QF7FK8RRm7bQtbJHQvawkZBWsMHnS7Pr0x1ctUSUSmp4YpR2MDRCCJYVbsBuEd7eyhQzYiJL3Smu
2k0SqSDzMNf/QW8gaC243edg4QMnW1VeJrdidHJwFBCPGTRIRWSQBdcwVFhhmMDNW5r1w5JseDSB
o9Bsoly5CyaWIZ3IzmsRLtALPGf5vQf7SAVNqTlsA/+2BoVrpQqVhQ48P29iID06fu9H4bnLpnRk
3SJo29r23462hgk5tMHBuiqueh254Vs8fPQe3mV3SL0Ot8nuOE9wMTkecpAhzqNv27p9LhpKUtjF
VFuuB5r6uvIEmRNQ8SQKNk1mJwNrEh+DbLnEHP6rgzzEKRtpz+tJYK/NbrWgpujXQL+JA3Z0UYY5
UyVaa50gbgqq1DqFDA7iNvjSM28bXFaZj2crOGf2ZdtxkSwaRJex5jZebvtEcfD8PpyTo6ACFlL1
Grm8CjKJQU0YeHZs6eRC7ECdSQ9yCtXocvyi3wALno8ZyNAb/5Toe4P497/UhyZAhLDQoPFJSmgm
9vqIzBM5oiNdB9ib8UHMjth18Xp+uAO/SW3akzUNGFttqlTSE1ILceh/F0b+nM1IBurs/w84Mf2M
jUwqARDCgxncvcWXk5PhWuX9I136xOXdgUEkBVFRcK52uZCp6VKmNSr5t2f5onck2SyFYIJ9H9TN
4dEB+Cl/aDfOgV4zHbbTqjc6Ylb7RJPZE/p9M8X3vT0qtTOU3ex3+QlueH2XOsq7ev8fXrCi5VIR
Ey6qCJgvpilFWQ7SgfYVGMN67HxCySz0UWqmyk6efOknw1gSauCOeZGFrxqmUEkjwYgMseLcsf0D
vNeSvq1qPtKOJs3sdaIAPRnh8NRQUZ19PO64KsfXwVMxT0TYdBQQv2q+vTaUJ9n8Va39LeynY6P7
VqsX+FXTc7VARHTXOKcmPb9Q/3Sg5bvqXNBK/Q3murBsvbsYNXj6mU4L3RF2rFIRb+KWUpPAVboj
eSdClIGqKnOSdeDWLXijRAHKgWdQpOZ2QkdVxdXWfzfN9XOB6JPe92Y77xIBekn4doNnbaqbQTSb
v4n/LyZFfJynci5q34jS1E3k3Q4XOxcpZU0Xv5iEsuchOl4xhoQpiQL9tA3jNTMIGYCHtZMrJs/c
TK1shSeNXeCzlnARmSdiuPm7GRb9ZIUnVIFwYBFCXY45rsF0KL9ZbmN1wxv9SZQ8JyGrxjxoRGo4
0XEbwov34J8tdZWZzUbINP/5IH7d+OI3No6rqIEUPAdHR6gJGE1jCUSehpdDPT30w8GFWNgU2qcJ
ZKWqE3XKHjIP1WMeOouW6PzD0GrQ5lmimDuW6CT5bN1Tm/cnDQ0hikBYjSt5rBozueZvp/KUUfMt
eKBewEappQDZNco7NEl+ZC1wnowwaeuspx+12zHUyHoTWw/ULfL4keVhke2JMXJnVM3p5c9lBbH9
3fp9h4//nVOLuiMbGMEga76K2sOthUMd+5QECJf6kcklf+jwLzPdTNPlfb7fbZzNySCvZjKBwlZ6
dv6zMAyj7059kgajrMQtF9NDaO0cZqrFaQHziaYuNgJkwOCA4g2uhxTH1G/2aVNt4Q03nWZ2sgEg
kDr0Ma3cYNu6L9k94j3TYNvIpyt6tFW6nmnjSk0xV6thogtj4wO/EIJLkSs/eYgepgIPdqT+wj1U
wjwKh2XW4X23hbS6OSeflOKoZMhYs5GCMKQs4dUstpXQ8547ct09wzaM9eLGRDReUXjE/XPiu3rT
x2VYh4Y/mKVfdU0Ep5Wf0fX+Cf8lp8+8SH2l9TNLQKz44pJjXqUtKN7Y3u4mkCosqGA66RXr+W4s
EFli7eQZUzQRoqi0j/ZESL5BL1rut66vvTV8lvJtLKkAasabF/81UVVk7NWsCmjGmVy5zN49QPSC
o7DHDXE2rSamoRfo3ANbDtQnnHZia35PNmCotSF0fl7RZekpChXCcAegYan0XHocpupSDZzGcLQj
1L01LhrDM9bDeUek6kZM3OOiH8EoqTtazkRTGQR8QPyUgQyVlXDREkiEiwewDSKFmgGclzCONTLn
oGVix/0rzOz5HaxfFfVY6pfhLmueAtyfdwqu1b/s9rZHxNU0934TAcYGHZEvaMDHWdJGOejKYTXp
Gfgi5Jb82b6eobCiB8QZvdxEh6U03+ET3MSb+YAfoqMWRCnclaDzVvTcroZvZ0JXBpkIrYY3Yc1X
PfA79ozNdokG9ZBXKHPuHjNV8wnxV9DMNst/GFlYse+duKQr/ZH55dNZ/hRQh4vj55HYpYYXKNuY
oCCkDnM14YO3bq3J9jIDPnHzg850pYAqGenU76fCASj45BYzwzofQ7v33lleU8RVCnYwOTZcFblc
f2y83PTZ3A4tGK2TEfl+VwqkphzExjSqOcFCEOYIy/iXONs07MX1+e6GdLdz0G1EQO/96I4n98y4
+RzqV77Ciuj2kCiQEMHRT9lA+Fz1wnPANqnQNSjBNViWPVSWOMqAqKTIsxQubcPZ5JRMCXFXTnvh
b3JXHlnjqIu0UAzG2PNmmaq2PnEohdyiys662sD822ye+Jqe30ZhdBjDpTmVk8dyIw7E3b58Omcr
Lf59UaoEt+O0DdcMN7G8zQdVGBr9NsQ3utidTD1qGeSfbVH+utmS3AK6IpFVhFO9vebG/eStd/5M
d7JoZHA3FRZfIGLH0d/KFv9kHKBaxjocjhEC/KWnLh8fsaELYQZA2DfJbBBqT3G/dq687NjTeu6V
65F+KKVQrg58nbdamGJnOfARote7iZsy0AZOGF7/3dg0KuJhr9itNlbXKk4RSbl+xUdlfGOD8VRU
t27J89mkD1aXRscjs5NhNgBEMyeBJMSlsL07UsuP7f4ffImqKVWkCUGmoBtOeAdprlJN5ZVwwqbH
yPPE9BeY+2x907bQPO7uooL+k4AOFKFG8DOvlVm1DvfMhYn5OcsTXdrx4Kkyue28bHaEC5wJ+iNx
024qbetqvLRw8iTwlN43+hPoDDaRdk5U+5TyuOGkxiNEf5J05mePAGFMLBGHCltkoXI5R/CJ9ty5
Kj70+IZi2r6IKcCngEZLhO289VhR5JsqOeETiE8iJeXMWRFUQCY2yXn7CRVwULJ9bi2j+6TfuG08
MZ8mnfzUk6s5Q+Qa/MkTAL0mtv7/I9RADMH0yuav40D/jsWVGPthMWwnLw82hPyPjyNI2VMkQnAS
HSL/tHLgo5Gqc0Z6i9b7t74mFLH2BnJABDFMWR5H6JM/zbiFNKa+mzq2GbYFcjzvNDaZeW3PLxzP
SI5gLhfoEMZlqCQfs9/jnoNnMtQaG+8qUM5hjNYOwLRYropYiJuLPqXQtWwY5xGVapALt96zOB4E
HItGN+X3a5l4lpHDh4Pa/XA5J6JlW6hjd7tGJO+StlhpIR48NbJaaTC9BA5xdaf/TDK8+vw92Iq/
KfCAbYYS1Nanb5yR1uY+sW2gSqBmqKrKVRLi5ou1QdMB08Euw1jH3dvl2u4nXR4RntFuaUj3efEq
YJyJcnlpBO5E3+XkeE+E8x/QKAsNP/p3EU/X02nIB/wBpKtiUf/v/QxXYOYMGjx7pKfu2aflWnGM
p2mUdbtDBXkIFavrRBQ2gLLnMNlFiR4tYohz4v0R7XLYRVjsuTE5VnHSxUT3LbBYVfSHDY+otLPh
avXV4KGIW5sxGNN13cicn+jDmURq1Na3BcLf/TES+EE1H3J47eX1cAcBwa8GYEQSFjVAKFLEn/3m
zBKFWcDGouz8ejT+nHyDeR7jFfNEinqFj+ezTEsn7Tr2ZdFPgfVm3iHSbBA2TAdPUjeLnfzGDDIT
2xDOQCyvuxKrQp5JzQ5JDhys0fuusrYcYDluT44EkAsuWjJyg1b58iXrmb2AJb4YAojCtufY8rvb
fll+M0SXECQNyDLl4/izokhAGJDLXT4fP5Uwinpg7RgBxZN0GC/9/Iuje1ufMG3IZFKQJa/eo5iw
Bv6KfkLvDroCNmGGxDdZvFEelsxb8i4T3zqqOkbUMySv2BnY/y3lfTmwVwzk7N6XSDT0utZGyNEG
DGR/N7RGrTo9M2fiJ9oMc6J7o+SXe8T81qdO6ofxp+9EpJmPIf5Z93zVragD0xPv8y2E1+29YdW3
/RPfIAc35ukThlRqes/wt6cacrFl9DFqxSxy5Mvk70+qGB+M7DeMQvsASWEY870X3dZy6GZpIAMl
fezQNNBklk3UwL2BDzNJyUST+FAwkUevz+0C25B485NY58BUcD2ezNz+tXcfGq8r/3X0CgOYtZEm
b0RdyntGapvV8/cz5Z3Cp8zvfYhir89urjs5hLN/gbGKtxxYFBJVfxcFHAHU5ivTlQbabyJ93hPb
ZZlqcb+afyphpoHu6dt05N31M7OIagqddpnq3W+hUyapJoROCQQ+JWBieV/Vy1sm9wk65sHqoPdE
3QVHTflEO4ou5KhI91Bu+KdFQjn6TgC24AhUYnLMQ6+H4VKO95N+Z/+xS+3K3JPIDdq0JVMJv0lg
IsOipGUDeeCcMY0R9B5YH6iNjy3IxJSdN2/Lt02NX89+ZzrhNev+AHOdoQqi1McRrrfQqf8xxzLz
oz76CMrhvnbWy6EsUu/iSd3HaCFDMhyNBQE/36waiPNP4kukWDp0YpPkXoJy01r7nlSqJjMt+WqH
t6vr5HRVqa2LWmG38XLpAPmOfwQAJRxB4JBEgfjvdAI+AZYYFB2E4ruQwJ93May0JK5MNpUr9Ddt
qSVVQXI1JpvViGIzmbkMvehVqHAMPc8tKO71vv80Rm9mE4MQ90VRC69YV9cAaJ11xkOdN2c4pKRm
XqPTCeQBWnizD0+iPygL3/8Cfrcng0WJE75RYVggUC8g2Bb6UvCBHJAvApQkdHrD3V3fjgXeznMM
psO8tye0c78PZAcmUmupLI6CDa84F1htAaSwYYXZx9IaDeiJA6uKzm5QCaAKrxegY5NlaTcNbzRs
oCWd43vV6V+Zfn9aTWL7o6+MbKCK5TWzIL0eEfmTi8PgM4HuZEgbW3LEFntxATpykCcUscT05oub
Q3ASQNAKNX2IeeNohhtlmBQX0IEpIuKCdplbX0MTNI3Vqgj5WW4hHzdetXZtCLr3hGWRv8mpZlQX
p45sGjptFiWUnfATCIFrxUxm4l6EJ6QuKIZbbBZUOs5IdUWwVmpUN9mXsdVa4OB3wOCr7nOZXG+F
g3Gja9VMCTLHGvat2ujsPiPdKgUXxjLj3myAjpwLs82+8nn05Ivdn4yqa5kxrLSBlWW9HzB3V6rL
/gB/SRH5suFW6IcSpBxFvT9QyxXQZTNAPlXXbjMuJ0HH+Td44oHp8UUxInp2WOtOf6G8bxINeI4H
oA2/QFU3WH1Xw03z/lba1a/05WBDD1YjxHiQKJq0FBq/LadC397v/s40ujGAZHSAakcq2g7I0OqP
x3XfgAwjr74Gf5vqRm00jqEHQkJ5pNZi1MMYwYfhIbU2utI2v8Vp3V9X3q/0cB1iwve8QGAanXLY
CWJv/ahGFIsSIFXYnb/wDt0qbwoOj3QS+NzPwIkpKWoa8AzHRvhSI5o7uR1VpOflotro57Y4bXKI
8IAuS4ClseImhCrk+z2cgHX5rxhJ+jkFT07pMxkCh6J/SAw9roZXjO2D1vyS3FpkPRo6xd5AZW30
sfxtHBrYDS4wCFILD8G91Cy5smawnwKSb5FjmLPOlHf2Kaj+2tGP+9Pn4L2jIG2Hj+JmpCsq4RmN
ENFgMYiGscD7suF3iDS4eNrTmvEhJNavlF1PW6AU1+Nh6feO8uJglQX1UW3BOTtpLsMSjgGSyGND
p+/mZz9RQce1G04be3VJkY9zAwx38eRX1rv80VluC6M4l1hSNtfKb/8Xkwbq/wH3YrXNBqZmlhef
Ed2KPLfLaAadxdyeg7ii0KtfkrmV17f4BaP+li598DLJa3KSa330zghs7esOjNaxlKty98+zieAY
gWzjFkPVl+2BGOT7IFIoM4WKzaMIG1Dx5o2mRecAEAcYpKyMSU5h1AxH8fvDU+W56FFtAWkYznan
0Tf55lCOr1/D8ThvIRz7t/NbyNyIRHsaeHp55benHPLOPoZtLjQVDSQsmJMCKLpwyhoqxhk5+tSo
d6dzr/2ckvO/8oTnAkgIV0NiEvTJvNSJlIeJVlz3kcuN6oZznNPe9Oo+R235NLEVq1C68zQWh/sV
m7ijbtD2CRHiefoz5b3ETJ9+qDV+E/07FKwVqXGNOg4AOnpmJOz51eodSJOs9R4fci3fsv0cPk2I
ew/7mlG15hlADeObqpqWuK3X1V7L/OZb6fw4De2DU+8vm15uMIoj9VxQceEJGuwrygfp0YFtKazo
zNwwJFCRP6o9iBz7wTLgO1anzF2BbbcQrTDJSDU46qJfs8w8VBkwU4KkfpSC56zv6RtqCKJPHI59
Fo8adAsS4S7RUDJUgHlb4A31YgU4HruNYAIeEI2ccrSawHTWlKOF5YQ6LWTuyS9DAwA5sey170ap
UY04buQFRjbwXs5xvW3Wp5V/b4YnSjxu0fltj0C11LRPH/jVu938TJvG4V70KFH/apEvxkp8lgBr
OQoamPfMHG0fcu1jQ4BgMjurY1zhOrE4L52lyKF5jbzEqqWT1MmZaCX8h1MPaUyQSSENzIXfRXGY
tbzOoNklrBgNGiDzBXHwAtklPhBJRpo7vxN7btCVs1jfheNOEJgKONHFhavaHsdcD7ftiP6wv0p8
b3GTToPE5ik6fIvJ3eTkvTE2YmL4BWJoqcGbLRQ+FB0vCo5bf3h9wWB0rxPGuohbPl7h4Y4ai7Ep
uUMomSWTyizbp/dYCJCE0OAeqjVvcXEeoxFsyfBEFtugaa4i2tERom6m8S0AbrpqzkyMrpgJl8oh
h+RIPxTqP5RsrtDfzVLF4tqx5bg4LAJd2RYHc0e0M0y+uo7oaPZlfFL3hp+epgsRcd9D+SuYk5/I
vKlcdYOJQZQCqU7vxOk1JSj+m4RK0rPbLpv0lUQFq4I0ViQjwn6VCBFpT9dhwvk7ujrG7OtB8YPv
m3zAfr+EQWtxMA54BWPaK8ZuZQRu8YWizgA7cS4GqsaI7U0nv7NxPDqbtUd/qG+BGJfBI3XRTRT0
jRlE9EXt5S7oZPcAj2jSiNxcMqBPelw6Fwbvfn54CMYVcBRcRaOfOpvYOT7KTLji+BQOQZ9/2TfB
DXB2hIBP6/1y+Jg1VQteSLns4nRe8ncffw9EJ7tWx0zJREWDA+coRKjBChQQMVFfHP5xsvFPksqb
C6Gp2bVeLgpDpZIciyBwpQsJlA4F8QCEO9pGFrE8hgLyng/KYPMtBabQjPboQ4I2G/kCy/rQJ7Tv
LXynOpKaSGAqWrr2CBOqERoYSVtPxbae7zNanho06sTQXSH7IkJpSDau+bzdy9HmCMiFFM176SCc
M3vYnAPTjKyoOpmB33bk/2Mi1kihpe8UHbmbuYnUp452wQCob+85pwphQwKi98Z3caIiosYhoh3d
XjIcc2ACShy64hn064m/xM58vMEU4DwvU1MppPLvnDEgTAl+yut2m8scCrbAwHwRGRWYHVS9IyW5
yC1hrZl+gdgnw6THmKPZwSBMhmbeGjeMeVNo5pk+NbTtXyoULqycU9SVyXlYr6TUG0MEu7uUoX+9
sTIztyfu+vhNaPpe9wBYKBRmJ7rE/FMgOTE1flajBLU2+0Fs2Y/S/cfIkQPpF9YeAg0n9awTjhIj
7A94bbMofF+C5e+aWKQmC+yzjiUSGJzs0AhroPExO0LSJEtiTt/3f3PfX9VW1bMXnrId9QRkjccE
MYlID+iZtHrMQJ2DAUxlup+EgqE2s9/t+UTuh+w6o7gkNxdhCcFZVFEdfmgmf2d+H47Nr00wACXz
RUbJI4PQWdp17xQFk0jP4CjX0YPB1JkUzfyrQXwNwwfXIvlTx9G8Nqhj6Ea8qs/JODqsH35WRC4w
FS+NFpTJM9SXZC6oPwdGfbyc4/tAlny9FXpk52qMVsnjaU8B67qhX6ajsd46u5vcGCcstd4j/mVm
k58HcfOwzYJEo1M/E/syYs2adO4F0sXAcs9baBDD9A52ElChzuLQaLWmnET9co1W0snHOeC5oQnv
NobDy82Nr9X9ZVV86UnFBp0Q9zwyJ/ySMfeS3EmMtFGATi8YP83XeY0XySvbpdkFl5TdhQm2Mtv3
PNT0LnWOXWCbVcklQ85iUljMpu6eV+opQHa8q0sIpp8LRtwveCkP4EGaYyaLkTDpb4Rr3t0TQrRK
TrgPj/QP0HM6Ej9DSrl4F+9rEdE6Fdy5xRiUa5Zo1XGZUjpvwu/geYKw4QruXhsRJWO++gi1uv0G
Lw7jknEAmEBqYQut8BH/adFPxCD2bUsDeKUHbIDB7x6+PGP8g16acKdsY7mWPejHQWMXkw1ekdNP
RWyNTDGYhf94kAuVD/rBjczwDbW9LqcIBmMwyU7QEz+6RrFqSLDDTWOxfnuVacwO1/679KdctBMY
bj3hGE1huRF3qrYtCk/MGFryJy1OhhS2Fd1bryOl9NA4ZBDbiSSQ0+w9mhovM0dQ0CLCLIQvoVtj
Z3IHo7l+EY0aXZnivfnbMjKI5VfuYvvAA7d/2jxsHb96QU1YgOfi76QRiLu1T5Klg6YzAkte0WYV
85HzCun5Bx5nd2/hnWZ2JdOTM6Gr5ZGYRdzUs4CgkTk3mwaR2/FoVT6kyRCBM9yswsh1eu2m+pDo
i2FPTzzJ16gEuns+mhxgZ7cQ/gOIGJltwk+9ua/mAr6IK8sq7xPNqCBYIrF1qQ7FK21N9yxlnxpN
zpFAQuLwsDotdc8AY6RzrWkpFqOAji6zciDgWrtmy7OnUS9b7YO9IAVctIcIOvZj3TgzX/e7qCV7
0NpKMXns2ZIDkz2Ld/qQjW3bBegOUTRc71WlNhYUoAMpZ+ei3X/3JiVYvKgoMw4qjbjUiKtDKq+3
+EH6DTIPNkf006724L8XXhS2izWlaz2zXbqeMdv3Y4CTXTsxQEb21/EeMzTtnSiZivQqsot4xvEG
6SxEsZnfxpFrQ2xMkgDE+z23G7/ooZF5ba2zKtpDtrkpq4xuBSu4rcHaofjq63h2cT0EzHj+hd7h
BBgqgTD1lSJ1NOST6jFKF92ZPhureZj363bzkWnBUq8hBqkTy46I7M6Y+pVn95yAgbppCt45wHXq
pmLfQ1UJyVVDDenymc36QxYp3kM76d0YCARMBf9T2528LBwOfk/Y9GkuwNxmU9ZcHa+FKgZqZwva
Gpp7T16W0+U0XH5ZAJ2qCms4wOaOthE1f5EbnMoTdPiHhpldWJMAkolRT7VZzrr1+D0oP/q8EihU
q7JQwu/RFSPdSX9kmk64SlUxI/Bdg5fxucDSaNsNGwrgnp4QGGbHpph97dq6rDLou6uPCCxpdM/Q
CvS0pKOFGou75IPpvR2u3go2lkO/ujMa4UDfZGLmU7DDAMTVuyBdpBoIdj1pSGAwp/BdTB1UAv0U
xVbSRT+ua3tBpHV0MNdiDOJtEUp0fcdBbYrH023PDQbV+0qcDrsNiwc0foiVv6MZuteDhUjmVuiF
mHjUXgXgJkPmMHGbfE4iNUgEeekf+zkswMi8I06UAoVmmvzDCe84qxIbMHaP4UM7LHTuUbhACwoZ
vfNGkkKk8GmXEMmkn0zWUAtij2fbv0S7xWvepQZ4kTFM+fdr3pSKp4Js4WaI6MiotYmFs5d09B+q
tNrfroM1dPiLRRq336yrFdrtHNZA26tT5ElvRFiTaU8ovIYPoibtAZt1CUkWTF6jViOtSaFVrwX/
BQrDWAlwCrGX9lsaXLFZ11cHpPyf2NdHx0JCV1ef8ENU8oH2CQQ2ZYr1c1ZksQRRj3mTGI8JF1Wi
IQ1HKd1DQ6N0PyCkcNR0uQzcIyAet1ggKEA9Kq0M5ADJe41Pa9jusjE0hMmjLAV5V/lpaMWq2iSF
yKKQoLwixSHfksDugE6D6WHXBZAa1RI26LPbBj1vV/PUA1xm3BkjlHckxjYgG14yk3xHfphwJFNg
iFPzH1mI56sfc1sRLhJCUc/FdScnCyZiMMrTQLmoakxkMl4CK/M7EWOxiyDic14VKr7UY/4/UAln
putKoBuGK7n4CaQCcEDFyclhhQHy5UJvAfh+wbVMkssxmoh8S7fyni6byOhr6RGaMoKtPW7O3HWz
2CxU8tqHPsb7mS3L6lqWzzeycq783lgUeAy5wlNCuTVAWP3xg04Bq7tntnSn2dEfH9sZYaE6zYJf
EzZEMNKW1tHzLzJOztD32PgrC2YBeW2LmPgJNKpBYdMbLJVQjI3bfkaMrdcTpWVt0EOVnLVDIkix
TVYdzl1gCOsKEcm7fSwJrXuIOJxj9I2zE3P2OsSUxfCRQE8P9oUfLl2SSGd4bNQfoRcLYhCZVJmD
qnxpQIlGrRU3ZaM4nVp0RAsYHgv89cXceBAHd2iGBoLTh5qeFXSYNmNNlOwNDPWDB9YAHcw0BVgz
q7Ml1zJhIYygkaWwYq0KJ00NtOT8WqVnkYpSLQxG96zNjazL1V5y2dFKVj9hpv11b6D1HVHZ7qSZ
EyARN0vh8+9ON/YsVFreiorlIujt+XiNoQNP4KLAF1cr/1QNKvAFFkE01l/4KEU0HcK5VmoZkSXE
rhh+mrxOwn9qt8jb5w58zGOh5OF97YBGOP0Emj9U06F0VyARViP4DGjTinj7LpTpVLO0qBKYFk1R
vdGVPziKf5G3tlkNStJPxov5jzywTbX4UO9fBWZfG3Sfn0tlBBEzOwgG8tM4TejByKu2dNCvNYeY
lRkk9wOT0XYmFI55AfJFrrB2hgmZUSTL1TzSrjjQyD/jwdPCucML6B4aei6uV5P6rX242gpIS16a
kSqHtC9dHCrOGNqhT/klgIIXDSErbB+t/eZxFmXirCLhVkzCpqIw6aZSVzNAupb2RzrLnaiJgk0c
z7mDhcwn5atdspymz6u0fHYxVdLekqHWIqflWel9MmxSeBm7eaMOl1QzvQ9jBvJlDKrQLasXc0oC
iWyBHt7lgLHyoplZ5F6vds9kPi2rcyPwgkLfqnCY1r4559TniIz+zGOFn/mEar0jsoyy6qLULHWa
+TzWdqsPsDAjt/8kII4lP6cV90Cw+vJU84UO6q3QF8XAhgAq3iSGceS19Y5ctt8QZc2fiaSo4Et2
OPnS5Kz09kRFSkrPk0IFp7LaySaONnqBvn8WpHGs7VB9y8PWPmE9/6se/LluzmsRuG6agKsfzmNU
qSDmwHMTDMRvO+pmM17j/az6++rp8eHpIfuYP0sDePP/V+SGfYKNDbGjaYNgUt/+1oAVVjyc7nsz
o3ddql9hCT2Imfr/DArsJIPZ0eua9SUDatArspTiozppNLigOiFsmIaLLi3l7F73xOlwf5Dd26Ad
ohMfMJbwVYoF1VeuHe2X1i2wGUKZUur2OqJz8HQnDyQNobWKZpXB/XW9AqdZSEjzKGgaS+3ipL4K
NduChS3B+zMf/KaYrfdH7lRgbxHZZ2R2sLwwOgdwt9eRK24ZTbCXozfpsMpIfTMHR05sKcScHpYh
/VaNQFLgBT87eARJS5VbWUqUAghFZnolGVbUIyV+pbx8deBtOHD+9uHfNti4tj8Q76615Lv2gguy
SoliQICqct6AgujQsa8qCdFLvPmBvvjz5uaONJz63+aLKh4jfGiVa7LTG2p1850cPLmpimBO3xbT
D1HtvrPqkhEhwWdNCw4cTtMD8QIy9Il/gZpgLO2oDxi1683P7X56IKvTRv6diPqMD2TD5Eadv2Mo
bF6gvFjiEQnXCAhKrajNpMGVt2h136nui3Zf7tKXBfQbCf1RsEpvzsXiJ/f64Sm2dmZGrGAtDCRT
YOdkJ2Inpy4c6LleiRa21KtAMrFQJEJRCRgzPZdCQzr33lxVzM3PwRFRz/WaIuY0rwG/KeJ1nwqC
fSYI6t8gbbG8+7qQ817BdznzOful2zBwEcSryYIUDdanblWGVYHn69ZnU+Binlg17iQkp1Ark8UF
7o/rQC7tjI6cEQYBQ6WYdjuuxWV3+n7P3Gow8m8w2mImmaG2aspc3kl4Z9rhDPsWj9IflSe8xqeX
aJ5Uo6n5uJVUVhDs1S8X/FaTGfueIDv4tqMbNN9yF6mxaxH22XevUs9ub3HyX8z8wEK4nhIR1Sau
RyvAd3xEygDaGv7BpB9HNgu8WgzUFmJmK9Fu63qalo+FX308SmN6WRNldhOYmlrjPXIO4nnXh2wS
dVAiQa2QJlPRKd92opjSOSMv5bK7Sudc1aeX8P3u7Q+RrIACp98sG2y+Ou87xUuz847JpsQ2Ejpb
6sdeggH9ZlRgeFbcZGKhpg12PsIGvn9ZrKkcxdLvaCnhEiqwUK0MAijieBG7JKtGUewNM5uGxL72
we/OxzXX66OUVIHq2095B/ZjUTEFHrbnPDIX9HnntKHo8tCNeZ6Ri57Vx5lYTIakUH96xz+BlQk6
AwKa7wD+jxIdpfdfDqB/O3WTQ0tqv6j/Md1xcY5KYGkrKp1GkepQuxZlt3W82QU/TxRtA5JscpCw
Va4nlfmFEuPNhSseCFwoy3Dk19af91eFSywNy9fZFxHoj/K2BO9HSJ2xXaMurPxTL2y8Yf7DVDcO
QNsgbpZkKFwBWvIZDnTP78PaXTz2iehU0rTEwfqF4BtkFnvrAna5K/3QYibXNG8pw2XZ14FRg3Gq
eROD2hEq4nN6uNKNmVsGJA2RB87U8GlJraCyB4Yt94FoFiN8v/GAkMfLlOFLy2tifhOtEisPm86L
spjwIaVRc2NWrVwecix66tA4HzGxWhbUyB3NZ+CkrvYd6wJ3nO2h5Ye/2Rn+bJok9WeWjGSA2yQq
1hgpmzthfP3GbYnpBqjVKqSm/AMmmVxNcm9OKEv1RPPXzDN5JXvfKL3WAE4o4HMRCrLkTk3bvwfA
sCxQWe56hEQ8EXzxwElILonFxmu14cDXQVxirb9C9UUWZgbMWykghFmuGyxyYIgJBgnHtMCM6kma
gLV83ML/lpKoMnm1IKlpNXrHnSm3LCE+/2gkyoeil54rlAv7ftQr36ERd7koRJ5vIxAIHTj/hEcP
pPu4bII2nqkDf2FF4x00oVyFHawjzgybA+gvWI4nXVTjMkjS1KNizdR8lt1Bs6OuVaH0Ia2OfPLh
A6Zq4cFQR05twd8mUO/ZCKEdiEfLnkQKLNwJxh1qiFTh+DHwbO+dYR1QWSQoa5dcFvS80whyTefw
UXgcVuLfGCHCLOqKusQ+kVki47bcFIwYQj8etJRgDnJgVdH/L7EZTl3GKKAZ3caHRrKXVfKG0GZR
JuIbfyif4zuQzIi/qJsrbQq+as0jdrIuo4A50ulgFJXAC1I4pKf6Hzq6x+/blmnT7ASyxnKMM3uC
8icFH8xy8wi5KHlML3VzlsvFMX3I72a5Vp2PtLnDOg12FJEzpoTkSxalzHl+1y6OBGvMDo+UQ2KZ
ODyZ0WvFWYuO/JN8Rky/KTm8Md5h7j5TwqQFiXdIMTgzYMEgZz4NOr19H0JtajSgtO2wWbqCKVhD
DoPiqvSS2d+35+MDwTuSgjc0ffFRAy2eNvJ58MRTH/wU33RVnlZgdYKFVjhCjQD4J8QfL0eVaZIY
oyXcCg8Zfm2+ftBnI5/AAAowB+AnFn3RFeTVThJA+xFygwsooNOMBwQYjxGh5UWYHrMDzLD6VP5I
u1TLhn2iG0N3Z3QRnzQsEQGBuaqSbz1Jm9DlpKaYDTj181nnRnD7lrRGwHnzqsdIBnFLnz7/QT+q
OgnQrLFQqd6cxHuDdcl02olH9Bsa9XmddainFrfSyaJdWrNSSIgo8Hdtd3ioCnw2yhLit2DwKvw2
QWZ+Y0+7PVL0gWvOcbqXZRX7RVgfzwHrQv8vYfkHPMZjZ/rROWJzwxNjxo7/dP+FPTuc/PqQDZrO
+gN+chScuSAKejmZ3E1vtlbqi6rw7P0woPEIIVYsmCfU2x3aztqnFp5dD5DcF21q1FqBxS3b3aiO
NidvIcqoR9oIbhIiFmRAlYYo6AKBCQEG6CLGdFtFqeRef7Rc6tM0sPNqPjtcQCSJMZIor8E0zwf9
ZbNgmB3UfA6/R0ZXU8kb3X+feGnRoIFrKqgiLP6JvbiAqevdHy6NaPq8P2Hw5TlilMp04gC2W7TK
6MiYKOi8JrlTuodA4DeJtbAIqx44sSON/sE3kw3gIsQDpkkA+Zx1d7xkZ1DoY19rKgjKgoUFUH7e
UreF6bLVMa7qu3PaDe/3jSwsKN704CVgN9Mzmvzw00+BNbsW6VKGxV41uF54IMyKP1EUeWWOn3Aj
rIQeDnt9UMMV1pN6ZOoBVIJ4PsmvVHQP/g2D5BV0jw+fIlscOGl7VLtKMkEO70HouqbRzgFh0tim
J8B1IO3O9+08PTLkoZ3v6YuY4qX6un2DQhHTjLilkkCzd40/vRjKRN2MUDfkzqwfUotl4CUlc9NC
zundguHw1aPEfeHl90T/vBQdouHX3vKOMTQ5mzpapYb5thLEv0Q43jcfa3sLjW3uOhgti8NtAnfP
m7y2LeIn+PpQfnEHptlUUb3yKDDrHxIk8XlJq6ueCvDepH5TVZtOUUIJ53GDsznJ1foOKXM8zKO3
iBSFIp+g08gdWY+y10QBzvntNau1YYcZIXuQfG/EXYLNtptOB+v//aRBjdbnwkwWh9fztLMFJ+Gq
EqWM+krUB8AFKlMLGy36BLBrf2s7jiDKpp5/OxH211C0AuD4lTarJoIrwhtMZuY9tZEgemAyzLAF
aNhw0b2P8RSxmlymr3A/7nWXoRHXcR9w5PdITKGE33y9K4tAqnagyoIHyIgU6uayFEyRObpKP6e/
i/ehtAbmg2QlDMkZcTWPQE0YjSUtzAyP6xRd7SFVynpSxoMA5wZ8MZW3fh1Ojia+wAeL0CE77/km
cIhwKjonAAGiq7rReBzAYloZ2mJ559L3XE0kFJZdxxE93n9vLKBpBhEGG+GZLmQL2pG5WnUmiDuy
8830YPWcwbfH7QZb6v8EPV8mYJJBzQUf1HvjnV+RpJ2alw8/PBA9CkObHUDQlhKyM/Un6MB86w7n
z4Z+Iwah29LQRqnpx4c2/1I850Jns6STtvzIcAfR1rA2HfpOn9htqfQjrAh1vDza+qv3+vSwcpcg
trmwYJ7n6WuPgtNziwZMvH2Ji/V8vIkYG1GYTnzMvqoQNP8GJqMtpL0DJGgJZibptXWBYkF7yAU1
9uagO+yX/T7xa2vRjGsuxAQj73+Df07jUQ7jgmCSIa32KDOLpvTQ1jBDlM3XHJrBGgxysi2Qqebh
cYZUePEHl/4muIeVncRkBbFkcK8LBbxeQoVzYnidBMVgM4nWo+LlHy0NLZFBhv5bfX57xSCAK9bt
i4EQ/dgQ37f3vs/sNReDsUSPvmyVbjjWmA2G4WA2G8Mcom11zm8Qc7DzpViA11/sKNEMhMjJXiOH
u/rlm7Xqz+1UjNjgYMXITDy3JytkyYq5FeroTTU9w1sIA3AWFgpr2DmSbJ2kNvp7Og6onI5Eci0O
J5slJSyZQTp+a51nKr1dD6M+KiKMtEoF2Hk53VtteL5osnubDIdiDjjGdWJ5I+QPbezcUj7umrit
TlxpjC+qcuLcFspTsJhtBvVwplD9bVedA+lIZZSQ5sGquIj7PfJ2la4he18vRmCpAZ7xGwVefPxl
LLrU/Q9Aczicsevc9kMOOGh44wUBT6sSUoR63ToS7UHkVdeEKKY3/oFA/jEropuf2J1s3tQ9tq6b
GvGqMBwtfa4VMitwuk5jW1FIYj8LHElmdjW4CVPd4h0542UckeXNUTVU09Pec4zAsW+E68qL2L9W
cXdemvlBkVm/xjzAFJCfbs3tsZHxt+kMX7H+q+v4kyqgOy+MT62HnwF/5Ss/yWjZ3QrFGDIi5BXO
Q+frF+TYBe9w212nMJVA7HQBaR6/+UEBTKuLti/7pJa7deBmLsDwGkS4eG5Jxyibu/TIdmLjdyPW
x1CVM8ZvgLdibaq0uc6TJA5DMF9US670epS7refpgtOcfz+sxewbRecAgb1CE453gcHZG2rF5slf
zSJX3FEKzBApF6bxQTnXcnG8K0UECRSdqIJyfjVigXYiUNioqm9vqAAaOJ65G0pqUFHirGYbJBAq
oGSMikWozyQPb1Gg54/hqUYikEWzzTOsaGu7P3x2eD7WV72DNRzSBXz1Z5e2UmVaABBVdikOS3rr
Fmki4qac0iPmcw1f+oHcwgtGAX2iM7auw1719XNNWsz+XouWguspElEbXs4JNZWX1p/g5Oo8G3rN
4RiMhY5yyP9v5dJ7Bmhllgy38P+tDNOZRAz12Ry3nylEj8VKXQCROdE3gszNj5jPGC0gd06r3FBo
YXf38r+NDmZ4v2pWDo5qx1BhwvMkf1lhksbZRSng3MeL2VifDTSusMy0S+rZkpUBN280JTq+68mS
iMLaVuS/s7nfaHNQGj0b4Eg2egkOprXV0n95xfG6nh164Z96bLnOG1sWaV1ZxOOjan1Y0YieJ0Af
IDorwBWBg9Ncv6WxWQl+I7R+wcSYScNoQV6MHXbGddlUdsi2XMls464C8dceRblwqbL8Hxf5AdFX
idwK+R7psPU1JvdttVJfx7DiYfLMFeve1WKfyIXHOHUZfug0Ldg3swo6qeNM4GMmBdiY8GuMzpiV
h09i6uG3BRTAI1/e9vq7uKg6pmD0W/ljDdg1sU1HQnghXvAYMQUaf2Z62vUui6prnLBAA7ec6YNO
qy0ZruwQGYtv8zpAYCtH1p4CBvFMu3f0kA7SHq1xmy6eYlQ3SsVd0+Wd6Y8R1IK0xFhjslGqbsBJ
mGazAvbzjkNAiHoNJAgNgD0YlNK7hwhX4fsIZfj/cWYxwz9rpRcP9qusKspXK/ui0CbPCZTckTid
mt4McTL9Tvf25zLvI0VeGyqhBeNTbzZZmrP2fR9btEQXaR5azj4CcnpI/o6grG6miJb4fEjFIWWQ
sSEg1XdRpWWSV1k0hAUoHOSF3zY61qUGbHH7emV6PsPgxJV1QL0bWmTCsvG9aV9ScmXIu0VMgoPp
sir0JdqzfBs5mGZcd0F5fuMYECbYk61auW6w42W6RI/ztlxaeup5i5wk0k9OAk9F9t/tVMPPtXOa
pMe9lTttIw1CfspwSHS/8LaIPz7Yif3+ZrdEX3pu3k7T1JEOiZ47XZRqROePB/Sb2ELfJWtsT2Zj
kHgLM8X+VHvjXHUp5AjM6quOE7s5gaWN5QU+RPksGERVzPuHJ5jlH7m//ajzbo1XqDNiELjLJKYQ
saZths4jJ865XoQQXDkhJMpv1lOHTrMVjnFVO7gb7bVyKRcdY0wXA662URBRkpisRcUU70qgNNjj
5CpRkcFVpvFdcdDYZjEkNgbdeJi9XsOEBKp7AmRvQXCuM/cCXbGncWs5hu5X8SIeL2Ytwh3UXcWE
er4vc7NgiXssHeE2eFtwJ7UUiTMwfCg/OKVhrGgfM4wdJYYbsv3SOEDGmdHSxG2f/5Zz4Y+30Gd3
lMQXgZSgi3y3EtvdU/P0SdElkiGqI8S4nwC3T62YYbu6jxHc7l+zKa6L6rzCM+OP/b25FOlk3myZ
jo20LVXEvNwAZU8zE3Ft6rsUjIhr8K4u7aPjjqXeRkTlke/17ud2egwj+XuN9ncmPg+qMmLU8pIJ
X6UKiNAef2t5/bf7MUcE2htQNIM8zSGgR9D5ccvjltdDulsTzRALBq9nB/hIxXeJJvpJhMTwMn0h
tQokonTIgE+WkDtZKjuiYrmKic1yOxHwKpfwINJ7ph4yTtI3ty/Ql2nabf7VZ1whesuHabs+7HXy
KI75NWhDqkckQmgB/PLLKwZGTRV/bxoomKJV5EcD1vTJnmAk3yvlJOcLjSH7R3OQyAg6YATOjdpy
oPiP/Xsi6trYM5YQvKFunBWtlfkWbbrzGZ73nMlZQb6OjxrPAjmFKjqVMnRsik7AFuGpLF1qgRkq
PHRBK8eFqx77yiCTuKbfs7qUtji1J9qBm9rVC9ooVi7r9ADF3pGqaBSHat3adCWyEgQ+jExPatNS
ejaOtOOeQ6dvkHqyNFMYFgUq8QLDf4jLzMRk9c4jMPDTCoK4LVwe2vH4H4hEZlizJg1DOA7bTAMk
BEFSuZB9x6Rg2kg9dAZ7GBJNqrNuMpT666FTbrqwsxNsoihhrQxNaR3lcPfoCGYmDsjdFsrjScNX
RfG3vpT/gQ/FazZwa1rCO4LL7e69D8BimAu2nA748NKND78h5dhGFzEm0DUUFr2VNVoEYgq1z9rv
JtdflU3yWinHadY7pMuw5aYs0uhiikr4MosFI3v1hMZYC+cnR47X1k5ZNyU9u7XhS1FLK0Nh0n94
/n5xEB/dBGj8RsHQkeVOSBkNFvT/HIgxINz8wPYsMKJKSHz6sAmILpJ0Eo38fZdzipa6MDXX3Cpv
Ec3NBM9bJIR0JuuOWodutaxd/dZ28Ahr5wsJ5EQ+f2qaoqBmgWRFm0llteIc3CvumXQXCpBXYhHR
BJxqypUOHgbSCttGj97AUKjeKSFfLcphvcnOZkG834JfKyZMVwDCY5sBpaLILXbnieT6ONL7Ex2E
9+8SVnKVCiW2yhii3XoDyWTkLLaWuxmWOdjzRxoo/wxXeOMxyG6hNLccOMlBcGEwVXC5grXyHAY3
T5XOMy9bVl68HY0uCfbtC5UDsR4IwzNB64S2Z8QgRqF7l96a7sW8F/W4mXAzvOvhczmv621wSL+e
7P9BJwYGsOQ3AYJ8tmkJHOOcT08Djx6QyoWX3wCMQOuXW4Ut9V0UC5Pt2HsFZRmydoZsldHGZV71
vg08LDHpaY7xWfWDnM2FYMZCHbpi+1GL6XDoy6K3HRkbloHHXykG7Tek96X9IYsD8jFvM8Mie8qE
e7XZxs16H+Nqy2gUrTaI6h6vhoQvvqQRKGSq+44kmE5K/Ehf7p4pFykm9PBogcYN00WP85yNec3C
Y3o6s0lANN3OvkVIrr3M6GqKQ0WDyQe06w2WJnYCixb9I1YVAl9DFWQXMCvYsmmqFczuyGbAwyCM
79pe50byns9fQrNqj+pg3qlTuhcx78TKcHZrAs4FQflseGJiO5N+7sHn+8h2MRlNWafm4+WLjnOo
egewhOoFS6EnmPhl+5XGiSBh9UQtKgQ1wo1wTHK9zk/CoPZX+rFUNttROVYcxIZEy70WvLVSQ5Io
dVHx+JZJlht7G0Cyi/XjM+giiykNP3tiR+4Tdm6imgz0XKsZLh07K/Ssy+UnnzBJhEJ+9WPHfODg
JgIwJRmXYfWXPTsNbEbV3FR0taSwvBzBApkriF7oTt2A8J+faYSH6deSarqIGuQ1SEb9YVxJKAfg
F1MY7x+nt/+1L9e7i8Wxvel4KdW5RlKzp3sb6b66BbboPpzzYNQrHZcFujzVfTtNsrL8zWORAPnk
bs8wy7tkSPqdyNJAbvWZsYCo0ac3RkhqLciM/k6n3JiOJDSxKbZINpusqLmvXlMqj0K7MpBeERvN
05isVrqAlPtJnS/6sgjgRMw5wU50yCLWNX/O6hXu63vPNhSKY7/f9gARgDYPI6V9Z2A0qO6pA0nl
MzYktbv78l9b+x0ZmKzkX3e8+HlHloEQaXxWoVtAAQAGj/yOQsJQ2WL55OLfCi1dpyhkmbbhs2lD
9Vgmavu8kKSCKXZjLcJghGQCHmrvBct6OjFzRyvBKfKROb7d4UT9FKaq4051KSDxoqchaUbxA/YY
mrn31AUYfYQYO+BTHKM4yN6GujKfg9Q7JteOna+WD16RY0cYkq6WJJlBYyYzjf/C63B2pnAE7wsO
ADHEYPWV771hcp57g4fidiZ5vxP1qFBRwliHrH0MtRodDiOZuSoypyaN1PMHvvlX5Xl8VyTAp5U4
0iPVqs+zIOUKqA5Zfsp65rHjWiqPY9hKPnH3TcqVXkgXgxbUuF7oYWvsU/R3WK4u3uK1EpyOIxWA
rhtqht2RhrBLiAqe6L9QcWNHBxuEwoQ0aBsdomtiXYJcUBmC9QAmSs3w0+b5CxftB68QTt1Y4ZME
yhLek27e4evsoP8bN/999RsPfyp1EUNyaZbgKWkRDlkLIX6A7OdomAdRxqoOMqvzkdP5xhDr7GO4
Tf0ZMN4KYjymLm587ecm7w3Jh66WFYMiSc0TaOlGVin86tmzU/cQhNqgM6jYeZXKxRgGe9kyw1KE
5j0RPyE4ehVf4Z94SlAcqmMi/79yP5qpayPcQPXFkvjM6MjCW9fMm6m9JYRRTDFqGBvmlTNpYSpE
luAzxcEWB4MVzQskua3orHclIv+y9SvfEd4oNI2wo1/sSwdmRhh60er9As4aBnA9ZqktJv28HlHj
ZmbwGNgpXiD7yY18RL/wFinZdnlR2L7OzGNfqwvXjAoAzpu2X+g92VnRdddHZPRFpANsNduUu4bA
T4rbqC05tLGfhUWE/z2PEMbLtmXor5f8+VjbMrJ+q8DymLcc1dGLZlBcCbT5dvIi62YMIjgHi6Id
wZFS+Yg2Hvuq5hzErtpEwSXYxVR9GuJpujVoPYLqTmFN4YlyFjoZZxXtZD4iBXRx7Z1nSpsCOvrY
CSXtU1Q2p5zrrrp72zGbQHBotA9uleNVjRpUdLgbEDLKy+VqPJ/aAZzsCaT7oCEDSnR8IRcaksQ5
3g8cM2GDiow+e83FtioT8mQnx/AgnCNo3DlPao3SJQhjjzdpU9Lqfw7i9SyBYDIw08ncMq3ItE6H
M8ZfnUhtUHn7zgTicyoWoCVMZqR88IycJOkZNOzMW4CK0dsN7a7k+oWc8LtnBXcvBx9S8YLTY40V
PK03W9gkMXj/U6iPnpEU6MoVz//PiE+tU3x9Oe/9vtP6x2Y09r1hkobp76K7kQwKyouX21i6LwMH
QskMdssDQzJc03gXKDvzIfr1/PgGRYAIoc93OcyzrJk45GUp8MYsgskEnogERo5K//H8IsQN1AeS
TIbOQKdIIzjSORz5r4/4aG6N5Fp62rbhob0XA5sObMQQni3CI54yhHeqViw0D37+G1hnNKmf3XWD
fpp5ShrC4Y17y0liZIHV8LNKWBE75CMJ2lZfT1fJULOfq4pRqUfeL/kkUkCXw3BAqySJ63GzYyUk
5YLV8MVQqmh8CD2r66dmuevBT5JZnXGxgMToGXnzLs266f2jIxehxPonYNU4EWQ6hLR5Rhov6+Sg
qG9ApTckqLdL6B3h7gOg4jRsefi4e/tPXnc9CDAfXVmsPPHGM5jLEz0KXIytgwndmBjJvCTuah96
0iFbDVLcOSoHeaEzOnJT+Xb6bdsM0/tWKFHDLt07mrY0m8RSkua6vcAx3Lu8AFAe503XZTqa94PK
rn3/PfPaXY7A7Av9Ldl9Yz+CRFNonidaHfd2kxFzwB7OQIiWfz37e/8WknzSrZUi4F/9gwBniVCL
IdfBtoO+N6w3S99dk6unbxi11b856MeuN5zZ3n90qLnr1z8OeI5XqjlimM7aGDIZAkFnJRpKkBBQ
NO2+zZkF4Nw7S2dcSVtF8dihSgiyF5zuKkIhym/Qbv9sD5h/me8JdHP+gVGsTz6fOJ09nMwF4fsd
HnNlO1ZR/FB1PQpan8nKFU6ybh8FKYChR0fwW7l4wbGFLtsxqWnRXMwnrsAXBCqgAK+HIgxZ5wNM
Cy0fH9r5HS3TLomQB9SBfD2iwOeBWa1Yyg/l6nz0FRb7D91RtNe3aTtw4ckJrKT/xJF7jvAdZbEv
wTQkZvxjwLPB9v+WeSBEcXIZwPD8E7dwMGx/V0nGek7A1FT0TI1htriFuHQq/vORuYJPSinja0FK
y5ow5wppNQ33EV8sR3Ez2iCre2TdRnhkb+TA/CdKHqO825B264IhuU+IcHFd0COca6QsXvLRNWnR
V0prA9Wq/ok6bM7n9Zlg4BIq2VsXwVqsSvTmikNjFCwnsecCx1U/ls/Ro9H+b3masj8EDexxHTuL
DN2HFtLWD5MLFPBHuCSWuKLIqXqQQSSq5hwmv0D8pba/CPf8+WG/RlaSfIoVh+FqONHtjc6keUta
r74tRZOHkR284fviLMWAMZiTpiYgOMfIVJmw+mQ3rw4VTw723TUDyMtDOzH9GcZV5BMxJxfOBs4E
9cpNqC5kRg3PeE3qt2Avh26p7sqKp1VWA8B4BBHqDb+EOdD6Ia11buexrX5zSpxV9FBo+SOQ1Vtp
PmqTzD1LQ8QK2Y2ubitfrdF/ldCagMQoMUDCZH++qAxsJYXvLU9alhIGA22Wo15r0af46M0OaCmU
7eru8Vehr03vrOU8Lv1Fb4sNZp6nM0lSXirx2imuMAmNC4XjPTke13Lr61nHsc9hbDaOmZmkIFyJ
OLiM3nsZkPO428kHIP88bsClqZQMyPLqMgcYL/1uV85VaSLJKIk2fYrHETXp9u3r6RqhMTzGdtNs
nqZBwXhjanjZPP1MzSkWpj0GHhx+HqJWtksHtL/PvyJmfAFztOC4Pr8QQRS5heA6jDmUhSPWaTZY
s7+oMcXVuRoilxMrxozmjTpM68XbNEkCmxz8+tm8z2gxHpOs2Jjhu6mf61imZ6IJ0xqirOqvtEUz
hSLqNBdY4kmMJmHRNEuKjZ1mJllSe5SYph3O5rFdX02TskKmsnJsjIKvQgO0VNq1O2kDW1fraIK3
aWksfOcO1GOADvCZauclEUsWB10XV/sP5zGiscaHRNSRZWqnFbv1qnIqm0I822FEjftLrhOjCDSA
nevDPFDhALCmLD3PHr4LpeSKzC8HeduxEFcHnf+j0zzQe82wxuh4G3Bca+XOapQ8H/PLx9iBGvmb
gjDAd7ukHngRGDIL4A2oFSVnkPStt8N/GTM+2A+a2fbvcx90WCzgwHWGozmZdxx39Kc6OTHQ/Chp
dZELyKlVTQJtelxwcsDKBAKhUwub8SI8WNz0R9KuMMv8G2NVvGvCuONM2U9lQpgO+bazqh6kKD/6
RQBPFu/36Mxi/4ARbcOL2NC6tpgRcscSC4MswEb3IwpEvIH4H5mhI7Mk9V+oHFi6otTeZrs4R05Z
WII+jphf7YY3opHAkwq9jUpKJf3CUhOH5wt+riwOZ7JUixnQ1iPMcZYFumWBD5NgcdPtJScuuBS0
m6/F4aCdlLq5k7USUXKaN8NV1oGIZ0mZVrTTIUnj78AtCdl4sO+6LKe5RfiNwdW0o82DDBQYyGl7
SgDACEy2ixQoc8HJl+Qb/RRE6PgAk/b9LQ2qPlx9ua/GrDRGLFsOJndhURUh5aNiBloOYlzYZnAd
IvtIyUr6mJdtEJGLaeJo957fbrsyTGTktxhWxBZoSrlbMXXfyJoQ4yOUJb+nbIEjOUqP2CHSKD+3
BB4MV9ZoonkDO//UHxtbdgLBku+KSFVqwBdm/ZGEjLKx4fL9qmZkRAi+J/EsnmsoUxo3jX5WOP+k
n/kykC32ixnM5EGem8aw59BYm2LBmqNhOBcS/3LE1FXwjryBiMyeZk14+Xz0A9QrDCtaEgoQ4fwb
IvaVWAx3zgHuEHSJcKuyzgPnR/c5xhDOUqGX9efgOGXzgyKab7KD5dZBFT7KvXH9NsyYKci9QpWr
UTS1ODDOfLZyF4kXD17M4Ixv2S3Ft2ZERZLiYXv+mPFGs3oKQnJDS5iK8kIM6ZO+u/VDgpjXb9Hp
iEkCtAvW9vnxOo4mdPqy4Puyb63u2Y801afF7/NqrF5xE0ziOciUEoUfl438Kga4kc5J3r+iGLVM
7mNnxLJfsYOCcfPwhTTfnXaJgxALCL8+09UscwIqK3U8mfj+ChCZ9ztNlbvUU4wh07+kPbM5dYo7
kbdi59XEaMawyMwSmw0k9HFrjf2mzgL5HY3nTtgkth7UYY0K7qEYlstGuSWpVJLzox8PRg+i3PwS
pNwVynIHPsAmdAiPsqUtHLA2ARufD9gxVTbFap4J+kzpwt1OTM6ye+/RM13WmFW4urBrHd1pjOGj
RlJZnlIM5TK06FTWnhB0xBSBmdjGygYBO80G666gkGFgiW7QF3qXoaUSOhycDLOii7lhNSIkbPQ4
FuM0+Uhj5WBDi4bYG6uhb40/3R0Y2onUwUfslmVvPQAb5aitz4JnU0XpYP27suOhnPmgOq4ATu4l
bqdk2sKCfwRHlItq8tCaGC8rVHR0bTG4YYwCfj0+QRY44fxY8eCD6uJgu02vlPyoalJ80kAKYSfE
4FqWPgHd/45j8RUwjgb6rnjzRtPlohvklNFZKwVz6y7XLvR6RQgfkreO9RFssGukEGD4hgTlJ/Sw
0dvfkPb0JAKwtdjbUOxaxnwCVnCwwFBLz1ameSbZQVBmUyjaE6S9BQBhWWDJpwO48PpwetpN35M4
SV3VSQcnu85XmMk0nye+sKakArk10lyZk3BvPIgcEVj3Pn05FVoj+5L1f5ptcO7BpI+IGRxRQNTT
1T0UFRpoAhHzYo82Yg4PvSbVEg77GMCEzcUbGagPVjGxt5mC4tVT7xjz82jYq9SCUfz4PHf/fIfQ
BIDfm0zAXLap9pGct9g4WE8g6O28iDK/urh03SFqRwxGAegPNZPt2LhovYihmNJ/f1FLFS8+5RKK
5SRmkecDYocrTAs+rCYGyKWmYdfl10ORiBE1hUYvEMwZUPdw2ahBSLSzLcmCnIHwxiF+sXvoTOvE
3kOpos9SzKlhszIKr4M6ReLKSNAP/b5RNFNH/xWmfMinuzQHb7PfWFbfyoqbelylaZV07egG9F8/
qMw+vUNzGKRNMpdBRFPwuD+M+wF9z32iaf34ll9CLgXKBCGfLAHZ5cn0PPi31uPH+v3+dyW26OuA
9VSQ6XLA2Q9rkPvm3rICAYUJZdSTHO4488FgiH8ZteUiBhMqNChgfy1Iut4E6yCr4jAHpUgHHGgJ
e/q5VjsGrRciGhYAp8iJvev5ph2P0d5MOqQdpiw08t0ynjAeC9TVmj+AnPAxzkEjN30rRmRNPprB
6BUsgN0a1bY6xHfc9x4hEoYOftUcnw0Yyc4OPJkeXDs9NlymxZ83ZKOt5uDjn6O94curlYNfDdoT
AXU8mdBP0rlcN8ckFBJZQVxgyhwS0j5Q5AOKh1hvwNhkPq7DTR+hml/aNNhlO1hgEhhxCZXPwY5E
EmUOd+bIT2FjtJJ/qlqvA6G/uQU7wlHG227SN91MyV/FZ61hZVu7CahVU6WC+aet/FwPmbsH0MKX
geLf2f4m8HEknkt5ZGZztSpA/Mwzo89PFVThmYuQhsZgzwcrO2FfgSJ/aTwgAVc2E9mzK5HTfLGT
sGSqLaS4E3mcYcl0V0QsCHrf2+JzWVAm4O2AzwZtvV0uAX8EyOTAck6PF1m4yJYg617nENpvzVbl
WbGAzgBgrcKl5TKBqg0p5l9hq7F4Hf7Z36r5LW5LUvbR0OLSowOre5OsNwCVx9xatLQPnjLIfhxb
LdAR/ayChqeGy38yI6OD43d7ksRDK6xiQkn0sBkHS0lfNwXM+Ei488Zwr5e+V/yz308qzHbodTka
oKNdx2L21nainNxu+SmlwfbwzPWNci726nwK33cJDdDXw8wwkBFWa9sMlItw+z05nu5S9gZaaBK9
IvcfdZA/d1eM5Pqfx+q+Grin1se6MDsgW8Po8+goaldL/fnUjPekmShQ5cqCXEMgjTUUx1GQc4JL
m7qE2bAgEa2hZW/821jXmMrYwBevpVL+cL7q79+/VQRW0+2A5adul/VusSbVQdBifB1CS4PvRJ+v
VP5B3CbaXgxXyUO9L6xvLGETdWMC7M7d7WGowGinPz8lVSMNiXGi6LzAyNAGmY5DkeqX1hJFI5dS
bd6GhlVS3sORc63Ylwjiw91IURPfSZMdCPEO3wFo9o4ziOBjGDBpIJNRFK5mKDnpQGR8GNQ3Yygy
XtfdI0X9iUjm8tPChqJicdt/4Gvr0Btg1cWMDyxyaFZu07cPgbZXOkDquc+bW2XKQot40wPBWenu
ilb5RXW1FyqPgIFjuYPz1pL9QbiC+lNKSaLZL62ECQ9GCy7h3Kso62DVNE4Pri3T8pdnLg5uMSNi
BhvcAdSuM1K7XpgPXrOECxvn68um39F28l46/FcL+s97igy64FzRziqXFE6W2APUKqQuz1A4JTKc
fyX54vG9su5NLeFSMGP82wCW9Eqi+BssCbke12dRlOmxrFbvAnfYfMlzHwASL3mxWZJV7t3gOWJB
bA7+o37OGMznQBSxicZXR3xBPGnbhN0sEl0g4bAGvD1Fgqz//qr1tvdmRBlAhJWpq7MLUjiCQmK0
F/YGKUXyA6gMMcDmuuaHk8uqF5jAyXlGhq6RA6nxmArqEIKm4CXc6RiSjq/W+LsDQCreG2m1+FUL
0Odrw7aEZ+gsewsuQ/FX/Kg2LA2LYwehcDn/VHCSsdzUwZm+5rlygVyXlPxVbghRGz2DAQGCShuj
xmSO5IqEJGz/rHdvBTF4Ee8ZPmIamxQ9kdioiLQOnbk1qW7NbEQZq1L8onoNPyZ6bdkniy7kBsTN
LtaXurmke/YgWCN/lfBLZKf4jqj6IZWevDU7K10LF+th4UvJ5F0PJ1THFhSwRmPvvSTA7Vy3J6f3
WSIX93umJAHC2vg5ZzJ8Al9SH798LRcdKBaHdNtxsr6l/kui9UbQHHXWBkCckHh9hyQBhFpeXCoV
lR4YdwjTmdHnt8SNw6kPgT+A04S7Rxtl1WGK1nU/lnwjc4vzLIu1mqgtxZQ+Rz3n9mJECqFJqAqX
tmN0RM7yxvXfwk0qYFvcUV8dxU0w0FGfybQiF3uiFQjknX0faG+LII/UYQX6WvrrrQxO5YCk0rrl
0tWlNtkA4S5VEUwwk2u6QVcftvGyzOctT70Y9A0Y2sMrpPYu3Oxw7XTTBu17INCL0HGeCoaXXL9b
I0jnfFVoW1PUlm7c78TZ/AyAI3KTMBJICh2iaV172xDGP/Vu4nRkQAqBIcSg/35Kf9ouNwde+vrG
cUJWhVKaqpj+MgibNX3TJpfujNoEH8sXVwl6LTv9AIktw3jwQpVXYRUgkAtas/UlTCdU0HeP9HvD
ncwEA18NBT0os0PiPrLrvBOqZ51JK31V872Qbfsr9tznjkVnetdj90l+J7eb6G4vC0PuOYp4B3PW
qtg/WyndQQXVIyzoJVh4VddyXcb1/906wonM2ZIWvTkfn+ZoGKPwBZG2Xy7EAhWTLXnP5qDd4LjY
82CXNBi9vp1B+Fdo5o81X5mOduuBE3mpVcSzNDhd1GoN8Qmdhgp79Mpwitt4FMA+5LERSK5bGx2S
yedUzoiInOBVn8BED+HeFk1Sn0oVD6A6IZzyKWmbgj3aDufg0PtNxm61j4VakCLILf1ImdOeRWD9
geX2C0WWRFBpRJiv29pxhNqjegorKhHdKbw/9EHca5ufAGco9GrUkBx5N/aMTz/17JFF/mrxAWHD
0qlRG5lLivdaAhQhDexj3OeOkspZi+fycZ724wl30KQExYsRnybZlnjC9tab7BFz+Axdkk3mSbAd
9rBRoJ5Y/Iew4bwgHLV/AwaMg2LXhcZhtUxLeObLEBXrfsQ9CyLi5x8xSnHjS4QNI+l5vXO3b/fX
v5EEvOyc8ZV77Nigf50wjstRsHRcQQ5ntBFxLFr3ci/513+nBCiiBjb5ZbKJvFtBZ6tQGkgvAKjO
gifcDcfuO9opnKKAZN+lW6CrQkw6gB7EOId35CI/IDqgLxInyZ7I7WZATAy+rGJ1HVLOpKKp5VcY
6cV6AbhqMPgm4xProaMPrVaxLGLnRJPyVvK7Zj6ni61x9sXO9juJRjnh1sui9KjrDOyVmRa5TJ/9
Bg5OSx3GFmQBBxb3a3fQb5LFLAdESP1+MmJ7WVEjQF16LE8Z2Uxsv2wbw/7R/BQtgYt7u0Lu17xZ
Xl0VwAubOvN7KGawZ5v5Waa2JrkuITV44WQ70t7NUubnZjEh6pC2yoGWIn/lW7VdkrKDQfGdrkZR
STQ3Nuh7qMiMxB4MT3KKyaDUpPF3eTa0IfdQdzEILFboya+ZkmxC79BADyUdexsz4R4HHlBWIae4
HNWRXTxdSf4JKZgAP6tI7xuqLo+BlUhwWFyyaIqeVPdSK8u+6b2/ZZp+I4ffAokbYFX2f6g0O6Td
4arELEO9cx1HsXO41sw1hPpHqZGIC+jDOYmowZEW/fjruWivZV++Mrdx540HOvLyq+/FfwWgTfmn
SngBpF3J1KnkaXGBuivZj/gw0hU7nfacOIog2s2g0+65pd8De3Sb/AzdelWHupcGVa8G4uryMds3
OlGV5/Ya/dsSTbcnH9hDiTzh85/tBniaQyuxG6F2c1cmF35/N8YojG/SOpbQGYJacxD2420H8HVz
LY5eja/oo91JEF0+8BraBpNIVUbFRAV1ZkN/3vb0R73HaalU2Y29fRJHjVz6102ydXcLrzfCSGvo
7ZHwvEoLQuR9pv1zmNKT0MkmvVw9byFUcw6iXMLv2KAt/w4SFa3CO4To9q72/cnmhGpoqs9P64h9
Xqpckd/3fGwztJ99lZXMfHG9rH8iWlClW/rB028NmKMysMAwqLv8qWmJ4MCTdRDy5WPNZ7kdXrPn
LgsjMA5kDb/HQGV7+cphpKYm0KqEPLEsfw1bGbD1m3rwvfC4IrqM7wWUYKE2xnobRo665GPvAGBr
NoBGUXLwE6OoaHcUS9sZ6OWRtw6gL6ynIR5pn2ja1JUQGQ8tcUIBGMbXijgH9vnkcljvYwS7Z1A2
hxBE44KV+clqxFrM33WWv8gy07/gbjOMJdXROW1rbA62Rl0TJ+P+XFAQgV5h5LoK262U3VNpoept
qwoOvXJg4jWcKbZeNLVZbjS1mTLRqgqXsbqtVhGIYd0dcUIgbpL+PPfd7EWPSfDLlGBCHFfQRRfK
wtQgyh2hiuhUtbSOU7q67kC3A7m9cA5wCL0l1TDA5+/wzgNaSla80sN4KHKCPVSGprd2AQUz41wy
qS2dTMpJwpVa+jahRRaxoqTn0om1XFjNqmqY0oa8c3U8cs/rg5HwQsTqR6V/9PZElW3s0175V1pZ
F3qmgyB6QM1eUe2ImIScfpyncgB0jhGJlRsOKFQPsu7ii5M0gog7bUueoQTa9YiMU4BajqteReln
vE2nVBhhXh/hgciE/8Z6a6GdMEMP90RoloDkBuCJIo3wzPbDkS9/xllBAynU4A5K0ydo7L8ENtja
EdLey9EHWCVuVlT0Fc76YNkkjjG2huL3K/2iKu0yGz/UGwbPqPaa1e/1koeHD4ZZB5bKA9s4Gb3b
l6wM57aDuNXJqQb6zf/2xFnUMdGec2rw9p5Gz0wXHbrceDhZBO0DZx8IgzMtVt0yX++ZPLqI6ua6
/t1DiAA79B8L+2KcMFolw0MhEPv1oY7qM0x3lC3YHcJMcccPmErpgOletuFdWcCBL12eLRLGDYCh
88kG94gD/MH58SFIoX1lcFdKUhmUIayBnWmu4sL19+avFi77bpcgE9eWPPavohTSGJn9hlbH6sy/
V4I9AykWTaJpBbfLXlffE94sCaFnNHFYtQpG00DWSFWeot0z9QZc+rpKAnrRr3l8P99FbQwKPkJh
GBU/5NR2gcD76W8BhKNkH7PIPe0CUGX5h9StlJNcrCvBAyeyPvbhl7Hy5ozOzw6d0tzQEMr+Er2I
dDgFkhBpM3QHN7skr/pUQkdM5cmjaHnOsj97FcoIMLs60owp9nBrsddM49OqKtaIzSRsXawv9aze
QRV4KU0mHQZW5clcx74z5171s++LN54nXlz3/gjs9NCq5N0lB0+Wh3GHIMI29djhVerXPopwjjBI
g8Yqmr0zwo1j/N33qm5ojO14LRlEQ3/D0hguOPtKja/HJdlSAw15RjkGRaigNPb/7+djBYtbLapI
YbgcofutuD3oD++xeCtR6cRJ+r6fN3VnuXyMfUPNsXxhDAsgdrvKEFpqbwd058tbtJGtU4A7jths
7eEyGgAVDNNq4f9xFC67nYrsC2R+MSdYtB/UVN2vxFjhJ1tzw/Z7mm1z36Nh4zvM98ck0riRUDsJ
s0AMQbZT0U/UtOO56Bz78BrF64DdE/AcmoFfIoOoebwy/c/eIdvG/drcO3Y79GHd0AUgPoJ8RY1E
WxlFH8N7BT4utvAJ9+3pYzPyZc4NzZke+Rp5xo4gtHVOVWL/gQN+3IhBy1vrwuh+iCDIRX34ZBqs
C+5Bwy/sy/gJGvde5ZkU+5BTBiO7Ex8DkNdSCdb3xHJE340X3wqdoGSdipm4WjTOQeV+BBlD1PAD
1IHD5m1IiozGD2B2Y1JKnwGwQbO++07rc/WuDkhoYtNCObLY5ZjkGSoleEZot803h7IKGangM9K0
H2dcF0BiGMacKoT2TdrPAxwqH3L+NhaPN0ounZJcFI71Z3jfBgvDEsQrWaho3gw425f6fXcnFMhd
kZ8v77VfytBFmg62FF8nG3KMkHoU/z/QOJlpRBu/YNtDCTAi5dUX4pQ9Il8ReWfIJbMqt6lidV1L
A4gW0TKcYAcHhA7uy5AhRNzTQd8RDmRksQiQuglyKcm58ODTFt4mzslRflj2SNU4XT3lNRwR9GrB
H94cFbBMEkpeQ95xNAAKqsJCEt/uYfaPy6FoSQxuXSe9egjUyk3EnK0pMi55rXWPKB4F+Rr4vz0V
cARn7bIsBjsVePmVMluaxeaMRvMwqx+A2dOjGalfwgcGCRAUEV6Wus4TgF/qllX9b4IaK452QfbV
GOFshmxhofsnB1tJYDNpEGYoCLAjyxuTpdVDLaYhsyomsOGZJ+IVR9LqxLtawSkWfTqzJec0v9Po
bHU6odSz/C1RM7VVjfWZ4fBmrW22nhp35VVZXZqUIdYYaQQtcK5IG7U7ATFSbjXIdLewtaybvQO7
L2rednElDgOV3bt4PfTD+oJItEffzEezQmik9T4HpetX3TAHaAKw3ltLBZWmqp9uaYkX44iTpsQa
yHEGLEK+Fe+7xJI+jTe2Df87kB088D2wMib+CYjbnXsHuLtIFF9HZf+BHzikXnXZCPQSn+cGvPX5
WvsDhqYTZgy65PTLRsXXoKqB9JQHTOn1jxO0+KsRGR9wemp69XCOTbodx5AqhcoY8DlXuawnD39A
Iij3rZ/rhHIlV8u0ZDAjp4H/DZ2PuL4er/SawJd8EFQ56hX14lFz5paCWJmYrzGI39F4LaNdjPXM
U+/su+sbJ7KKmgf/i9IclxCaw1KVwH8tpuwnex6U5jEzOHbOXiNqAt20ptC8nvkO+rKpcbwCbWg+
0Nqc2J/X8EOngq6SK2iYTicjqNgLTAKXmLAHU2vhNjqb+bKBp1HS2+wY/NS/3oWFFtaDLoQOW3AW
eKQyYC/D3mGZCFXLWNiP7rRxp48n5stINzy4EMY/e4AOpXFurnun/qBKzmMbpOs3CZb1eCgCHGVG
2I3mGhBAXrHyn5w2da/OpAy6kSQpBlb+tqH1sGjzBYS/516gC9vWx/fw5QvsR6RfhQTCFYxCXxYq
OBmjhA4Gh41vu3mcpUaQlVQwpFk5b/28Ls203VHy5MstrgDhxClCpAmQiWYE0N3C3maIgufFqjku
7PRF/8N61rtrtFIVmDXdcNeJHlqjHTOo4hTZ8LwVltibGr/l1K9mkS+n7c3zNelyk9ZNwC1ELfvK
jPHz+CIuAMNvk2t2RqvmzYePdlsHiE+ofDhyq5rGfN8dPMUBGa7gPCcMsjJfyetteU7owJaT+al/
Wj0Grwc0wLv4OQun3lUT5wuipwwy5sc/s5uXHMmbH4YUnoxSdC9VW7Xl5pGy1zLGHqmsdQFkL8yA
rPEiiotOLD4O29Hl1j0uoOYEkY0sdSM7pdZIPDIH0XxU2aEAnfNt32M7iviACzFA6/T7S2flvnCt
Ti5wBN41Wj4fkoyt8t21BcIvbra8jV0b+KomJfKXyW4HCh43/sXv+wAD8yFwwEWC5/DNoaVKfFsl
DMASdD6ycZEjVmMx8PZBFw6jozDQjgjc3/Dx8J61Oss9sDMcI9GYpD0BvhAFT2H74O+LOLIKKfAp
TpLCLPJVSvJiopoPX7U8zeQVjAomPlVwBb7nxJNSlIueupr/FfPPa5X9wPwYgw8v8HLGfz9Xrphp
uzM4jcaurbaIiFxh4StsJB0iE1KacH+1qRDznsl6pHmxADhIhidCzHVLMPUbAGhlOK+e90WCh8tV
XWLjmhWu7ktgLzaCM1enrO4jD0Fgfj6cqw0UJrho/9prQTpnWnOJ8n1ntYRozmCbWKyuKUmTBpxN
VDpU9jJa9GyE2MSpEQT0sck16v1kjxSwAUvOk8mOW3AZWvHmuM3/EXx10khiRwB+z3MFGWJSYyE1
UJbqPvZprm+HBd0o7z0iGZCjx3eQcbHv/nKfDQTCdv0IKQERndC3cwT7mBSdUCvAVG9zSMdoNFTc
MN9JGp4fAh/QGYUOIeZmH8j3gUTowsFBtjkbYorWWglY4torNr+Zj+Nqz++7coGQqHb4DiW7iABS
QiUPp0JwGx/krcGj5qZxBhfVtoc7p7OOVQ8vRohi29yncaFHU4Y7Eqq7erbLUdjg9FHZg2bTTVW3
9H3ANh7M4w0qD/H/LMClEGVJJxaqbxDlBAo96zv2Ow3cw990epy/FikzqZW/deoOaTuEVU2pgFIZ
eyTAq8NqZMhlRb43TXO9ALXwf00pWsYjXCg9vIVhrYG03G8HL+T9RhF8DsmNYHdcn/4NYzwYTgYe
Q9qeS6EyGuehxcK4iYPOS5YknSd71upFtNEZ6pGMD8oYBEbkzybJnthts8WYp/dOLwi/11rj6eWi
q4pTPjCirM+o/YSlKQBg2xWIxSEKl0flJavBVmBMoG3euM087muB+Wqk1TTYSsBurzFG9Frp4GU+
itNUi7ybty6IOzmmxUG2qSHbCh0GZ9ie659OVT3RqAk/Y0X3y0IMubk/Xi7hkG/keZyFu5K7PIMt
upGgcQHqjEtx5sKcRmkNQqIkbCxpir3V3H0KULHLxfj9p1pCAmmRnwlMA89v0WbvqqUN/5qoJ9ZU
ViIfASw5KAxfyFUhQUi4XMDkKlqWmZtDfpg3uzkoe+6ODnI1onAHN3z44D/z/GqsFLwNj8+I/iW0
MDqmr5HbXns/CdeMJKHM1fOY8kT5QEYcIdZCIBZcA/hOBvRYESru/RGRd5padZklgE/i25lYbClD
U6R9rD4bPcS6UB6l10K8rsGfkPdx55fnWipNBlzxl1IJ1MBfsB26X7wWUHlKinQBsjP9H4qJhcp0
j7r2va3ukicnIkeTw7bBQ/2Vyu7tR2Ms4oqTpQ5sKFVO6R9UwMhycNXn3t++O17zSH0wyT29RXwe
mN3gD2N34jO87aP7OIzgJU+AtY4EUlyqQv4AkLp4ijSb8++2fwHITSv8pRkgzyzwO5DFTEP4skiH
JxqIli2CSp/Bpc0OYDw+995AZvygNkkOe+pPXOhNH+scLVuH3aJU6Dq21RqHkFp5thFGDNC775Ie
IcPOb3tAgnwrw+MpKlx9cHhgxMl5C3qMgwoIfxUvWyhcc3esag3FyKnNsbW1murZJUFY9Dejb3bZ
26B046z5MV7SuvNYuFr+S6XGNu6YCxKmf/w4AkGf2vqWMskrskrJQWZCItFfe8VZfxqBnV1gwZ9V
4rXN1zQmqRuS4yGCWI3UGaJ1r7CwdK0FQlPKk0WhMkQ0m+LTQoPO6omN/bZHTbQ4dQRS5qu94mYP
S0OjEc/FjnnWPgA1ltM1uzfzOznGrFRJEswCiPaSRTvoOoLMW4wIBGPfdz4k+8o3fvSGlxU+Mxj/
aad3mSf+oUM8CUMXDW7oJ1XQ0Y5kqu9bDnmuexqo9GTHGsHO/py1MDWbBZTgrlBA4ZvT3i/jA9xu
Iyrcis78E/4+yKJ+gNDAembttiz1ZItAoQb0Kmpsh6+wK3tvMbwkLmqnd4fAHapua8JQCZDuQK3C
QybS8eLHZzXoV3lrKU8WJLRGEjcmlc0fz/KA7xyi4aHk3h2GDZC7quCBqb6yZgrap4IiiWprh8xN
kOL9iTbGjWSo8aL6ovj8JiO1j7ptwgH+K5082MFEPxgp8junbA1UKTuij3azwTJGaA69b5xNbZlY
0axsdscyxAAo6SaYeq3O3J9HkG0/YXJiRHfObKBtLHnlg8DA98227DPeEQh86SNQfdtD45ryFPVj
AGgNXXeOfWUWwpg1V+zeL86wALCQryWhCokQ0hx+ixJWgdUuGuhaHnALo1795ic/x0zT0tefiYzk
htxdXAh5eztctoMNJayKbFTydftfN+x/ng74pT+iDPQFgiEs9ED7AzOKcvHS0U8DYAeGg37qvTVQ
PSA5BxwpFbkoHywRKTZu7sFqksKJ9/hxyyT8BBotbhEMQgXDelc8IQScV3lWKOXjqnnJPIawu8nf
NlD9rFH/uV67s/nFWMHfFuFg14TAYPU4P65XwdAXjV4rrQ7G/0/aEWgzpX/YVUpHrjn3VqyW0ze+
GZlCok52xtN9//RQBKFyKxtKi0s4SPOdMwa+ggwE82/hEAQkr4dTy+XBrsFlVu44Dhnb+3WkHcyH
siim75WBxLqq2gqvc6j7hsRyHJkU+8YNqIFI+IssoX9aCvrwSv0+5Qu9n/b6kF+ed0ZI2r2quO2A
afVhxrHGWOTzjqzfnaKfdMiZ6wSUtni8oXRvh+q0BXFwcbRk7keQbfkW2YFZz67xffogQqIGvvqq
EfROp7NKjY0MjYf9GNKSTShJduHUPGjRr4k1bxr5YLLkduCG9wN4DUyfc1hpUx5dbEhWkad999C9
eK/9on/bkm8k77H5rSAEmBYgigZzOQKTQ/XOklFKXKhApuoLE5ImuUjH3Iiyopjpr7vavo4aqqxQ
gRWv98zD8lR9yVyEsnOG3ehz0N+2BTyfyU0eYriZwFqZn1ABb1LeUZ27CVC9MwFXNw/sq+DDLWsU
8Z/Jc63LSA4EUe3bEU3JOs8q6EkixMhMtzwD3eBM0N/jn9li8vrrM1kCvJcABPjCQDKKMWrrgH/S
z/db1ymtP9ul85E37wVEuyLBllBhrWcC9ICROY44ZWynFddEn8PIWvflABRwbsK7u4Ktqmok3iwv
6egWjwhrm+yDCOlGnJGEuqaNjuNBoQtwTRTVXDVgtworoWGSyAIBvLPT1OiyTmjlfD0WHfqEdGRE
didUrFOhuOLAiWAdRO4Rxqi5GlpdTRHp8UVjwfJepAUZOp1zlw811RRqBr8naLFaDS64sCbOcbEm
Hk5VeLcKAwlroz7Kxubu3n9nYxI+RqgCNuXDpPQw54GaOdbkRbyEgla67rV+VExXGvHp//+f/RtC
MmPtI+71VCRbjxWnMOxVqN74vULhDH5pR+jnpS6Zub1CVlMKuTGoPYZblvdJJy3WYBBSWEnvwzaW
eL1exc1bPZiaGIh4ClfKZ7Z4R6/f9D5srNsxqi2cg22pH/HvhpKK/9cp69RRmQOay7jH97/P5tTY
3fQZswzfcX6dzSB8AIY4aYKGlAxud/4+MCuCPqjiqj8nWtV9Pb7pvu2xOZgtFA1frtaTnM5Obbwl
Ye2ToQEjA2yg/esTwPWvVyFz2/H7DxJv2SsPv31ZaTYujOOLoBFCtmKOCchOBwPS+DRoL8j0NWe2
zCcT6YBhVPmFSYDC600QdLWJkyknG5lNfMMDYfaOqd7UkpIQla3gq6+U+Z/aEU7cZc5uU27BWjgE
Slp3hLpkI8qkRTW5CfD+8DohvM4LLSRfKXfG7SQA/a+AI6CubzNlFYBgLfR4f5ua8J7jGpcaIZDy
rgpdyGu3J59qDcdWPlVnPDzM96xL9smb5N4pISGrxcP8YghRIqPmKVCCULWxd8dTfVjpfzW78yg2
lRYTmzCXu5DxwvgdZAFq7SbkkjwtI5vLdvkHgVt1TL9wz8VzxEB1+c3HV5V6yANeYWK1cpIlWVd/
XEUp6qsllXfdJ0WpBzxQEalnt3OLJP7JCRUkeUks8Vr0V5XJ2B+IUjCUY6x+QIYaruhaj27sqzQc
JRjHMPWJmbXYqgZALaZnjo92rb3aM8GqIGd28mMB4EiIuzo2dwymkqw9eYX1M7/kxe2ELlCg/0uM
R0idZssWkzCEVVrMRz5vMh9jQuBZmZx/4hkb/j29On3GF2Q7EhBKJvnRukAoEC0cBKab/79gzDPx
HBNdoni3kiNiOWDThngGJ3eAYYVtO8QLE5OQC2xsUbwcJxYz3xLrpdCo4oSetH0RhX7UdaonZA1i
ZqQ4lLN1Pudi+V5nDqhAHRP9HQBfCT3l1PGcbSBLarkIsvUh06BcU1CNik12ldRGWHGNEt9UCq0d
E2W++WjDcDcvXsOSujxkBNkal781twQTrS/YwNonAow4h1g5ffwJ2lmyfIQW/ItRZHTYeqbliXh8
CXQftoi/dRxMz9QH7vSougCpJzB3YmoDrqdB8Q9ZkZGEb8UHDp97W2gRdHJ6to8OtQRmR0QoL3/e
tVrv4bF8+iZrkP8s5swfMiLFbcni/5das/07/qTNz5084ShbU2DjmRj1hUEk3yOHr21QbTKoWzAW
WAVmAgcYbczV3W+OtOp2CDrnEFQeL7ZmTLG2wXM0aaR3TSio4BDtLAfDx4Uz1JkEnPxhk4pWDSbH
fUDXdZLReG5pp09dwVoLdVvTO6sq16A+ye1wdRdGekuWtt1+IQ1xM+DDohmTi3sRAevkANCShsLo
PgeK3T9/Dp+9Rtb4PYAa3iMGRc4FKOd7BZnrhVlyzDyPyZhOiItfeVJ3VoOopsMx5f02D8Zkauhc
odm5MTwKte4X7YSXlrwywRArfiFtNoTqt/Mf/v8SrsYGenEzIQSpfhRE+xGv8rTNZaEQEIb1HE4F
wPU09whrdcW0OImIIPV78RmePF8F/EXAv7qDwz64yRQipOC69TJ+LHXugZWUf8Btw5d9mwzhBsgF
HnORwZ2Upwt14UVzWvAMiM8iL67mR/Lf37pcXXnAX/qVvTAtWz0fmh1w3ThenlTH1RQtT7DZymq7
jVduMEv7gOcYV2nuDcLCgp/z7M2JC8T8IfsO6FTWJ4znSc952AACjf+EPGtrQnlM7doP25WM2SHi
1PTHNMYs18Vv8fCa+vxtG6S/IO5cyCljp2OQNN/ci+z+v62s90w0t3rrvpcBTCh0CN2irub1QKsl
yQI55kV3pJlhIOqnslkw5xFaafowhbmnpPnTJIq/fHKQUxG+Uy/NmUgC0lW+DV+FEv6nB7atfXqB
aYQYRWZxaK7xzWlv2KPwuW7S0/Rh7VVBYBhjXLSukwn7VYr3ws0iH0WAgqxKgR2Cv+k41rQ2WX1R
rIEPLdsvpbJDZthb61VP0WpVebQv4aZhA9lv1y56UbG6oB/33CIrdfe90qQDwS7yf22C3LgxMnbN
MMekmjyCCu5p9S8q7fGibpIkxMpkG3LwhkVb25GAOuiCV+T6lwkzTK+ltIcLUkvgwBRJnRsMiopE
vndICdX+5qhfKFui//krTHIUjdl8bD6vPJegFpjoHQzEzZvTVAPt+v/CAjMXoUJK5Q1j651XNXhl
pv40cO+4H+SWmCv048t2aTksGf5TYYjYt/0MlwEEyaiTw/FbC9vgex2ebl0KaWf+3FOIhnVcuLwb
v9f1j55XbKv3umuR3VxqdY5HXhkRqnB/4WwqzLI72GxSHb68kIr6WlUu9JaplQDCUNTlkRZrZ761
MDzOiVcTppBSfWWOcppRy4eSHdotCdyK67BoTc5Y1C0P+L4bF/jDh1qP0U9znsqEf08ZKSIvYzVv
nWe9JZeH2jG2F1v21SbUu3XC3gzrcB3t4VxzlAtKZOFJ2creqRjZ5FnqkWv8p+4wT5jiQoc8hulC
mTs5Ny3vzrK9Yd+GZeqYVePaAWB6nk1TsxpdjiNP874GN2hp+8CCKlbYFhtiMol7RZxt7to/llmz
B6ABx9YWyisAYLP6P9Huwco7aRyic3FS/O9+PjXXDrO/u0BfutRulXxEwm/IR+WeFmMWtviIrOkJ
7ErO8ci04AeO03RC6Gt90Ty0I5ZX5u7gHzK3Iv6AQ/zq7J7s3oeJvGiUHP0QK+9EpSv4UnWIWMck
yfh8+SWI10KHcqOsd5KSaKKgfuIEodFHql6lo8E2pRujltbZkdmzgwb+3oWSPQHRkD8g9DqjaNdi
j+/opLB/WU45jH0WTrROoaEqKWW3ueq3D4tZniInenS/VJQFwzRfF07uhhtdnFzWy/vBcbyNM06M
LIKLIYhy+cr8m8GnwPusWdifN8Mjn5LvrtbNmhPYQGn7pFt5wO13O7IGbEwRPcDSVSee/D0D5F+G
ZaN4JcMSyvoOfydi9k05iT3u+vNQ5xj+NB4Lc+1UyBB7thAiwTydld3zrbB7YCKjdZj3Klekg1sn
pdnW2LUs2+DWySVzgxo1LFanWCNRzdA5wuPNXvong4OB79ciYwb92u8P6qxhFJd3nwYQyGKkeaFp
jXM2Kb0NG+SI3In0n428rK07SMEEXPm01FOmILRhWswlZ/T3zWe2SlFUPvus3Lgww6ZggU2xagCH
bQ++NS2cd9/QvIBz0SRwuFnH/j4nkWjKbRKVlOe38uhIxXE2zJizPa7X+i23wDHfG1EYNwlma6w8
eShMbE9vC4guqy6R6CBO0TnwJaxZ7HoUAcoi6xUxETf7OGftpjjMyjQiprQynUrlJhV5RJimzb6D
VVHzedBF3MK3VWbmPcQfgmFPD0GM9E3JaiT9CUmo/XQsWBJOW0I7mAkP9cQ0ivVuyBVk1j4gLoEz
YiT0KhH6hZekbMPJXkkvNSh0CM0WDI1LINptEbt3YPPzNULAJB3LLdgN0/fe0+XVXjda5zCFVjnl
EAtt/XuOr+UQCHxXmDoavxL67LKYSHzqDKRXGR+pg2wPEik3UMNcch/Woit93oZFGwT38kC7dJWs
aEOn6HsOFWa884bl38wqnN4uis+zEDy5Euo4J/Yyrd+GKHrK7t5iL63X8bPsaZRS/YG9gufmK0Sm
ogV5zNEBdDHsnqBFg8OkYKKtXZ039M0lbibl4MMVTvdZjSyABcsDt/Kx6sVK3Rldv9NfaCxI3NTJ
+TgpMl2hMA/tv2nPLvg4xrn6LJKFvO71MwmR9eUNc6bmZGjcgv9t15hMg+w2zFlSyDyHjDuqIBgb
ihO9BBBQBi+dDEn+STGmTe2prMEp9C7SvaNX87SQ3+AT7AjzOiuvavYkoXN8iKNCGppH9oLyBNSI
H20yNU7LjQ8T/wEo4OqkHyZ/t+csCDtkFkiYt+Qu0MwAytfxAtZfFK/WXcqsIAMC0xbAVIwR8qiJ
llg9HdXSWvAc5LhoFXgkzXsMGD21jwk/TkLcZQCuXFq5uWsQ4LXzZPmYDRY8T9mYhEnk4T8zlAd9
xTYDDnVAIFYuh4oWoLWkSgnU0YZu9VHRjzZ06s04nILsgDTQTdzOQxS0mzGMBU/BPbdVtmPZDmRc
qNWUMIzP1yAAGCC+b7E69qDcHtuh3GEH1eubCKADrGb8tKp+W1LosBCDe+rBoUM6qElkavIWEESM
tQF7ZyVoTVzUFW+c2WMquTE1YYRAmH64YOzYUdxFAYP9jqkDciAw0fwuWGEsLRrXU42grKSBzN65
vCmSMv/P3rYV3zKpk+jEsJk0ryo/Q4AUaukHzqFf21rp1CHX5befnLG2U6Ldp/azcLbAz5PQWT7X
BnfSPR++2rSVbQpRx4e2fE3Fbh4aR+WxnZ3tR8vd+IpFQHttDV+7GToxhqqK+baS8ZoOPxpOHnET
wj40HI1AtqvRfd+QtgHQdtMhuM8gP2X68ZInydrI5VQXfad+CZGwM1nqNXH5mNguaa/SzPdo1iwR
Vpz+yxktFBn+ZeHh3XfWhMEaICxWspVWsM4DOmhfjQM0xVZsJm2SjRf8e9xSP0M6tCFbrS5cUoi9
yAr/x6ggNCQHdYqgI06XMiJX3yqg8CT1Goylkz8POiTVcy2B1/HOlJ4anTb2akMV6ZAZsPBY1syz
izX22KVngFtQnyGeULGa23iHOK3y/PUeSkR0mmi5Kr0eK+tNCVMsTPWEdxr+YYLMLNNFUefQtku9
LvgXd8jSuo09KKvzETf5wK3R2bv8KF4PkrtHTmLizgjeWIQqgr0T4U/4ABUliLu2dTAtyhJxiv8b
45POGQ2rwUfknODgVHz8T+84sFCFnUmUX4jeIIbmQhv+zkbwcjT0gkuT/tROrDhfnr+nNiiRmCxX
gwjxOXC6kOLjccZ2ig0CzeMIz9r7rEZOp0Zp/4tjnCmjpRGWIt8UT1ckLomyycIYSLYuZpTHzWDB
yMxsVJG3arj/29Nc4GYDsadileVsq29ikUvldnrkrYLtr+Iswqgrt45+jPEW9SvpIyJxNUIlsv/G
KclIWVpdTYDLzZsfvad7EaJbnA+w2Sfsxs6MBxpkCNPJPpAGO1MPCHLMxi2n8lsJooiH++lSjq2r
X4mdSeo4umliUYsyPsiIQpB3bNCKm2m2tIBtnxyw+pvA+RxSbZPwZZGmPIASfs8Dt3EJZrH4AZYA
ELNyTSc/QWkhI4p+ZtBUUDC5egrZCx8tLyCWV9Zus5wtD2gTMM9fjiXaRUy34mkljxLp4P7YYrFZ
s/z1d0HMcCfi91b/L3J29aTqPV17qCnhoWJJxIvAwXyNMjUU0F/SnZWHaFs3QBrHMiVsIjjnd3Ug
JM1lS08e1lNfPV38xxJfFqgjoBU23kquBu0WsbtYQgBqKaKSFSwDDStm9LXZuYLgZxuOjhr9aBz+
EIB15NqJHB2nMTWz9CEwtQYhqsrBF46SF4OTSC3VXSNL3tC8gPu91Pir+7GMieuiFVO29y1Q848J
JNXDcpAoOh6M122zVuP6aCes15K5f6UlBfJPF1OKhIrbUKKyraWjRxD1CLN1M0NkcY9zX5G/V/Es
sVBhoQpiMX0dao/fXfCi/W9o0Qmitp+lB8KoQN913Bkm+dzmqZ7u8+PklWmA/JhMMAsE83JxQhMn
xWAD4o55nZNlYP22T9EV5iXTRNYU30SgIKK5VvlZy5neZGy07lntkiTBT7PtpX1MR7yb1Ls/EGbR
9wWjhmO2FtxsZd3IeT3/i5Z1nC+b3zKol6Y9ZJl2sMZkO3hCiTBeJubRxF3CljmNU+ID5hYnz/lG
XApJv3LfL7Q6vJ+gT+lALPnJ1mwyzu3Zsypd5mKX43sB7nANQ6vjRxqb7Mw61j9Lv3RBXDOG8RaC
dTvLgIMZWF7ILc5Hm+pnKb1R0DkYATSVX0vIRI+1X6aW4l7aYDeVGmbe5g7zhyZJy0vMucWhuMk6
fHLgrjZ1bKI8/aEhFomO0Km43WdMp/5suJZVmOLUdYFtFe+1EWxao6OqdtXTL/JhUxsjsKtHnmd6
+s5RP0csFPLQaZhNodtvcoqPgioGCurcKClH0kCK0PtNLONsgzaa0rfEwuPN5g47y1FROwzLFUYO
gf3/i+dmo00ibjTp3ciK6dBApAH0EVXnTF9GL08iUQNQyk8C5f568ntDW7Fr4peEf3pohqPxWGjl
1auKAoWfmQSlU/4Aiamtd8C4ggiYzAPY6Bp0YL9OhjIpUk84JpwtmTs86AKLD5/pT+pjURPBT5M5
ef9K7eCGyLgadc6O5sJwkPtWf85A8pLR9OmT6YBLMa5PPpsudLbO4imNgGfVdC0HzgHTXNdmBVh4
2df+l560mRcmHjjsQz3QoKHUrcYqHF+jbPdVL79hB3EpLp0ocOBxwrGPkfB1Y5Y7MSSIbn5YeDwn
JkCy1tojsaQGcpM7MoAxD3/HDJIP2X5VxlmYdcmaYGksIolDcnebrm00xijvCb9WQUC989gTW1HU
/k3+9v4X3FQay8NMFCMKI3yIdZGdTfDb40tJyMHj3Jkhj20M5a+FJFoGI8Hfga06lMuTfFhTSwAm
VZftRCbPWTi3HaNbE2WCxaU0QcjAKBTpLClWRkhm8d3as0MtCYNt/en7DgWFkUfjOhhijCrRahCn
6CZnW9C9id2Wk6Tc2TpjaFrjyXpQlUl2lVdAJguzxunuUpr8+YEA68l7wIJ+NbXpLhq5K633UfBe
nIpfeWhpfRXC4MOiyJZfIMaIj+VYzkwnWOA9DFupKhoLJFKbWE9EpRS5Bx6cqjqnusZkktqZYeRZ
FJWNK85hy6kjiqMT2EEcs0PNEoki/j2WwANaMM8DaqhorRBwr7IODqsL66G4bkRepabwLaVR2OlC
5K6pNjlIyyKwkvoWoJWrVcPRBJ9r+4HnaQPeHzU5WM53q7nkJlBEFYhBi+KNP1+8a8Iv6Ysb/kG+
6JMsVRKxox8QYrEmEJlTAjPKnUfI3wlMKPQTtRu0onYfxYf8y4/JnhrWjh9/YrRpuUrQIffN7QoW
yfg13frSdCS6B8/vbGAvFPJz248H7GuOuR0iG5QeahMbTdjuuC3IyWeTeb8SRlI7Vjwk/nRBGIG+
hdoSMlAY1ONQmVVXfDqubGisnBunu9fJNgB0CcGHY4zjxqOKsLCAj7X840MlDI/z5829r2dZYvRM
ogsBbYJDMGJqfVbzedA+H84v+s0aXsWt7TubeT0slsXko+ACouTpnTgkDQOsYecaD0etBRjciovk
VMVm5QZqxMQkfDtWbLRqP8ctveEtBSa37ntlsXMfFruU4MbWTVnZHuB+PVtsFGSbfpa5YPFkQCgj
CZPOkixL5Y5E6OaNO7+7CVeOid26uBDSkWIehaLKsI3LAia3T5ar5V4ybgrCUU1K0sVOluw7Cxcg
KUWiXqJgwSMOmcQ23IqNRzIzOMwjjmC8F9fre+LNXks+iNqf19T2Ovt/bzNGVRjSDKYcaDEBBRGQ
T0tIILrJXc30+3W6mOTgEdOowCVPE927nhGrmw29o5wdwLiMfrZhzJIV+g2evMx4NPjeKElthikC
9vJgc2JTnnZmze8Xh4yK/5Eq5XrLFgcrbGXFvFM1cuKmNr7em/dF5OTb3bS8Nm22i+INqgsfM4Mq
iM7NUz6PX/3V0iLl4ibKNR6h6125JjbaDzE8ci029Nqjcq6vxY1ZFG8PWRU6SfgkDHW7QWAkYJ+9
GWWredbVrzlcoz2ApJBYSpfQLBc2HvADWfUXl19fZPTkHHFh/kz4CDECeFbe0BWXus2qLFrT2FrB
3R/hHnWM2DjS7tkOepRyKL/wNcUNJCmBNB+Dzfb20QF02aMs3q6frwXOQyajpRHZ6+A+0Mb4952i
sZ1fivvKQzpaRStXZniCoTppa62nu5OrzmtxpOXlOYGNFfZZlsne7VWeMl7cgqcYVI6waigfyorr
i2IPikYQO+O7ooXZ0pNDX8ti5JPRv1TXCe8rNK0aMWRy1fRuA4NStuTXRuQQ23DkStzEq2epadsP
YzThB5m/xepHebqUDg8JiHaYnJ1XsOkg6x5dLuZA8WTmLI2e2OUXhcWNBdzasGSBmxbxtGWyi5C1
HDirMaty7fR71lg7ABGuV74bjNUF8cLtc/thZgTDJlWbkS/FZgBiD3PlTNuJKlOJOvQ2b5Kv+kRi
tZXdDcwa8n2o6brANvGAtfzYxDvTCRR9gi3UVaCh9Aia2koYzTtQQDLoWZLFY75smTApustV3pzj
2ZUNPf8DqCXgKknHDPcZ1erTtfMqU4Ntstg3aw0nntSqURetFCMUZNIA72HpetRKwlZ6vTSdCKb7
MqqcTEpY7lBCmZxJxnI8ueJihNWQGJVqU64c2knVFmDUKopBZaYmCRToNihQ3UUrUKzdeFiWMhwW
J6QKo6hrJC2khQpg8ETQuS8icofTiAeFllkjPinMRo8TB/o1CiRbbHXOlkGabI/zN7uj2KCWssB3
DulgjYyZ0hD4cabn+MaiKgNsDb/hYbKc4rNgV7wW+aFnGlykor/mLGH1pOVcHzNZzqil7oQTuola
7d+dPfQbr2M+FdHBlTQ4hkqUOduVCs0AuV0TEpBcvd/STbgVzaZxhZZh1+RNGKCdvowxD/uJa/3F
Q3HZFjZTau0I6iW/8WrG9u/mwxAvg2Stj+XXP7LEQffhJljMCySS2rzYJVKyUb36CMmCzt+E+MbX
ZGYsNKBVSi4bQDUfmtWoMZo4/9XH8a8C+lDZHVFlzhx13KQ5gcUtaPmLeRFB9WxWXGDJALOE/xxU
M6i0/qtKu5bW0MZbdr3UE2gAwkDZPjwDZQbbrCuiKkS8WWNmRnvmsA7yNbWDi+QBb7pdPZAmdmOc
c+r1kygPgJhOvnI3WQNVezSE/n3HosS1W0pZTiMjkt3KAOKlmGHZ9BSx3f4WIpPVB+u6jCLqldpk
5PFaWhpTvpeB/EStz1bG3Bhz/G3q6cdAwhb5GIc4IS7YmHXMDh9S9/JuNJInWxZW4t/9/K0imodG
G7RHK7nvGkH+BjNpsDSDDvHWkVIo7wXk3V72zKrsdY1/hIu40wrqAFTfwExJ9uCujjrUbFy3VA+t
GVwh7R0/tDcSWpvvYR/nsl4Ile30rGZdiFwoJKyctn3wJu7ml5zapVzVeT/IkLdDXjmHTFs8F1E5
Ta4gnO7VenG+B29Ie38O2iI4fKU9oh8cfUBWjv1GqyVC49L97QqeEeS8C0Y1eEREjbwMgNLqBP8y
bwWyoWMJaKHvAO0/2mAcquSR5MuuG/oJAPe0KDD1gS87Lo9MBBTCqeIXTFdThPJ1ywlpz/D+/cMM
qhlagkiGTcrmBtbZZkMmMDNlhitNWysMlyAl++RFGJtxcYMYdM7R/jEU03EUNf/9qQRvmxmHs+0S
aAB6JcMdvOWAnxQy3PTHNHvrOAdyf60HHAx4gdHodpQUvM26SSndVItEHcA7zLsSrajjoILe3FzS
5hmYnuqBS2GetcHmvsuYFuyZe0tSUeGeauJKyv2uAX02jRo2gGkAR7l58H5ifORZXW1IDN3UXwZk
7PgfEUscqJnN/kcNoTE9bhRroYKVe3uIQaF24YuiOuWnx8buBlZ683uWddVXoTc+T+pGKGdLRSlR
XERN8QR7Rr4lCS0D0uG1WRJI3n+95J5yiPsmdcMUVvL6N5E1vkGB6tk09k++A+YJeJw6f88MevoS
uf6ktFWcXdltzUtYIaL0hXBCVJ3e8r3tEKQi04Ue+3BtK83ML2GUEI0onOvuJjG4IxGEFS1msEpC
jGMXsDJzGgltM7M1jY0RGkz58w2OYHSMgngSqVbJYm5/bAkKyxliSRiYFPT1lM69G6rLcGlacqSU
Gzrony29+6/fd2WagWQE7odpK5/mRy+OgGhdXVPKuKH3WttdhgYsj2jS2MB0X61dGhknWSl7N2PF
9du6tojhW/bMsv3eubXblMBnVc4ezEWQGuStngvgFUme4gP7jri4elJngP5Qm1YMZczjzLPm12iE
fsnopYNJaK51n8v8COllwqggIKuEWkdFtRhz1gbW9z0C2+cx4si0CoaxcGLaKGlmuNMFMve7GMB/
gGJtT0TaEhUeOoHUhWvbCn/Z+HatxABk/LB51f37j78pSduXcs1G5/ACY6XQ2iIQqwtu/1bw6o+u
MYYi4XHthQXzVxNDB9FBhcGr8NhGMqjcMlw8mFSXIz0NRwPBUQBKMu4MH5WiQqOWzzTwJgJUXHmS
/gFbkkOqVkEvqDGDQhV+C0bxl/VGw6h8G2oayph4Ftms0NEe7lY2jWydafLnouu6iwSCgIRjJKWh
OuYgiP59fIGM22DeRueFmlPj4OLfCOHh0Cosdq4AB4W0kmQDqD0Zj9z+Wpcyz9Pb1pAnc6R+6hoS
/QP8hxDPJPe0S/JHLFfph3jGHFqWOY8wMIURjkKwzsNDTuf8HpW+D/EUzVfjByva3obrRcyF/duh
y8xQOioXlGJWQiJ4vec0KqSfRBXj9Uc3FlZ1JzM5FnrC/beaCnkttPgKX+IA86OvNVc8qOlw9iPV
p41TtmUI/rAB9YSLagV7Rpo0q+e5p2LjfkXGg/USXlMPVlDnX0ACJS/MbxFBS4ds9hsK4+WHZXD8
6IwiTADPgxm3cDUJR1CTGU5dLLxsOwiCNz/22+cJXa9tJm83W/P18kbQ0r17aezkr+vaptbYDI5R
lcli6e0SdQiCXkEDB7RHSbJtHfvbkZeQO5VYP8LR+misV2D8Mxsw0OLrCB+bKpuf6bFk2Z2lhyqF
7keVOivao+V0dSZzoaREtTBEtwRnsuGSQISUTc5B7dce5n55wDi9fhF2RCp/4zv7oWPq2JOZjW5F
B1q3qF2qenEEOnvVPLj8xFHbeZKlzhh6D3Hj5iVklFrF/si/IqC+YYfIBpPvWpoxB6B1CmxeCFkE
06rBSJgVVuWbGjxRzIgrX7pETZ/N3i294sukfqBO+VUPpQdrGBnhLDJoBXdZNSiCuZj95Ymensmp
dBkOKKhEJhQrN+/YZA0SzaCWkkdXLUDvn+Ir9yCwlqYcnnItJ1FjDz9E2Wp/lxq2wkSMD4IV78gv
jGWokMCtfMdsUepHV46/TR2jZWRjV5U2KCJZTdNPVSu0QG04NNLsG3YwoB3yQ+y89FtoNlK/XvMT
ZWFkY2gilnNTgMdt1dGMMThHYfhRot7MT4tM7RP0xKySg5fAt6f6HRJBcpboF+poBkYwcXAhdsgq
zWhFF3086eqWRJoSxt9VqPQrtIf1UuuLklMgwEMjsiePgoaqiw65DIyZJOsf1F52R5dKsEBM/FnC
+VnroFiRYd7ygF0jmzvZvn7QHbIe+WRFl0525gCDzz3oXNL1SnV6NcD5jIS31UkOBuD0inEqtwGn
oaHCS9OePKjP+CDeviq0Sz7mej6sV0BoQXHxhu0A1cK649a7E7Lr39anV0E05akKFybVSa1C6BJx
wVn83BufgY0muwZY8zdhIRMkREfADKWqVNfMf0/Td+WHR46FII15N4q/Ib/iG9N8uxa1BsJTqZ+O
RNcysg0c1+Y7GOGxtZL+VdzGvtTvFu7eTbDFUFiDtbn6SEQVULi6zSTXslNO7XZ4Rb/vRcOeT+cJ
0wzeDVVcmdcb0a4flTS6sPMYLKUiV/7LdD3pcnK3RGC0n2OCYfxytbHSKz0KjPBslQ5km1tPbstC
B2foRKlBKDX7jhHfc5ZrjBtZ6zbKHKEPvtDqyP7drejN7x/XyBMqvgdwBz/l47AF/iOeV3pZntqs
oddF4ioXKnGFHKB/VvISqjCiSWRKko4ljGHEe9wZxy8F7e18YpwrK+Gh8gWMjhSxr3LeBIDXdjQZ
2Tb+WtWKdnjIMaTV86mMAUXVZYhYduiLfi7I/QsGboTXgxI0RwGYzq8TqZbEhPF4Cw8UlhtSeBW1
OeI1OjEsGAc6NlQa/4m1ymqSZtd005eFxbrjMrtoq/1hdp/wabas1uf0XEcME72ekfj7jaxOKW7N
sw1dzdbXHfmi93lc/vjB55sIOnDOvVWUjd6FdFuUyeGDgjt/KQ1l57BskzW8Evrbpe/lYVOktLbD
0uA7HdA31DD3mXpScbhdN74XIQcgOU1eNR1VAfjfFoglBaPvVfDMyK7O7+OeHo6SB0eC0nEzJ2y3
IhZ6Pf6xm3CLNf+uXMJ9mQXeb1PbT2QIiZo1bD6WncCJmKiJSZM1pDF5/KG/2f/8nNfG7+21I0nx
6CVltAKZb4Dq2ldiGphYfRC4HT015dzAN61EQurq+y8JJc05bqsyypSxNQTjPOZ3kpHaNdqk86+k
PHdyCKf4HXMDBYQ0WgwOJlYKR6Eaal5UVeOgF8IPq6tuyA4Ue5d8nKB6lehgLw4UjAcV8bf+gylf
a8bJUbeS800MeonZ+ctsyk62zz8AMuUeCUgxfC8OrP5TBxRmflUuUukFGU9v6wzY5LUfXY44S8L+
OImYZu80OW9ptRkwrYSmUJBYEtomEIc7sBMipJXpKnPWYImnjceZ1j/dizpzUNpQHxQ4i8qYo38J
tFCd0TgZoA+B/g4KWePZeS50KuMKoqlCFpai04bjhFh6jJXviF++EThS0DWASwaZf9VolIneTB4v
YOlIHZeFLUshy5heLoZ8r9Mdelln/cMt734QHZkZATCkE6u8R3t9N56eRhooK4EmoW66Gq7/mIYh
oZ4bA5o3WmmjKNYZ9TqMY5E1fuZW4hC2hT/TGzXZBhLPQeCV8GlyKYp2EzWBCQ1e0JILyvyqSVyM
bgqgc0Rm3I7itXvRd2FyZ4MDnUwn2H1G44ssjCkV2Ig4yY/MT3aJSO0qwWNp0vSLedwLLCdvhZbs
5O59KzwoeUN2bDiIDO3mlXtOqQM+Xe1dZiyeqNbrPt32q28UVBpV5CHrmT0nWGAXLUMzuYe3Qo0h
jeVXFqvrssK1Gxm4QBv5u/3NCb2A+f8+6zROkY+N05lMnChoAnrnhWQ2YC9bDX/ZL3hcVFzJCwG6
eP9zlY/4hzK/rahWQASgGFrECUTqKEIQuW5g7cUeQatyL0ppdMihojcXUb4ypmdYBTDQMOwH8LKK
xnl9xR3MTohU7Y1DCR7b3y98lKjOO2rxZ0JgVTTN96yXxVw5sYBsXYhJV8AeqrULvkSkY/o5rd5A
Ws3iEGktwQ3PcePzdMW1qwM5uIPO4PyjwK7+I88Z7c0cKvlRM9VTGNV3i6uXKxVUdK6H8wAhTkD0
BIgXiMlYVjroEDnYKhlagIbR0P1x93TqGagW5++s7eQYCTpaFa9B9dwWo4ZxSxi2vZoZJsQs2MSZ
rGouL71yWc0eMPNM16pursrEMBcYEbb9Sh5StXzErFBSFqRJ9CQ2IW3Pd4+FD5uDP2Zi9pBb0FQ0
nef+wqaVS3hYArgUGTfXwQLNWOefLL5qu0p+FldsQ7CCVno2rABkXt72NtZooOrVtCdocQlPK9h4
ijjMUYc0AUltJzFDYEOjZMs9l0HYp5BVaX+SiZ8u+bitp93uW71NkLNmB9vjd/rbSZTtFDp5cgyl
GtuPeeRRelFzO3hdVwPNdd+CGoMNVpUTYDCh5sr/y69aMBw24beQRgltwV96m4Y5o9coDHLs+zGj
tcL6zkDiYC+b/ONfstaMvhAKfJKSV7fMKDVLRn8zCtfA28yZr7IQLzSLj3Y62J53n11RcYBdEs6f
/rMoPSldjSPsyRDRMFaqlD8Z9wHxogIDLrLqNkD6V7sMxjR9hwxLW6Xn7NVhb/+E/IiA8S3jnl1G
tAmh8j+1GqUmoeb8q3vBXGU4g2KIfbbnfDFQ4LorsCYMKMP4WzpbxxQOpokeUhz9yfCzsee7r+tZ
Zrjhm25ettkKj4mLkqEcuJdSdBloUHeMvBtqKRku2gVQ1KQQFH+qUcPoQaIg8APbKOWVJI8FGJ1Y
08pXsyw6X/KSTVr8NorFAk9gfyPgklB+TCbWQ2ZI8vL2lU+4MzAUEwHWtZokFHyLPf6UcadwuGgV
AlSAg2iWcacxT+9GhmRZUfudFhfmKXgHUI5kVDH7veL12F7sB2SovJsld54SyAXauPQoK6unTH48
kYKeSz8URaO08iMWPz6AZQr/jRLgdByZBr1QEuOKDq4TbbYelyKY+c5QHXrwxk2pheNY8fb89pNq
c8+CYmIaYRrGAxA+zcm9uRNnkMC2IvG17nwRsmUJtvfvg+/v0vwDgVAnTU2BFP03twlfoQXLt2Jc
Y3IsFRiUBHX5Xxq1DjWYefywPZty+wjigr6DiqbzodEqTFYqFo2DkgyC3rrBCYCWAQJWQhvjUs0m
exsggzIfbctynNUMZjv/Eoy35eSCbrZ4hEW6gsJH2wQsZ3NXni0JCx6z26WNTwr4daU6cqb4118h
+kL9cTSUln94VjcYRy7OpUin+6bnQ5xPlETSEbUimykq3+5QTsPKAHS1DYwKQ0CMv+Ldjgaib9d9
v4d3J+SGS30oEAPg7C6C9KqlV0q+QmgySsDdBD9AF6EYLCkFRYZx6lSk0/eLK8PNRklI87dGvOwI
bWW8V2ukv4OTm50I1XUsHY3e8OS/EEDJE9si9qnTY9aIrG3zVFYnZyN1ocyQF3Y9Erfk7n8u2lT1
X6AAXRjyS697lzN/s3wQ1OZXvl2dJqizWdeK8noFva2YDz/6HC2GH0sqpBAyhgsPCmj2pcTBPn4d
nQfXKcUpi4/afioGXgqeMaoSIOQx+HmjU45dFdqJ/fhyopCpg4tpafaUJ1p+myfvz3auUGe372o7
irT4sJ7layqtndXl6qU6NqNOn0VTNNA6ZLS8v5pHt2CJeqkWb/XyleWTjfuHfbYV8M5b/lohXf0X
iXFLm0nJD7euMW30q0cphznnDWGxtR+czp1DBbsuGRjDTqm9OI5G9IOUFuDrQ1wVc6LZtJVJk3oA
/VRuq49f8/xtJNc9MafHY/s+m1JTfSKmqF5TMzFab/4IWwlIlMKwK58uTCAyNY+pybAtLmk6YcEq
i7GBHQ2Q8WsCNQS6RDWmlNoyboEdum9tQTJtIMeWKgrtFltQ76vNS6uQrjfwAesGkCgyCOzcoCF5
50UVvu6/JD6XlSEqV1A2haJx7Z7Z3kghv/oOptAv2tYEVQ2fcrNK1c5CQPDmxVSEOEOSA/74G/RZ
XLfQEB0lI9oJag1OZuQI2tqvifnQ8ylR+6tECEanRjapZJPbV6JfzEC3R+KMFOZgXB8b/FSVYcFI
UpmwLEAPm1bsG+dhrFoAUtgmeIKSQRileelHzEJhEBu9+x7nLwOUCGRqiv1AjaazO3etjAtdrm6c
j/1vigUcf2fCLXBgRsbArRDTZeT4LLJ8a041QUYDNkU6g825cLtuS/hknh1eESpcDqUAeDEbgI3i
b1EFuw0MVm6PQHu6nSUBad1O1/3VAMlTb+OLEZIHmOCks09P3MXO9VZ2h7I3QPWl5unjRJY7xa3o
+8toiyFj0ddFZ52IlyRCTM7m6r9q5Sa+K5qq8EsEF17EoKI6e5EY9YfwSnAdyClfO82IYjDEwR1b
DPecnHo2ReToMHs4+/j8FefVydKtGRSq9vLdDXpyDA8KudTjgWltuqgs8c5Jon52d2jVTt+MJ5Dj
S8CSlH3enn3vTx1Lu/HCbiXUgdZGFZl3BuktIYOQv5kEb5iZHn6N9p3/2HzLrXa3+qNLp6I7aw+J
FxXeQ8wSyprHvZWMS8zbep21Nh3sJqSyzZ9JUhKrE0LrXaVwKbSR2LNENmK57FAX2KRp5eyRjB6J
KTHddjM5k6mzuhgx4ch73unsCkqjJBEsBJk/ow0XdFhO3WC3+ySsiR8W0yhSNHEt2Q/6nwKuaHU6
yZqAk0VvQYiz2hLI8RqXCNTVHuRjNEVRJm8z07YngAm5mZZHy0s2hy3KepFn1ag1JNjNonwHpX9I
VI6bBLi2Cv2ZrpR0zLi/CbIOp/5cAwDXhc5alzVJBAD4j/LBw1XCB3Qd4qlgi+qufYs2UTM8Ln3c
qB5DAvzxKGmIrfJN8Qf440k93TYFo+MO8ftLZp3tIFmRhi9u7eLigxIYTIFsQCWK9W1V24pk4Nbu
9jY1ZRsnKKg6LIneba9gX7n7qMwUa3sTJAKl9DWVLENdjFFxqU+knua3FSHrMk2t/i0R6u6LD8P4
hfut554bQN5X5bUr/xgKM3u9OQOhOG2z7MIo3R/V/kgTa4o+2mV3xcuFv9h3G/nd6mQ36xasyvpP
nRGMAnXrk/pGuZMZMTNwupOnvom1ETr2yHsoTileD668WaufACjQwINuNwfSbLSjYxFvcxnGeQEU
GDoT9q37HDduZl/ziFRBKCe4x/m6Kvyq1sxoNwGhVMfmnd02h88IKBGOiDuSXf/eEst9Vws5Xw0C
gTSoWYK6meBw0Yh904Yln62KQXha7Y33ttqExKNJEe2or7shP3m2uuEOK+q/rffMk8CiYj+gKzQT
e7PsTvgRuAfSfnYwG2YRC2Gj55DMenur7nk9qS+oUj3YR1zv9ZgbVZxrjO5NpaJQB8Ix9e7MFHO1
4YueQ/kcd+iX/ywZJNeWREg/TbA+CMev/CmoIf21hys5BB+qVRTvLmfTcadwTeem2wXwtkG935vV
M29D1wPiBvl+i+OtKmIiXNl2tZ7i4qHa1d/xnMR2uQL/+law+Bto4vSNG5IN2RZoEtrG0PJBASQ5
lzXKwVhd3+KsgHaE86Ccgl3wQy02Teqb6HgIOKyS9h4AgvfGwhFmppB69uZeN2fdgmro/iJIyHya
JvIgQuXzD7UZ+bJZO8FlDZp1pn5cHAmwAVFA/eK9IZ91gU5NwO3VYurJSg4i5UqtnuaqKKfc+iUn
OVMxVg8IJAlC7q9gHxgs9hH1pSZqV3fz/jnjZCJ0WfBxU+emn+v9yu/aUjoVCUEQyVj2Ek5vmYcR
664aDg2HneC9/fpZp0oCq0YkbUWvg3TmIWWCoklfOyTvT3jw1rQXEqKWuw4C00SzgeeLBA1Z0xFx
GvhwnVLwrGtAPhRN2ZyyWe6PLvENGsms3r2gXbF4dSyLWlO3ORBemBc5kshjBG7JeBkZpZoZr+8G
DUo8ExMrSReFFBJSnVILpj8582AW15D74TMONQ6RH6zTbiv4fXqE/2S3sSd8qsOQzq5xZYB0QTRE
l+SqAnYKy6ClV9Xo6YQuszQNxU54OZc2pIEHSRa8tf9717cimiy5H7BLEamf97eSDDxVaOliQckv
24TXJn4ilud8DsaNn4Nxrk6FrumvOmqNnG2fUtyfBhPWuckCbJ/Uy4TDMOpPypsVqAHUd4t0pyke
Y9oQ+CFGsfxq6UqKB6e/jcGmBPfOdMrGTQiTTUaGKAjq2v+w1cctczhcx27q13F9h434M7wR0gwj
rk7BwY1+wc6cu5y1247lv0e2YjrKGKfqpRSg7bzjSy+gWGRvB8Mo5EffyStKY17EmBVOQvX+dayw
KAnpF555thCUXy0yzhM8mWDPHLzibdUgu+uWMwyuk4X6rge+eEvBPypJ2FQ+ETwLOkHYURhmVByN
nARBhgM9B7SsLGdUnXtyNd7PMN3qr9+FFjy8GPQB7QjgzR2s7Dmeb+34JuZlceDItwFCk907g9Ta
2lNOFoLmofCMLZrTGwBrB8tWney68LS6UR+P7KtlWPwGZBRouiR14CdC/1iuFg3wy1dQ868TYVnq
ufhQXR07wgDXmOCoBmh4Q8GzZQFZearKBHQs561JDUo6lifkYA2MH1VDJjqPF6wppTnDXEWbSUje
9X+aNjlAHIoQjVaqMyadFcEiwsu4x5gWp/jdd/D/NxMXVvL2lSs46Q7Oxs1zDlWDkpBgamWmcDLE
2FCYvmA/VYg2FsCJhbE48yHrm5Q8uPUlC1vh/g9aKXgB+wrBBDIPKf1Krl3ZPffZ4hUNlTkeedy+
CBC/PfnGNd+0lBAbtdcnLfkwLYBvcpC9GSCgbuGw6Uu9XoMpQRhMiIFXxN0+hXrtoLSGGk1P84BJ
O2vdwBzCnlNb5mK57/V5V9uQOh9XOEHMQsicVSHD/1wtECExZzLgxDNJPEPj38MLZZcBjx9RwFQl
DuWvveXyecfHiHm5EJYcOOxoQ7eiUdf+Pv1MTPxCVnloWzmV9lmDv35xGpT2ZqJQfhNrplfDNsaE
tYD2iCMfIHs2u3Kh2NtRZbgnNVken+/8ghxqxLoRQeUNBGSBHTYZ2O30kO1r1zMcMW5yy9hL6Ayc
ta3XVdkFX64c1ZqVP1aBn3A2ESe/k9UtSB53OYgVqiOXOrLkT67rpgfi+OnLsAjzdBm93BiyYdzO
uS2bPG7zyfeyXtI90DXskIi7G7yhirVp5dIXjpRvq5qRSAviuOTekFHYFhF/ZHdDcS/2Id8KPy7B
umkpHIF6KlzmLgo315s0w5cq8qNdapILMd1wDfwoC8fu76yjtYQXg+nPyBdA0jbxZaOiMLgjb3sq
nKDNsdseNCVg6kFX1IP9EaqPysFb1WrHSENHfF/Y3MkrvSkWAIexR79+H0EFtheAdOK5xE51y37z
1b/Q88kE9nl2mvoFe4u+7+kxUlWpODwrjPDwe8U7/xK1uJnCmNaAaqGW1+eBjaVUaE3mxuQA45yS
Iyd0CTgiRfg4x/3TmNRpV49uoNt+D480FCkFcjCNPjhoUBQV/GprU1FDPYGSAj9yzDGlAkk3LkiR
K9xnhqBU+8PqGZxQmF9iDnY6/FfZwEONn3+TT6vpi0K/ixGgT/ey1yCWhdnlJDXzJ2/VSrv9P7vz
cY5T+WXW1xfpZXgU08NgZawtVeC19ALswKC6bvAPtta81DG1WjLTC6PfIGLewmsIF00F7KSlHvMq
3KROLjs3thtP2vxXdi+IG15jZDGqGvoHufkwjl8o1E8oC4yHyrka/Jz1DEKKw0XBJMTkBmFlUG88
Px73wZRNyetRE5/1DQIh82Vd50QeNQYIsOFNJSxgQjIsoh+ujE4erhwvDN8RSJSk8022ongZUEEn
1XlsbuZrhNZql55PYEdo4ZPbxMuTzzrro4XjqJXUkAilYl0aa1kIeZDARiaRwuPIuqT4uoaWAKc0
5dGBZB7mfhf6xpShpBmiobr+44FOGIlsPSaX2o3gJPQxqlRHww+DSP5TdwiRhvgYPuSDsPlNd2dT
X7CQ8jRMzDsAloeSIPHietks+T+rrkZDt957BrJ8Rlf7CIarf2NFB/b6Qgf8peT65XFoOIbExiD5
EF8BB3NnfVm74TczCTMvwFhLp8yxOe9CrS9MX/0dnHIJBjTMJWwZbT1iYjI+mehW+g2rTOmdyqUu
u9tnqXgdTL1r4lJ4OZogMrpP3N8CCE9gYk81v67FSKcTRvrI18tVhKpJIMeUjKu1BQ/jDr/a5/tJ
vuNSAZD0Wr8tGmZCS4/I/0ZBN3CiQG0cGthSXgNVDt7JsEBa4j3JiXg+Eot61cAoYNNMToTz/Thr
aeOcCLLhMYv2+mDMl7PQ2FbWUpfWkXzmo4BWzLQgTpnLihPCcYbjdBQJQvZmSoI7jbno3MNg4Eol
aBk8xfn5XSe1L3UHQaOLJC8DJeBNN3q0aEOuI5RWTtBbvwEjhT8ElPCPRYij5YxOqxDetA6BQ8Wc
bZs4OOgb6PBKoYBEmtLx+W1g+KYdLiUNuzs1V+fcl+/RMAoiSX2CXejb8hZrUTQXDjmNMJczuq/M
r3ge3fWZV5J8dVwEwGm1goPX6uN9rZRiBB1mVHd3Q20GEmIMDw/m9LxEIQnLQIibmwz9i9jpvC0b
NvG0VLTcad/286tvpnVpUNGJGY/qQNwGU4PVW/ofxUnPSjnYsdC1W753zGfAxUnp7NwQFmeI6rtY
gb5pix/NqwHEOPHrJdJcul6hLq1ixtRd4jQG6qkpUucDdV9p0pkkJNtdzP9rJyYcI1foW4nHHPqf
QN+tfX2t7dlQdJQoFtKUWDrxXE+nWP6cdG6L25z9+N9CDpvC9A6uRAb+OockOZCE4eA/AbQn9meF
GNe81uBKga94UOwglS3AyCkt5TU5f+WfsljNEMG0Su7grsdjfQ4qP3KScpsOzPzCHzMY2Tpgqmya
wjflLTSS73sz4EE+Z6dKu980Jm2ldX2LjoGrW11uOLgRqROdDFgY2S3HOhzZADX+U9BTPVMe1J3P
RjOlzbDGyM0osbl+c766nv9vFlYM45gWcPG5IhNpYL/x4fofujoSlajQDLYUKfGaD1mfA4OJDjE9
qVDH6ae+MWz/CwyqKERcYLVA/dIyY+Fj+3WgEJM6foc6wzBsZvvnm3TO4OIpHHERmD9R0qgTPzs7
XRsS58Uh7nn9p5qVmqtSDU9XC0PsiwcoFMw57hPFRXo5+k04XS5L15CASsC/r9HDkTfXczpMGOYw
LC9fPtX77kPd9FwM/FmACHDso5ZWIXxt4sqe32YB0IkwOVZEh108D0/DY/zQkXxHyRghXNPoHgK2
UGgfe3Yqq9qsxnjdyT3v5dhkPf0aI7Sos8BUOZtNx/gm8HFlAOXr+PWj3cuJqTlY3ay1YfChlqmP
IcsS939YlPE6+HcnnvkKCKPoSngqIWBCApS12y8MytV3p0O27LL/4vsjtF2xaoQEehiEd7Vke4si
RtIfyLvQrFx6TmzzvQKbHwgMOPmFlZV8geE6X43Nz0F3whT3wHj/QbTGO8K7mt8eOk23B5bqzMGW
iX27Jlh3ICbEoeBQ0gyF6dPw1g3TXk6yXCUCQg4EvyG3eT7JLf0gNX3102K2A7JOcoxBHM5i+xVC
ifioCJiAK4dKDmk2HMb//B2wnD3j3yItLFfcLK4WESmYM+sFG/rdzW9l7jo38eEfksZQhxANZQOS
Xz2z7mI9yKYrXCgBy4a0naeZnPtOdbosCu2SgB1W+ejXgYhWmMJ77qip3+5skUgpm1IRb/4ITdSf
ZDr5PLqfXdtmz+00NPYakjLxuma5bslqZeWl7/nI5GT9TeDtopOJl+qaCXdUpvghFz4maVWFXHrU
smxnK7zqJL5YBaLELtxfd8RxVJvuq+mJWrvefc4Pt+K8U9UdDyzfrIggFxE0Xf+m/69w0cZ1uwzF
DUeTV4UcoP7LPCUMlAi/M13S2SiY8cBUU31jAFGps7g4RjykfUMkndS1cUAkX8MzlHyGgr3XpfSB
E8BW4Ntr+FCimwFxAsCqNv9mm9LBWGxfEyDeUIjp4s8HzzHQT1BR07rr+EL9HumcFh/2l9HVgcB/
UIaFOYBLB7hawT4ziHTLvwV/LLwU1ICN1busrCgfS4NuYj5O3a7J4jD09lFoYAI6rq5X3Ri4cOnE
4j8FFSgca1riCkTTEfU842U7J9tDNN9ncV5Otm7PpESRUjpxkXQiGTlWvYRNJpjv1OICd8O5yEpX
4aI8gYo2DHQdOtH5lklJwCdYppPT+5crcf1UBwZqw1J1YmrOrN4uguuOVqWb987MK2tKam0eUpp8
L6YZ3V6k9aTh/pQO8+i6g8DfQ2pDEGV5eUAw7FOyp77TAcHTVdEiW2ML2pB/x2GuZJXmDTDjFgSn
WTu67gP/Plb/rgXkxCA+0bbUF0GO1fJcPpAK6FY4KrYOkgy9Vrn6OP8WawLIj8r+3uvxdFbWyCPn
W87L3PkB3AK+32jPsWh1ZR6W+YES6kPN3SRhQz4wsnLZJE2q0I04r/MYzCj2S1Hoi/EGOyBnM4Ok
JTTbMw4yzQTVeySjRpEmS0GMyYf9PTgVGLvimddRptImTnueSuR/1Yzp3m/E88b9E64Ce2u8y+EY
sDDZvHxZ/VU76Dy03QQvLoUYCaOFb/26SBIOG5CP0ipoiVKfSeZON4KeUOnv+ZwwsL/Ta8ui5nqx
PLxrK798VzgVm4QR9F+VUQbBdaqrOmWD/cWcbymD1VqIT5eyPDIsYwDbLKv1DgegmNzJnxyWiRUm
+0PhUQ0caSr2n/MOkmipFp+iUvrQUPU5kiEhUKGmtaqKjj2iyz9UQz8/m0M06NNHQU+OYSLCQjkM
AUfxTHqn8vtB9M/FTqB9s92qaF0m2+uFV3FUSIeurXv+AEz6b03W9U9ktlGkhgOCF13nWHDDXkwJ
M57zS6jwxhP35ad3xu9uE1WEul9417W3fco+P9agHd5mAr4n7HNg+LK8oX1HnqhxJbbINvS/Ccis
T5ZB9k/srNoD/By83P1OOC6SdctUI6pF1THKDUz+OSNJFRpAMb7/OuFIYLVRgs2jwHi8YvcApl3J
+rzSyxTiyPTzfV+L+Gsj1ticewlKsg1sZRlswrhbSEl+xjvGu1PEFdh1xdKplVpk/mv7Qv+etWRE
bYnree8j9aS+3hGt0DjV4DTpKmzuPVXe8OSGIYXKiqsfiHc0uJ2hDZzaEBpXZCNORk2jq5jonPMd
EzblM8Hd9tY8NFB3tHieKSOZ8ZpqYt7wyz4fSl1HAXLRVLFaARZYAFNlcat1yrqwDeLAKaaDD7n5
HU50Tyz29wrEqqwXbBe250CJo/wsw+u1v4FRT+FT2gY1snNXFRYqyUTl63KFLffV9CnmfwaaKUZh
PLmZ9k8DrWrelggPdYHLa+CHv05p9prfL5ev4HUil8YNagyL+T2PsNOnZuIdqCK0/ceYzNyHyVQT
BbAUZv5N5nxpiqXBVByEQ7XQvVA0mwyeBJnfWFRlSAUll175WozpYXNftTukvaXG2gGD8qqn1LvS
SePyLq6lK+aY5u1WDuEhRGiuZ2vrwUrWrQAVMKYSY/ohdrOCtcHN5pGNdaAUxSmW+Ou6GIyRi4NE
uXsreS6FdQQvmjpJgaQNrN2KC78Rm/JOIOVDZG6TeEqRovmKgduqMu5qx8LFRsyhjt+yIeu6EyAl
203MNlcVbYltfZZuUKbSSbNauYU7Emyp0kanQ5ApTiR3RLdY+sHkUHsXtFaCqKUGMNaAZpcxBUij
bgECX8TpToO0A8UPt9oGqy35Fyul9zZ7a+v4/8pSyhnuC2kHdli4dC7zrV1NLsFJ6k0Jk+krUqCa
ThQQdGlSJoeBXCvL863vGkpVPn0lIVrCX7NqEoLKLdAUTFpF83ekeHBGLC3XMM1Yq1jNGKxe2320
2Yq3r0BcRTRMKtoP5WtlU6UPbWfFh0BDhSsqdWCL620ZvrfbbkzQ8ptCdY9xe6kpZJrcG4pUX08s
y0G9p4ur3X/2vi4QmobhBnjG9xIAxpe2CPWm66N21dU8XVgoXhjHrjgtTdtkszA/2qa/1gAn3XwI
Y3jdurE13JvAKknGID70Y50S2yz2TEnaX7RkKpwvltRO+4gaoe74TviTl111Ay9pLZJ1A35RLed8
5aeLOEwZYlJJd/SvwuF9EYPlCtLrf9m9JCvOXFrKtQAbwHCY+V+Jvo/Wo7zDQ2iEzeCBCGkWpCkD
UxZQ+vgrLO+ZMUZn+llVdD2zoKg1k1j+OqciaeHvacAByFWRMKOoUvc6jTYl25/hlr96iH6vklao
Kc5j7rgqfKWhKBAchEU/eXi/vy0zmS/KJrwWh33HmHy4U0ObUueWtE4qHGKKdfMMBqdbgjR0Rl4Z
A/RzB6zGtaF8dd6TOqQEfd2GKytCNs+NAxcJra0kTYkrRXmt+1+6clZhoHBQEX7Mmss5qmbq1qSW
UoYEj86/YxrigevIo11tDXIyAONKJj64HPLuKBkuylehmDGcnXi5jxXATxFBVuQS5bTZEdkCfmTF
i87XVUNT6qarG7z3u8ZP5xP6MA6RcdhGbeALq8Uye8L9FRkljPDOUGftPxWQAZVWCrlBAQkoT/pa
02BhrWoJxqreHrEYPPKd2ManHfdWuBzsoKF/wMDdfjqPoDENKi6lAUbOmtk018IMJZqALcet8NuA
7ld6oj6eIzCVej5llqGGXmKLRo6mIZQIjm0usKidqn9MlcwvQoBZLuICn20YXNPerNxVpfc+NXup
+Shec1C6wSUe1ugGn7nBWNF/4PNBgKKXswr9gjt9cP/gxr91fSXaMmRdZaiao1CjnpPjVu8fyzK5
LMfRL2rxXOitUpe0LuU4NQBCcoaL0YVsaU8Yyt/mThzrgziClYLzogNpHQ3+5gTGkB+9oEvn1YT+
kq2w9m1iEp/KyIRkx8VLTaYs62L6epjp3sW1QdlGtI8c6S6T6xYmtXE4zC1pj+LKxueCDntvixFt
nsT6rO7EnrsO9flTbj/ErPVxCMwmNYqIZsl1xnPj0MuIRTISs3BhQwI6mq7QH5GvlCpoiwj7ORG2
hUKKIlzmBN7/p1Q1I1ZGrSuPZ0HrYyDWs2fxO58kJ1FKt8cQpa2fgBMzVfEOkirmEgySrEstItZu
vIkCMsuiWHfvn/30u3nAEgFbod71sdshyxstoKeT0RpZCReAbeEPNQOWE7C8fTlm7HuPuLJY0GO9
NwDV4ppHvl6hLm1NBlS6GX2W3wJvJP7bAXRqzPszKx0uLMaIntK/Ab8ZeymQNZUuk5cIvvPcHqWN
lIGMWAGARW8tGCbrM4+Y/Q4eXuDHgFFAAYJgmV+DRMuLWO5EQwf2cD/VOOlF9oLiZW9+PheGkGZV
t47rd3B2bAAhHUDR5Cx10BUcN1if98d4YICBCgQbutWsPi6ETlN/srBY4lbDnKWmAwFCS+SpmnY0
lDJ9YvFnTdM+w3x5KERFVk1LEDaUEu5b62Zf5CPcCoGZcmTPbDUWt0nzxKaEQztBsgoEp0A/qQrB
rqEcR7T8xkqP6aZZnpxAiRqG4qNQP4JOes/zAAU9Xz2qGbXy6+OY0ngHK5btHA9UMGyNHoFX1pAw
vMjFS1uWFi01WDC7Sshp6DKYyO3gEo+guqW5PiPhAWsOgDcGe4L+OQEhZx6wqtxWDYfOCnF5l6yJ
64WfIztCIuA+RT7vJPdWoUQylUONcO+b0zkEGqtc/YTSPRu+KoCXuG9ZFhMMIS0mmjvYvcdhX+A3
ImQoG0yynM6QoAyNelfyjBm/YdEWNe7z8WUraSKH94IEEEQ8UFWV9eeqWF85XKkP8Um2KQjyy7wu
ov2zPz4z+B/hU9b7UW0Tmsfskbbr5OkpjTfarGnt7xRts5f7PGRXHoIgvdIirkbJ7qz6Lk8nlZFm
YCvlBk/nE2UJOc9qp4cnJaIPuypUctylvqdcT8/JmFWIWN6ARPhoZ2jyncBDcfsTh4sId5KRYs1q
5J13ZWjy1ydG4zabbsFIDLIV+8q0yhARSeJ18bMby+pLo3QZ6EYrEEy31sdKFIka1YVU3bSzfb/U
Q/QF1RcTT4TF6EEY0G9EfRKGLVOzQZp0xly4tKeHeWfk0o+kB+WaAJOCFvB+yx9hhgM2eP2gXr2M
RxInnY/8JHWBSCfXrx+MDiMF3MasBDHvHerq/Xj6AWIqMwFKLZOuiH3udOAVq2Iuk3PedYoQOf84
rP7nLWnIxscKmWa1BV5gzSNdvUi2ZFJIk3PKGjtaNz1sOtAE9q6irQdxh/Pc4U9debd2gDFsSuUk
4u+upRfE+AqDbw3YPMY+8ksRowerQXE0sgCsUv5lJDzC900FlqmOi9kayx4MIDAMxZ8a+v+O9Vkm
TJOBZbzL1eFJsBaGViLC3zeZTOfG2h0L3KYdHtpjZYpsX1ThIarqP2WRqxjo6P03FD2VJagU2qEV
ThhWnySnb3T2JPaO55aXSShQi1g4bwtqLMVhcQVHTfmnEm5htpgbgYxL1F5H7g93WB8VZ76LvFOn
saQTR7wOOniUlpayILe4nI/jJ/vqaTK3UZZOQJ7GNAZif7WW8FfHKJFdEtVGcnwxOGjwfg/yn+gA
m1fgSSyegsUOh4ycsSWHhx0neLSP2EISMLPMQdXTGj2bu4aqT8vQs58zPc69mo6x6KieprCtOfSR
neGGSux851QONdYu+o7Epg7kloNqRYolULiwGbnLB4g7CegUBcaPRRoJDmGlvyHc/5L2CxFhWI++
C8ycZRoSjW5TSgNUCfmGYM2mhkEaBwapQXYeju6xZkA34yJg6uxcwpbf5ghchwsruoDRNjJHV6Fq
lp3waM3ea7oilq1b5QdQKyP+dvlX3ixwYH2yKk33qlYZHxFDTkEFtXjV8QL3woic2ZB4B2fbRoIk
bXbsP8O9C0B6Qwv+OS/dJFGqBx1vD0uHLdEYlEP3yjtpSUg5C8kpK70JQy5+0sZkvuPnttHo+k/5
p1qmZ2vKVOPodWpKpCk+Z3AG2ObMPdU9VYxfl2SbmprZFj7VlBd53Q0b4mSY0K+1qDcI5Rm+9Lov
b9lG9anYiITwLITd6FagtcI25iLHR6AhIPxCl7TJvNu7meUkFsZRWSw09adFJbqkzKwYqWI08iQI
qYh2yuVfIgUrUVEsJj444HZ5VHq9f/eQkQu3OC7p0YChkJhSG0nszc96axfmw126pV7xevyMMDAR
jk/2sQMjk2HQVmNpgPcKvUMmS6cpFR9j/9aYj9RKeD3TbJcE7iXL2L5YvGWhZgBZ1TWNwyInpOcm
Yr2jH0Yb0V7cIb86ZQhnUy8WVOeU+BxK76QzgN/TjkxfHh8DC+qxfK7DBeNN6GEQ/bMsj3VBcCQ6
ACq3VPMKBDjC8LqMnr5ksVRtN4dfGZs73nI/ZierxXAHltTCtQRZ6A9RHfnpHY2+rMEkodwsgc0Q
d7J3sZ0b2S4O9CdWwz1z3fpVpzVMMLP7CAo84P4OERMuot19pj8+sF1z1fl8V2OvTq767b39As6V
TxLTPr4pr+x76iuuVztnsINpc+U/hXcBIaLGtMKgD2wJ3MTDkFMBkh3mK1A7sfwyD5d+TKFPoq6P
8GpOKD6uj9ziXJXtmGyFv6XZPaAvMyk1eSTemJyAoIjLPoVPbIkBcjo9x+3eBInJmXG0ZpFFIaN+
nAkfr88/IsHW3GfSM35N2B5fCoEWHJBYm/AL2NBxh7cMtOOkI9oHqPSfkEDZYc0xrtKXoNrOcPvX
CPlI/pMExNR+gYxkLXcuS+m4yKEiNgyoDr7wAL8nEiMFdVw5rzeN1iw50LzGwZrEr6JK9/gD04y7
xmeVn63kEfsE80cxr/V8VDuH/anmwd4/7HAO3rKw/ADwD391NP/cKZMxw70JUcZ1+2zxCsx79ra1
6tSTYIHts15A/qTDYeFUavFjHxI/kl3Ilwm8ft10zhmyT0RurN82+ymOcbDmRANNhb2l879QW1Ed
x459tdcwjUhHsRI9vBueCV9VhOMXxwWo+U6wHxWfXrvdTwdAIqJCGglScnDikcCyca5G5cwBj7VY
rD6b3NNkgDCVee6qRT9xanH+4tjTmuyNr1NOMkPapYOCSv1o2LUVq2HWzafEaOeE9EQfF+3wV7C8
2ccGtXwvsqCQoSFWOaEblFBxoj5Q0aqR9S9t714wyRvtwJ0zuavSzV6Qpx5mniF3K5Cnu4JB6DS8
EC0feGy0MTXzOE9TN9m4NEv4SGQQYfKDGyCWueJyIPaCKzTiqU/d76aEBkBZRMKTVsrpRKnEk1m7
qxu6M5/oUu/PBtPs9rDBYVz8DOk1nGQKffWdGARRicq03Ku0xR2DkvNdDuM+64YBu3tgRD92fDWJ
+3Vw4xkBBIR94F+5jD0RvaXSwu7ZM5Mg263GNbqggZnN9WJwQ7eqQ0PyDmMIcz/W0g2UrT03Mvau
XSeHZTTrfXWS4Ph3aghx1YFRXCcMAexiXEYwV+iLIvlxY5wPXx4Qbam03BRsykfVgT8UaaAhoNR7
0n0U7NL3nwDiY15+GFXYvjCqz/G/knAXztPNLIEwnAYW1WndaN5R+lwH8OkrjUB56QKuT4bJZ4WE
QrZUOmN6mbayE2+/Iyxmr6V95MUojilLUDH4e3kMeHFziYSxYRrYZZym8KG0OJDlv+52S94ZrBhy
G39+SVRgGp7LjyteQcb8YTaSUTJQsa848YZy+Fd8NwkCFdzA3oGibXHhi9buwFeiyzvxGfB88U6w
xZLUaOLIantBHKwpRn9Vfpq1Y7SUwtYJFm5t68OvTD14f7k9uzu64tX34Y+6wkNMSRgutJLtyl/N
TFGYf8TCTC0w53wvMFjntAyHeUun4d2QkfW2oCd2hGwN3NxfItLizUwjIZMV2Aq74g+DeJYVbp3l
IBnLPQxyHMPLCMYW8++pyaFY3RK4nJFo/ECdVUD3Huw6pEEG7BfIGkFP7V9mnTq7Qttt6QCKCmy7
10HdWixQcxmxw2DdfcTodLBuwp/UoWIeucckre5G4FMrJugst9Eh0YnEhFVC41i+hsnW6PAkGfQu
AvtTah1wjQoKrlQAA2z0YkUBegC/iaAawJODSytDbkE56f608o9tHFS731Toneg9gC4UBI4iJ6Zy
cj6tlpbhusb/8PRvspy8Hk0ia1nSceDcCdSfP8FXKw+pxZqGtq+W6+AvvrjnMTWNdDNS3pMGh0B2
FvKIiJZ8sz/kIUlmtG6W37/ipegoI3ZaW5l12A8h7sLd0CdxNrDHTD72HB6Ufwh6e2DJS3P2m4Id
NF+keasqmF2YGFt8knPGfOr3BeZWwvwB0XavEdpy5J0hsJhqgHo6gVfNbXNSDEWVk/ox1K3JJVRS
MRNdRH4gD67ttbYj9ZLnt12HOKwGOJ8ngzned1YyxyZtFwwoam0qVCJ73G7GbYKDQlTn5cDczTe2
ko4Pmbw47vmT0+UW0aXJCv153MjtAEmK29ihH05z4nqNyswPGSSP20/4hz4lFKhRdu5lV9hYWx/M
lXipSZJIcBf19wi9z/pxkl4Y2n/nIARXk7lVW2EKXEnybrXa+Kcg5a3jUSqldVtPt0gm0HhIaJNc
lSJTEcCZ6VUN2V7KvlJVutHDxGkSNTdKsDV7IFL0B5QY2jVrwpJN/lXVbne9Km18NfhNMjN8CVc3
v+PYrW7r/4VPtBN6U2wgyqBS0osdJwE/O/HYp77XR+HRBDbMmKYW9xxbXnNmnQF/KWb2OYKuXcuA
MnO3jHySQnwMohI48Z0dyiuAc5fzaCh91Vj92B0WoU1R05VivyrFxkj+gjkRsxW81blTYRHkR+a0
wYmZjRK/9q9Q6vnhOxbStr+dAcFE9Z67uhR9KDvwu7mNP7LEN4P63vGQnswAHix/6ESBWXcNkvLo
X7fPLu2MX3DjnDFT8gdGKQu1w7DWpk65mK7H5piZMuEPRVFyzRpsPr01K8alVphArVZCDsmNWcpW
TtahiYkajyrWizUBkg3RC2xfm6hL77k98MKn4/+XEkYVvMmX3UgI2GmveqQNHHs1ciwCp7yYn7g9
/JFzWBU0F+mPt/ETaDx5yvPonVEPjBGf4/Cp/rn3pbFdcjf1xWAp0zTCbb10+To1ilu+kMQ6RY7z
eVGDqPP0PXoyjf6KBSEZfYvTf3PQBW6qDZhBa1JAJiklh6gYuq/vJcgg+Gxhfqi5Al46VhhXRwvi
5OYJ2ozaTk2SUxSwk0zKffxWXGOEMbnqDk+BUsj1emNDDeP4S3krkAk4XxDqkBSVwIz0Q0b5EP5D
UIarc8mMDSg1zJy1SAYAa0B/dvZDnYygD9gGZsscCsWnrKP5KC6xRe0PX1f4fU4unyfbXB0bO7UQ
4XEwP9atlL0h9VujUZ4R2BVm8vFPCyLhppPnU3VMimLV68MYz6pPTAH5+h6FCS8D4UvXke0bPpGS
eCnS3cjz9HazsCVqitMFArTmM7vOlkjBTCn+A1/G3BU++8VstEzkSnSzbBpToVTvRM4menyvVVcY
KJwgcbyum+VBPv2yDA33NPjzx+hpidJzBb2bisOA7h9oqJjgPE1/5/NqHIdSWkJNgrNr+jm4YRRq
vcBz3donnaL1j9+0jdT7sHGYNnfDE7bCKFvk2H5OfPWdPZZdNyFgFmi5Ot/Fbt26Or5W37Z9f37H
19hvWLy7/bu9dRWi8iiNND/Nv8xzSjyMWeKQKosV5DvPkWMTMH8DhDWeb+ggdTN0EQFdEiyZqQDP
honfFxjHeYuLHG0tzADakJ9F9p5+HKQu6Kz5os5nD4XxWxnUVxjbkLfvJqtNPNt00Bsz78sG4/Ln
yD47ZfC3SMi2/CF/tvGBwq2mkH3HqdVGauSFsXSdGW905dY1aW4m526ze5l+6JQXJPEeHveyCINp
ES8txZ2NkLj9ZZzq2HMfbGlVQbPjvOYA7kmUbhowGFbYHzoEXsYdAFnvCObl5ilaPZGnbeHqvT+v
knRJ0ACdEgFgpnAg/Wz/c72gHzi23EzaiGtznxfHZnv6HUdu0cgunjnpdboYFukG5imX1tiVIujF
kt/LgRvaLF5fXByI4cF8uQmm4ck22eki4nOiQ2TnU0H3QOCPXnb2F2fXfwBcM9k9uvQ25eftvkOU
awLkSo3zsSvv5H1dVEGo115L9LSaSJet07+mEKMB665vU3Rnarg6h8Y382uAtmrzo92tnu1HnmVZ
AvmfKYh7caXyVRaOkTYi5vGDav/rGotSu6HRynhhtPfJgvmU8N3Vj+odMPLKGmndbu/WVeqpOQYx
VQNsBwSALYlHYFKfZZ2W0XIPPbmQQdwChdPWW94V1HWbKtcoNzhKlSHGW03d0IbG4oC34mAQXzZ7
ZChl5tbWG+plLLeG/pifSMw4zLYRnCj4u6ASp+iH8XtNI1CnrZnNYUvt6eg01D+ayS/Smwp0m4gs
RDHZua2ji9cEJdBx7cplZrwwJiFGl7F2AdUy4h164QRhhKJcQGNkoGKAWC8iDLAMLsKxR48PtPh3
R0/57ZldGjTMBriNQPKK4jweUXQBobOkNb0Y7wnsaPIelaOURDls+hx+87Z3zf77+U+NmUt8buyT
UqfIDP00754sm8fDbQlhUx0nhS38MJYrg6l3DMU+Fdci5knJwZvI1AOFFnOTa2vmBfBaCnk27+Rc
I5haFotZELVFXQV1lOn7vJ6TBcyinYTSqK0usA9dbzxKgwFEWfTtnKSUpHpFOq0BkdQqyLh4jDqQ
D2bdTXvNVAiAvulgBz92WICpyJcXAFuA/59RzFhq172X2VbiG5K7QQFo5P3OYLTBj3Pw3N/g1h7X
RMy5RJVPDyF9T58v9f9/xOXUo88nE/1eGPRrpQ+ccYYmNN/cEMMy+cfGxLkhRxHqouExmn1xrFfW
7DuXp4Uad1RQVUM8SeVF+u9IHoKk/5YCuBrbzBPPvBC6wqAuOaIFY6vmtkfSEQj5DwMaAerCiQ4L
c0YwU4gNgQOTub8AMl2e1xKvuj1ilveMF4t/BSIzHbWr+eWiNzxctjKxnjDqk63ffQeRWo2XJc4h
5ksvlsXtqYs0rlMIBIgxW5ZGJ4DjE39+Pu16eTHsInS+gMruYKkgLhfDAb0RXdJzUrp+2mmnj28p
QTSIVBocND12/OnUtgoQabBPhT24snxc6OTxYwtI/aOE0EuKK1jE99OgWzB+4Y6DShxo5G1PM2ky
gPuCp4iflKnREwAfhM0AW3YB14SY2mOBoFAF6WAiyGdwk2hWbxBAoxBNcli29n1t43hmqhC7jOqs
4B0gC85AH74KOU6c6QLmnz2ROJgDWCqi1SJnri2OImxwet+PKTgGP0JTnvHborLYqdzvvUvTlpQP
ukoeqqbpDF1gf9uhRzNXqah03iJRcCbd6Eyu/Gc52pVU9ZNJHxxoF5yzI7YlpC9yPm5B2nvC1S7F
zC9cYlkNwcyUH1Swj6UY4z6x5Q4uIRSo+QAySKE/WFICa7NH1Axgl8lCEiuHC+UlGjln+IEspPw4
7CTNDCeh5Rm4QOMiBr6jVHRJi7qrHdDi/2n0yCXOozc4zIT8iQRS/XnccrgxFKdWnYfbXpoG6FGW
asUtjGLxsO//NDuSVkGJaTZ3RyLUPbzRIl1pKkltX0eeTuxzStqJyL1Tzy2rV7CsWzB/0BuBtTqU
9dfEofM/eHa/wEi2Vjx5tCmfZQ2UGTubgTuL1Smf+wIooMuK1UTuTjz+8+Qe0gt65rYvN82rxHBv
oEa9rF0uhNAqR6Hfg/DQ85QHMctTTCLX/+4SMUY6RUtLuhazsGXNFnp8eKteexcd2DyS0YXNF4vb
AmLMSEBjvNPqCYhXvHbEOWpWfztiTXca46gQ2jnTtP7VVueETxwQ+cYwYn909ZL3mGRgUwHBujsb
OgFdRPhK48eYPkrCIkY1Tb8FhQOecbPoGHuQo+5iqKAgkFF9y/Dq/40I12EnSnxYNs4DGW7avLfp
j3/0uT5m/ZnJYiHwUr6+w8F47sSHvE5j6sdhxWgijt+eWqvcxYDt5xRVESeKxvWdyqkhK0gk3xHr
6rOTmhO2KbA45J4pJ3pqEIMeRXLlpYzrvnfF0o4sPy1hwLlcjYnV2mrE7bpDt06aVBtd/plFxF91
ZnbrWWByXTCiTKxGn95OaJdb1n2dVwV0AN8nl+PN3QY9IsUCcb7cD2ncDFkOu0APgl5io30dHgCL
Fjw3QRvZTBX2SQ43buu4bRKEuswm3hAxAFeqcJVzKGeRTwhUW5FNA7wo0tXgDUAOBVKj1MkdHuUV
G7EeAy9kExMG7VHSjh8v5Vli+hqVvhT7IpUqeJJilzkXs2hbYrADwdV65mFO2iwxyBNTYOQ4zOP2
5j4CR6qwpyDBKplSWdy5fMzRx2ThqcamfRg5+L41aPSrFo2FgvChnuIPSCn0Q4FGvN2VZWvA/1mE
SVH9DcUbiIzfAuchwZ7FFdrf/L3vsGimB4yL6fC5snB6Qn1i0PtqA3pvmNQH7XZs7SqCaK4nBneB
bVzE3nmVf7iCKIgtnYkTX9JXpZACb9OwcCdJE5cfYt5QLTSXjL3qDEH1qCZHjaLzunowCDKkW1QG
fjkjX1Ew0/t7UKtatPw2dHNEb0lCm5eS8Eb/wRMvJeqFrhsO6BArn629aXtPeZ2icMp35u3y/3Qs
VvEdjs37adwnT0BJhIpKFS8QwTQAC+iPq9RDZYWHzzA92evuyL2KUyAQO5JtKcI++ddK5b8amgYw
6gJuQfIvq1AyfNz4WkjKWh2+Tnn25cRwl2V7GTuqHWbKPw5KSWAjNPCGHFVRNXDyZfk935S1YpYs
rhOk7M8KvHeK5l0iv88/PIp8Q1jPgZFkmhy6csixLwdGzEAA6ycfXVbKrO+IBZA0P1+pkLC3a5mR
8PA6+8kaAHgqfo/nJ08GZdlRdJ4U8B+K9w9K0Y8sOR6Lr0YTe1HV31dYOL3KASpliZGQ1Jez00/q
oaszoaNNNikDrcqhB777WfnFrTlPh2inr23mhE0LroTNhpEE6cfHJEUDLOYsvCBeGk/vvb2jEEpx
LQv9mEHDSuvMhF4kFDvtWUK3Dgf+cX2TQPCBDe+a6p5iQ0zHtTvwv5hokSAmGh+Ha+f8FyP9fX6Y
I+g+FWLAOWsk3yOOyfO5G6OBRDKs92Xi3+e9BGFYSLsImRJiVJdfjzMguPa4aZZfrf0OaiuFsagd
2fGuRnF5L11F9an7LTuKVMD5LLTpBvIeM3nVKwOE4dcPE6wbYAtPOxWWyB+BV14o0qdAC7XbBJ4r
v9hzQVb0hwejwzSbziuIzdPTjyfKbRrBe7DnrNFiXL9soUqgtk3WU+/VFdxmwwrkgz3qPLJlqFHQ
xEGP9pThYLJPO2zF4G/9sDdFdnbrHSr9MmaADmVd1svsUd3NabLh2n3hWZCKQ3m0ZNA2EBLGx1kr
S7RCYTJC0YmrzwFYr/EOH6VOTWctI5naRPI3dLO3017Ce7+RXb5B2E9ou0K29fyb7ZgAtTiiB9ei
bQ8iQLFGIfbLGYS2rZkFnTnUruvmR+EGHbr2NGiFxA9CHskDht5i701+B40dV0ZO4YZbcJAVJDZX
a0K1YDZoJKd44/C0dWWyLuFY/pzTcBnR4i41srROZ/mEF7Icpwe2rvDRSJxETj2/JLWpIgA0IFvY
JCW3KWSH0FyM1UxMw07eNMyrrg/JvX2eTc+RyGYrsWxydGma+SVFn96OrkVi971XnW00eTz1AzKY
PbYjzjxlK6GoUG3k9eOsv5Ri4YW6/rk+EcERp8ZVsxGhOqBQxUEws2SpC32pOgnxuDZ20K+EU5RM
TbJdjAwzPxtXMfh4n+2uwkK8yNgs+ptk3AccyrDQP44nTosYEudv0kidvgUL7KB5MDH0H55WrGjy
bbmJfCHoQ8uVH3p6uk7MlKa8EH/rSZCO1lixXW4xZ3jqo0zBn9h05rJ0yWsSOKMhD5AP92WRdxgA
sO1CmQ9NIWoj/Pp5w3R9rNAtoBZmoLDcl706jNuf88W8Kvk9Y2NBAMDB4D9I2aujZA8HxberP2my
x/tpIMyVtuuUv2RDyVHUqAWNpFwQgzax66PfmSHrf1FFZ2Gf3g2//zeY9hEtAGohpefEQBh4LW2L
GaM+rxn4vKKPz+uwXK/ZCy22X/Q//JWJNoZ+8SG15Vhk82OBkRjYQUkt053uzI1y/FpHXlKbIP2F
RFw5Z6S/xJdNs9E1Tu6LKsKzk0YKgXtT7fZ8ttBAApvE0i6TDAzvHN7I8UXU3rFBKbOy8CB5bhmU
F5BEe0azEyjAw6tcr8cCPDoqMyTzag4/3VSpznoDVwXGG26W4x6U/scrp1jp0aa+M6LJ/0bJJygp
AFewVRtnTsPN/R/9KwpaQruTJmxuHkqCQxybGRso0OplIc0zLeZO7FtfU0Y11VP6VRhQr2BE2KU+
+JlwvQO8S65h9mUSCygT+Np7dGvFGIvlhQZIfPy5xrnA66/7IPJN5gOF9ff/arkcP+9sXNHTp2Kh
Ez/Y1cKtEmFyli3OxMPWZtW/7DZEfyzjkngfmwEUAZij9z0BP1daxW2zLJYE5kI0dBhguz5xTfn+
cELEfBk2Tey7I0yfB8wXY446AOsT4BzxpDQtofKpch3LBlsHcM/Mow+9+9H806dyNNDlTgZ11Usk
ot3OUDnS9LpNInZqkzK/xXaInYvgZoorsQYkPC+eofzzzI1TTNjPatAQHl3RF8z5gkjnh663t+I2
M3yUPrgcPXS/HbSaibJ/nus1hl52rUBh6cg39ttdr3Frvp/GpjMsN+X5MCzmDhwH74qNZ1S21o5N
OX67GtjXEf+csLbSqaJf0PqCxuA0n2F+VFUGp6EFJhIr4HwvTjxGdPh3bC2qfZXjycAHLhqN57kM
Ob25jYJByDVewcNDiNyFrniPgXzTEiTDqpqKZVFd2zT8ounNpZKSbgNbrjv1QxZRvGmF05iViasi
+d3nriSQ6pbe08griYuEz2axx90it3rj7K+AnDHJ5tTea7SCRDFWIN/5SIbOAvh7vPyFauWk8mVu
KMEaBDRwxghhbfZfZ1SgpgN5sOk7PbiaKHhVMDIGNC5YG6pcW3VEdrMUQu+QlkyqNlFwZ5Gi4Rhp
TDNG2GXIaujH/6luNjr2bfQIVHcbzH/UeQSHxFMEBap+FAqpr7RUrbbCKlhCMOreOndNgNqFVEvw
bYMJCO/p8Z2LeMVhpIUpE0RzLjH+tIFBC2F/krAr/iOyrg28CFk8wxhu/YPSgjkPirXtiYlgL4dx
lhfwPkanmuO154dPXpR6EjuEjLNOX/QwBFsf4oO2bcWlizAGAuspW1n0b/G9xiclpb1gp28g0pMg
7mun6nSR8JjhO7blp496y/ILFmswNpZdujVFB52UyWWvVSHxEv48ZVjvL1R1R2obgymfe8LW9WSN
JNg5uQu4iPOU7IyBOFXxProAq60DIsj5vdn9AHlq5XKEW3WFu8uC+QFVPtdZhv3o18xtZQ4Qn7C7
p9j2wNRIokcE7XDi+rGRZMeoe88XcCGauYbo8OhlW5oU9t4Mixi/sycrHzKyHIR5iIj6Gp9DHWPB
7buw0NvjndXGPMuEP8zCmkSN1eTrEFiHyJK3OUifO7py2KVbtb7134iyXjnrLLBCTSvmnpTU8TgZ
tRC/q2tCQKoTVDoPBHq83NjsJXvUFk8gqVmHk4H1eIxgH0amlTIm+WVM4LFN/0hV3ckL33UB2mcc
sqtTy4kWNa81IfWOt5fxWCTfeddTvpQog7zDawGLCJT5W90c9eZ9j6ZmplwXpc5jW8LFR3kuT0VG
3CjVuF0wRFsRCY8wn0P+OCteRQenA2W/bcfgV3QzW1fWwQUSHyup4V7sOmRzQukq3X1N2y5vjVHi
091eQdFJUVcDmnsZW4d23GYG8op3ss36RQyNF9GWujW1tTPUZKEUfbGiHbcZCUzgP1i48CzUBu4D
M6XM6w1+1EyRVHDnuSma0Xz7ACOEq/z7ifSSDl04xyBTAeJpsyEonio+8WhGfIGJTz0tWJtbAO6b
EAFk+aBa4eEowioYDy+J3COgS9Auyu189YBBBBZcUBwkCM53T4o5WMxWqPEAaO//qwmTPW3COPPb
4eEYOzbq8yEfP4gvHcwWm5IKrb1PerH6++5cB/dm+q44KUYi0YuX4rpZSFvfTFJ6FiFvnJj/5rMc
4Lq9pwInvMKPYIobGijPoRU1L9BaaqMmGgWFETEagRvZumwyRCq0uk8C1F1uNElGR0x22R4fpc2M
61sreg5oBLUFq7HPZm1PBJr2/ai396NXPMTKMBdk8me/ziXieUdGX/YKWoOxCMZtgz/3kxF+NPY+
G9o+hHonsnE6QcqvdoQ29LhtIDmuQ8+IKvOX+NJYqRV4BpUU546iH0q10doX8g53CqoDLlE13cdK
AD1aUc6D7LsQQ1cCsu/La1bFyAI9ixxajrFBifb/SeyGTAfhO/9+OoEC1w9+M/OGcXGHWNx/58Ir
oB144TvbsE/o/lc2rC9kGsWzlg6e+wTWxACkI4K7HRTK54awKx1vWs+qADHKot7BzSkIJ9Gn6xyC
g06SHR5uNWVSrWdTnViQ+f4QHyah8M65sYaURGhwmtIm7Q6sXKkEpzWLMkYfWYYGUOn9cjrY+JzR
kQ0EpRldj2lEw1CqRpEse+/ZpjVuB0BRrT8QrTC2Y+4j/xZRSBaNwSXxqlub3I6K+TXA3HW+xj1n
8flAXcw5OTEWcZFv2XgFt7dFpLG43QN18pQ9TkrL2Is957pslRsgPk5rOGBo/6HAEfvQmuGMQqu5
NfIdnS93yzEwkHsdpqXJX4j3n4+54U/YAdF6xVVe6hgXjIsrXY1QQRlikFqa9cGNlZt0+CEgoE/R
H/1ME7Gh2tmuviKwesfxVsCUQBUna2toEXgQZB0iABt+aX/qrpWhxJYuU2NOdGZs+LezLMvDjq/H
NNFZwxm20Fcnpy5xXwxXua5pmOI3rrDJOItaWyyaEYg+b+ljJdIJrHKOQ75mGCJrx96GAP4V3fM4
MbpRDC32cimXN7DefIGzYQrCsBAUSp+PNRGYnA9YvH0PL/Fo4e+BomMQGMpJDZHHxep6sqLs9fO5
13h5jv9yWSbUYeVlvUoTC2r+2AdiqYH3sRcLl7+++bZOJrO1/YLPS2ITgrgZp4opLUyjc8Aj6X40
VFXaNPerl0LJB8v7GvhchO2rSDc+dQRlzxoR+hFU6JDcihUC+Atqx1v3NoSaGJxNYGxFRR9z4ICh
go+ZdEowf259GdHXgviWNTrUVPupIO/NnzgRbjkqUjGS3QsblbII10ih2u0pyHq3ezjU7Q/PjNmQ
qSy3FJ6yfosANEE8zXddbvxkxo5osJKlgkHOwebAs79n8MsXUrC5U9SIRQIc94+VHZBrZJydg32W
T1ivNEYv0VkJD0VrfLdPMTVQoeZITETXbOarXTrWFH59CDugdU5E17T19SSU+0xxewso55jI+ZCo
nQFDWNsqIeXMKhQRqAQWXeru+PfIC3OgIUIc7RJPDFYRZ6hoVvBHhzALmFHqZIHzFW/3N8NGWlA5
L3yb6wbn8eublHQNB+/7jZYk+K25ASG7naDdy6uXgnQWpjUwiOO9x85rfHBV5/HjAQxzINtCsEF1
ZRtk7lFtiJQRVTE5XqKv+4xi48kmsmTzMClDT5ivCt4ZDKO6DnOvx9vL76jfHDNznadtHTWADJTI
d/QO8nkDksRrj7U1sfEsWV/nUndqjzGJl8MtW0A5KSFMAWleTe5L2wCWlwFsUjVbRsF1LiDCsW+j
4ur5uublGuiSZkqNKR0SEBvUoGtej/hEE/ACrDzd47co3fvt2ApJsqXq9Cmyk+4nFqPC6lE+xGcM
0seL4kq1wbwCFwVcGxkwqLmp5Cr9oWPCX6Rqd2rQtBxVXvcADA0BhkN0y8pnqSJNCTaBoB5r+IGR
x5Ld+uQOlicCi2B5W4IbZxsyhs1Tua9EkVYgYPAKTBGI/6M29tiAXmjjZ2qQ6/vq4/9x+MF240MI
hJyvujV75mz5ULI81MhqVjBYX8c3wJFI3M56ur4+FLfJzapQGSlSBl5pmkXbg0bTpizo+zNm1h58
CsOfT+ohoVI7sXI46ylnKd7Uk5WG947vdBr/Bns1uVqVgGruxUgTofKjwGR8qTOvai4UTtJNqwMj
zaXXcf/Mw4bKXJUbn902Im1SLA9FBDQRs2nVBD2AIWr+wZvjqa3+nUsx5CwUNgJ8hbzVbm/6MpmW
MK46IRwFW1+TwA74fuZmMQpH3NNHJV4eqAGDE39zha1rvzahbFA1zA2R7Is8FWHsVu9vvulURxFc
71bGt7XPfkeGPltHTmD4kHNfVcm6R4Ew492GGkDSWmhm7NOz5NeVWyXEq8R09SGDXxs3hMgmfo9o
BUh8XpK87T3+PJvFNrn3jTtcC/ULm/oOqieKp8d7AUUoGJ0Y+TaAncu6I9uyGfB9AXxCwCIg4Xpj
7TiwSljO398qeIZmxentR7aHg2iGJFTnHiAy+jlLcYNr7Zc0CIPh/8wBR+AX1UNCXJtWsMayDGnx
K7mSUQzL9lyc10tpnV5BZYLpb+nxfyfeExwPbn3f5+k1r957y3446TAsMD4n/DZPUGZu7Gh5duKP
3WayV6+LuF2VnzwH1o0XP/EUMfCkIUzk178a9OgZ2kzh5/5LObJN2OrVlDcfrOV6bp51H5TBKkSD
s3lKQWJ7BIBl4Ju5USZA17U4gaAFaSMMqkJIuXfTHV4rB5Gumq2iuIfKBH0UAWZDtse68wUFSq4x
Bob5ucFzilmdhaR3MMz+ITfE1bkq6s1+XtjCklm104BjXsSY3KY61AEKM6YPoq5WjAa0VVUQ/VeG
R6NeehD0qVIMD/lCmpBVLJRpCCb0/8GvqYb7gmx1YfbFsCkTfqeY8WKcKFPJX1WT/9I4ngAqQiqK
teyIsvrftd0kSoSou/nz8/yDlBLkdemMoJwWYVS094luxTX5FXptI9IPlI0MfWOXLx4SJJHunMQe
6uNjySPwkED08hedciRviweUAOR1jAIKAsLZ90Bwdc97x3DS31pYt8HTzUGS+IcstKTkcOFICH6f
Kj+18qNNE7lGmjfqRAMdXUYIyEZvFm2L4blVs8+yyQGvknhn5mj7w55004dQsKKZzu1/kBbz+Kr4
etze+XMtqGI39IKDFL7CQYOZqGex6bhh41cGh+glpCHjs06d8Ynl0h+EQbizhlVUUZ3tXcj1Bi8P
Ebp8PCwSzqvOot/UX1TsXzsR3fo4pWRnYyp5hqg2obIiv9IRdaIxCcNHZ0Tum+/EUzHQd2Uph76G
bWOnugzT8x1MaPQOdxqZ3DDihI/eRJZbPvJ9u53+4Sc5wTD0P5fJHt/8R9WLqomNjU71l9wpO3Qa
+xOck5M3QxMIqyHPGk8XHApZPJxLJFeLYNd8Yxex+JxYjqhT4b+K/XhMDS4bzTrZnIylnaipjI5j
H0aP0pU1VAI0tPrjg2x8+gC8DkiZiqD/kbV0t+fJatrAhU7YpN0jFO2I/GeRPy7Fq7yafzNDUg2Z
pRfESRJO3m+PKHA8S/Yo3ezXws7A9pf4M5sQqJ5ekB63wrLk7P//suqirnHxPDnMiy3DePz1SWQ9
SJyzeN4mz6wCPR8QQhPkLsEh+FuXPxR0OLuCfbktu7FPj46e6p8bVGeJPtvuqfBnl1MRVVe2auuw
AkIs4SciWmj72QdDPPxKRJ7GuBf3qApjkJmA2RZb2dTsGxNs7EGUBa0m4RUhs2FUc6Q8/hz3NfTK
JqpRlf1l9n8Rgi1Tl0r87CrXOmvhM3qWccoQ5z/ouv7CuRkGlpf6pNLCtgAmqyA0Cig2FCJ0rogi
7DtwZg/Uyq38iuELSCuaTkyeZkyV5RseHPOwO5VyGwS5Jw1BmbBl1uRA9yolYio8hPoNqutkzfO9
0y/LImE/DeDW/ZzBo/pnbEpgGpgrpF/msyvWu9gmyBoIGdMke+H/EIdyiqmm1nPeswiyNkBBL2D9
qPxc7mrLKGIgW/yUwCSZ7nwxZKBovz6vYy70f1wTcL0/7rG9roogd+blbZMbRjvj3Agig0+31hF2
1QCCxN+jaEHUvq9nzujLInXRTDtPBFuHPTGV+G7Zqin20cM2WuHIA+mxu/TGpPvCSIh6+QVqdk5A
av2d+U4o6DokMM6zb75WLEMXXst0bmhgJ+Zn/n2ceG2jq+1rkiLfL/f83euhNPTIAj71wexf6hVY
MF8kkk8oGAv1Bmlyjsr2jN8s+Vp3UTjs4o1x+V7HshyfMxAZ3ttn3tp5LUFZegwRpOdji7KBIBgc
UNoROQ3grBUzbRGlSWOQzruiTQvSnU2crQhLgDgJdntCkzLuI68v01GQQoL8r1+tNVf/GWlxDCq6
JhiK3991IXGyzWdEZrLD6SWs1HYvGhoNYwlXzNH8fauCXPSGU1lkido5QGFdiurZs9YGTDBasHZm
4GrwaTFcbCnL0ZoJ3SHMouPC6C1YsYH1wk8sKHInzhB0oE/45quI84xGRK7uI6KShfpRbtULEmqj
5tOSdx0ywcGlTgTY0UZ5ZiaBblmQpW7HPEeEaXNq5hGOdyoukFvF8FIveKnt9TgD25WgzUiKxvq7
46IqTxLCx5W62wkjN1rZjXD+dGNyTrWXIAuPRaOtZ9TO4KffLA0pIv0OB4xYCkPlCA/FF0mHEqKF
/XhJAQI0wsN7kXVUE4xltX+0qX15fRYsWIuFLmHxHKE5E6d6m7Y7b5O5wlJT4ra02iZG2flW2cy8
iNkCKso8WFBh2zcAtqCTUstFWnQZHELqNfULxaMpz6Q+7SO2YNTLSHFeWjfhEpM5qu8O+tJUZfXx
FXeeWJ2l4yADoq/QegpsygmGuA1te/w0FcOmzWXxOSfXReq3eV22+rY3nTJpJefzB0hNU2QmnpT8
z6d4TuU+fUv6/wQ6GHo8DPgoyT5fE1iP8hs6BY7L6UBt9H5eFiy+Aii76bZQO/mwN6Tc2Eb1Nkon
+df2cYbdrkh/cCf7EHUla6qvyXJv74KgqNIiufY+y4bVV2CGCgim9B0cXtxxo58w7q5iKFZ+hQ3o
LVGVUHHa+AjFVJMhAdn6Vh2E+aK2jyhGO4vBoyC7aZjbHQFMfwDN+Xp10kuLn49t4ZvilMoNYYJw
1ZX8FQTf3+d+N1LRyJfoqrdsa1vDUY7kksFVoryARenc2FFOX/0TC60bUanYGOAr2bDFBzM+reO4
+owuHnNOl8sGQRIYuY+52Cscx+S0CP+kp5LBQR4NGiCDsgVHDxOUfh/XttIcvgoAsdSSPTIeLQjU
Aa6kSIJ9Xtuu7pdB+WIgnyTVlgyvqHsQXpYmuIK/t5dZOOAZQxQ8nHZdAfaMKzI/KxSYuRU7DvGW
YDBsV3byujdI//vIDD0unrpSzDplGNY97ebC6/sqTS1NglvjHXI2UM7dF35uaaIZbPyvJuD1lCef
PBMrMca43BTTdocog0cyFIB3aa3/r9dXvwSdqzNmwb0nFvzUANIGXv++UJJr4jwGvTVQR1jlOrCz
bjSM4W/ZwGnwyMD2HENqeK+6EjNnfihD04xrhPJm0Tz78pbgmlGSJU6+FUyFqK3JlEY3Zer3ac+z
25eGu4Nl01vFxCb931Ze35S1J+QIgoPmR4vrJTPxfiJBF/LRntkJJjrYFbj0dS8v8yp/40yIcBm5
5PPpeRhL8EjO5QoI2j8MDEauRpzvZNWdDRTlGkvbLi9PzvMa8eWSgL3gXJdCAjks2JghrlIer7cN
epmYJPcMxN9AUP2dlLj7OrjPO7Gp/r6w/f/ZcartpPh5Pl/eKHq9oGmeI9cj68shA5mphbO5auXb
CdovapJX+pZ3VzBy/hQh7B+DSJptMo28fy0ZAmR9tJWHXiJAYVkjxZR1eWrGZi6Y1unlP3IxiDmw
18BmE1D8aOD7GqTeRbQ6Gyry7Z1oTgMeY+y1/aPTj5KPOboJS6HMWkMvBIdnx5zVeWLGwbv1r5ba
0TSsQ28ZWVcTexnrL2S4klOvFcmDO9Cc0P8t79WSrBwq7IoiYAZoBRGNpBxYpA8H6bL1CAwGKagJ
jUCMKsvQ3BY+1OFsk7Sionqh+IGxr2o2bFWvWGrBhpb3PjS2Zuj31YUPayqXvccuoPQfDUHsQp3h
ZXO8BvYWRtYwpFrkKhmu0EeA5CEe+walXFIW+UEkQIPRRaQ6uUvb2q68ueYtuRY8zHbsuVAaOQvq
Xlyr0QAMuhclz/AgPqH5cI+V274dxR20IhLJo8jKt7bIfMpl2T8y/wJYG9cbwRu2I+dilgf4RguI
MnZ0ArKLDwpXkx943W54hxmM9j+u5/BXnOU1Akg4nZQMSKmqlICT1tLC/m+XX7Ec0HsgHG+cDYIH
oR5hXX5vso2XrwaUGyfrO5CQcNS9go7jc54K23tDLNcmqgf9878AwRmVpQfv4umgZtGTRlpOn4Rn
U0VxgmErdA+JwsbTPA+38Ea1q44EWPJtrVqSmFf5eDf9NxW7BfcCAgjr+AjlpRpzVPKoQRo0jix5
c9QQ1UdPPyufGAQTORvdpN/Lca0lZM4UGvTuzkmO8a6gasWJ/BsYnFbTQ2X3umJBGp1aP2lmUP+U
DMzxYjbqzLR0Nk7yeooiN72/RC1y8SC/aK08naZs921I4QTNg9mO9ryRfoi9hkkPuyNqHLWpacoG
24sSfS9XA4sRSsZKOxm+8qycAsz/eqjFkwzRw3dxGr4lsTvqUmXHAu25tvUiSfvfSydlaPqhSwns
Q6yUpYGBhfHBIh1ySxkhXy4iGfn707JW06fspq/71ccarwsbmLAgkJVtkmJh/v2wRLLDuCCb1ZOH
i2gmtqEfu4qciWk5IpLTRrjplmZ5VuVfjlaEI83IHlTkXygopZZ2x/mdMlW1e/VxnoMWeSI6KiJb
xpxh2sYlIFXr5W4ph3xMZHQz9v6mXBaq5PU0XKapRJHYCg08nMbXnuEcs7WyutZyJoxw84Rd0136
YMTk8pnumhPxIIVftBO3DQFSaPuturZMfIoIO4kQR9XFFlt6XteUUYyz3QyH6Zfcm/tBfAwfbWes
lmiA5mJQZ/Rd9sTMcgG6tvOml/w3Wo9XyF6l7wutTb5Vrzcew++/I6f+g7NR80vrtAeOpmtPRsPq
ep7EKqvVTcY7aPDFUNXiQG4lz6nm0UGqjGvlIxQstD1SbTnLuKwR1g3eiycTiRLccOR6H6TJB7mM
ZC8kPAjCl9OnWlVFNPzrXSxUWPHnIfjFsO5sfgo0GFt+T3hl9oEbBcfLfWdi3DaqxyNwtJ6m1n1C
SJuIR7m0ts2AA2sP/mkNr3qc8cVwBvZynQh60Ygld9wDLLUAYveCuMkMJlRSdrD40t4dJ+0ia8jo
w1rfLEWSa1Nu9zrWKFL96LTlTQv/ImI14f3AzrB5qkjXWkRivqzdIztzxNaYbjmKK7qceVjgEvAi
a8lnnxIcjsQ9hA55pwwtfm4veIFQDFQnB2LqX7j2+lkjbdyVYM4E0ep8j356IFDlMTDg6oCIpgvc
+l1vuMqMYF3FrYm1MglzuT1NaChWBk7AYdztVGD68mjg6pqF8etP+/oO86RH2QJAP09+obqxi0lR
I+7m4sj50nvuziPXKXFqTopnlUd8RePxn+8eHOnVPEbGAf2dtHrxKFfnmStgfFvXRgaZvXvtp37o
H0Fo9OFNlxTmHbVDdHXxLjHGROxrUc22z78GwEaUDjMktPsyJwSgNDec0cMS6DZ0+WKlx3lrpII2
GYjDT+7GBgKsPJQhYhwGu4AJfRjG8RW/JLzx/9JaYuHefGMLwT8SYFXAT9QrvOZ/qUdtHf4v4oO+
2tARWYAEGYxAZwa/tfk/2ie/9PfKxBOzplriF61z0KOmhdUlILaE5pW6RlXijA8ie5BjjhwZAQ98
XzSOOAhWFTdkbKlHDLKfAe2qAw0GR6yvPixg+J/yZMlz0mH21xOdP8R4rhjMRTdupMQ5ebwmbGXX
dmjQI7eP89ffLMmDgSz11iiShgkZd+WPUrEECjM/jYlApYg4xRDp3QpD9k/hnCtyk2sRfpeB96DZ
2ZmtlvWi2z4IkS+LJj2pQIc5sGpWe/tENebnbKvnxBhB5BkEw0ycVPubVEcV1078DLlgqvqkFE5H
2CeIAYGeS72rEyuziY1Y71PEW5IbRjoaOxduyUUNhVO7YGFhosZ6vPt1v4qbGPU2QorUhXrHeV73
gOo6vrnmijiqi7q6R0s2S3ZplT/otkPVndLn/03zIdNlXrJudZZAroKnOR6PYvEj4IMx+smE+3qT
cblfA/5+bwg/pXTaOO89miR9lZpVzZs04NUvD4AJTg8Jpy3+wpKKSPZLSe2TEKEnihYn/YS/wJ6m
iU0RfWnQYcjmH+AD2yMqCvV80VACScORG6lUa9CyXwPTyQ7BeWBGjeCnNk34GiYyhML4DE3YWU93
miI6NbRvJ85rL96k/ihRr9g2e+OiXqcQdH3s1R3oJ4lb1M3w4/Mu4AmUvqpIzyszeDobje83qmdp
2kBh+FZtK3v30Xg8oyswUEF7TlvVEJbczV/Sf/af+ZixUZGANvO26q6xXlC3ryNM/r3JU3Wu4Aeb
rLiluW10XVf+I9QZra7/JiVelKR0DdReEE5wNGXgg6jxLNiaNoeQCduvghSmXhFK6+wNNtESBa4H
aTPkmNe8Ls982g8iafGtDHftZah469je8eo6HOgkyHcy214g2FvsVoLLjo3M9REduT2ssXXYqKpu
kIWA5fVIEsk2/00bZaUNRyv7sMgPBUkCxPU0LU9yvx5zZfwK44HJoEfw5D3nIyOy7pE/UdTRRkZ9
y4mSSBIXZBe2KMPUry8tDxpFMxB7ATFFTbvw1hfTkvGKKx9hkC8ZdatCVVIfY3ys9WvvUh3RVFcf
vwx1jaXjCJGWAj5rG15wHICF1GfSqk0JoEDD7pujyKJHXgkL0l0q8sMFhv74z0SNB4KjrSmw7Ypx
LUksLZJMq//9miER6Re+42BMJy87u4SEmcxf4nqxmpP5EFZpF/VCI0UoO1UOKp5L8qQ/COcrmapT
0QpYod2VpXAoUifhpKyg7TETIgKHZWX8dtyOTPIGtxjS7UWvj1W9saGSaO/Isjfq36+q/aDy6vY/
qvSoKBGJjOkWN7Jgm0Tios6C45X8PZoF1qzQFe5BmPr8yKHcWje4FK0IpFSpsBALVH15Cu50PFTv
KTY/9wqLQgn8k+cgNobKHpsaD+xeKrQPY0X8/L0JB6mi21dhdpmiv4eRtVkDelJMTmAvgZjda/fd
+LuH2TeXVkB882r8fsrW+ssVp1fh+Pj956HlyT9M29jFjFcy6R5QyFsb/R9gL03Skvksz6QMq8Cg
ImddrAzCUxWGaaV7qgnIqDPDm80vFGFv7yooPmh+onYwQ+NNjbRvOn7hicvhCYzpQzc042ljg/78
hl6JD/nRhXbdT+SCsnX/bL5/b6hMkLPXglwDeLQfv4FBBOXxDmugnZtI4r0CSK9tRE7YIEF5UsTy
1+9O754So/HUyzlYXVfaZhAOxiNxCxOHbRE/P0ojT4OXgSYYRoA97Ras5I2+qtP0PG71pt2WxRlg
cGYtsvoO+1ISVoVSSnjnP1AkCmMzGZce7l8nT3JU9JRWva1KjObAbb/zMLbkB4Z/ggwNbZiWyhs3
orHBB0H185C/pRrjOTyC/Qr6AuoZsQsOxiaqWUJiMz7kZShBQ1/BaUQhnDSCCaR+D1whKUWuSE9j
MbX6r3sqw+roUNDr6fsB/RFJkUsvfAKDEN+5GnBclPcVN1VFlwaTkpZGDfPIJ8rSCpUcnjrgBqiv
7JPXKuHkFdY2K17Al3XABpJvwlgvEdBI8zU37N0YUx1iZFyxO+IL+7afMGmTXoGEr2B3iac6B0+h
yr7GKRe2+gGfk/PcBtVe/rwHE27+PxyuyAkc48WMNOmHAZChNmcuDBYR5IzzudIukm9JdVQsFS3F
UUDxq65FefSh410dmk54/9hfn+ujWl/GPSVj/lF8aa+n+TSe4zkVrJktSXO4j9QFDNXhpDDIW1uZ
tvxHmMsygO1UvcsnSjoiTEqtwfKbYPT29sV70Emrx2qa+65CaI/y1kpt+pkZE8mKpFQ6DmF9fpBe
flG42WZfSI6t5/kwEpjs7CxHX6CZGHQ4nit0x7sJ71pyDqQWM7qiLEuJ9d9R8u4Sn4FDX0NzMmAO
I+NlE+oXfN7q7sf2tZOxbbr/Ox069op0XxYoSNYEuxPyWK3HD4dOmTG3qk6FlMGlXOul0p+hTA7j
+oCUUBI0DbG/7ljoPiYIprgAhQkseJ1BUX3ZOMNegy5iaAZ8TLa/nYFSujiRD2K+ARfHmfHJBe3f
cdVrXwRDKC0eEOUS/ru0PvV/qvju7HuJi9TE1/HYDclkgHEngjykSlA6zS6AuTtEI5ZRmSTa+nWv
BYImOnNKFjGt/BbqEgeVpZx6nbSB6j70kCSI3/ZKHiNwCiwg906VNOhHkCXeoG1Px7KO+nz6Ic8G
5jRSoPWd/aquIhbyALMBewbAX6xYQrcNYpwsW3E5osirBevKPpWATY2BUTE2FrgY8azdB2lMCa98
lMN1V71sPaJUwdmBoj5mW2QCHTejFv+EopPU+seWgYIbAciCeUw2mRWzGrGLp2G1Wt4ZzZkfbH0+
Y4551vIhMhlViD048Pzbl0ERPjyU1Bfl5YHYfMY2fHE4YpotbedPHR66wTGeFmNpX+kudfQoIRLf
dXFOH9ifbJQ07+D+h2fsEKC3wWsQz07z4+HKow4VucGtBDgLzVN+4y1ecpP6XHgxoBTrOgvvCwHh
G+9H45XDqbk6Yy/smhT3lKkT3h/iOBmUVUkl/WntpkMC+MyilatS45OvKLCrVOnEifyO6gWEja4b
TbQ7Xb519sH0lY3m1DFmJGb5FJ4N41DKH15qJhcgIoDtfjDY1jOhvAInooS0Vp3gaIxcExmkLCE9
vS52fjEtMuCyjIGcMtp++kHanui1OjEMKq2mlvzoFQyJcU6D342RI8yRw+yWzjunhM7W4voM7wTL
S5WW+z67Lob+8GNyC1+KA2y3vlXJ5EzO2OhkClk0qLzv0NH88QZNwTnBKjVPxZDQzf9Effc3tFoG
LoSssfexmsQ7Mu567WfKmiQvETcxHXpV+yUMtqHbCp5z95jsMAmGuXoKNxjEv2sUn8/YuCGwygSe
0uYX4yFWZb0U+bq2a0n+rWhbKks3zsmRTooqc0RxQfhsnBXiIaNY54w1f9qoVKUewkjopcHgmO8u
FyPXqjaVHdoo7cZMDHavBOecnchmOLHzkMhWVBJZw25N7oWFgVxJaAn23J8Fs8Bts6X+vqLn9nXF
KWQqrfaqsbnfLpXLbaGZiNScbPTw/9IVQd3T9iwSs4wkxfmzPhTs7G6uxrtURY69s9/G2zqQR0BZ
92maNnQD8NCk034YTsGXzyLuCNAmW1DNNM2bKuFEp4TiN5Kp/nWfAcsyl4M83uhaAOfnGFXMoCES
hhQ55jNRyDgFGz/9NqxAVJvGpLPKOtmqfQm8zS7TDLFdhw7k284rtfb9Egq3z5sko2l9gC1VMDZh
56pHBe3p9BmNPu7fv8EnNlfajfpdMOx8k9zPquxMJvWFeIVpk+QyrZrD2giVaEDVKny8pKBrEE28
7HhaDqNjjKbrwa8lhKwud/py4Wr6YAcFvDA02nhRRxtV3jhlNGXaWh+y2B/n/otXCSCnM85i7iNE
JrT1tXBXd/yxSjqCGV5k45SBDDWN94PpwHsZ3tYAei2iGrXke8Q8FM1PJmEOWBVMl5xwVTYYTQvf
gxzZ1I/SKvF71FcE0c/n6ko2CbdDVSBkEZYemOPHDX2JTOQ2RyWzLwPSzxDZe+y3cCgrCE+hBz0y
bCFJq1LC/AG477F9GTsYe41Nlk81HTvYSI9Bw3rgJbVVIxkmdEe9nsvajNY7UrBlG20fp9LXTSZT
OyRvIDxi5hbgzn/aEdYR1vR7NQp6v5ilMCe95d9SSpY2+qDxOXOX57fK1QSS0WKwxFUcRKPPgNKD
tEQ8yAp4Vy5LN6nBvWf5MSAtm3f3+FMRX3YNYbPfx+rzIEkfm44/mJ1SwqMb2VmuT33N5TM2fcGV
k3ZvNfvl0VOg2ZSbfJNvgVMWSZY87EhBjwXeFB7b7iQDg1OzwUQo5rCn+GLNtL4UTU9Qc00lsDZ2
kCQ8vGf16UOjX9LaBsubNntivvOl7Bzu7cp5tIoJLiIeoNtx2rFayGsQntqLKPhll/o96J1o9Ei4
ol8DGTt5zD3hARdsQu1+2T/2+xd6iEuvwRFEHazM02fMaCFrmRmwmujZIkoFSWDvFjWUgJnfiEpA
//eFG9w8HUCgZSAJFg7MQdHOKYvT/Hdn0MXtkTA9qIFZhwcV1ecLErjUyViCWCEarCz6Ab3WagHn
t4FtZaiidq57q+dLYVmLFfCM6fhscfsBUyWBEKuuzeWUGBTR1zYUQBUc8+vddy0pnry6oB5gDPQP
+sCEkmhLTUZFOs5CoakQ8UgsqFeKExlMUbDtnD/ZbYTZmqBRpxxw+RUM3DD3h29SFj5VqsgFQOeX
mUdpVSDWoAuPbDgHTGok3od+EUDPP82gzty8cCsyQJeko/rv00BrzOIH68nRTd+ZxYUe+eq1cwCZ
izz8rZ16CZYUiJGTjSpv73uYNZ1ptxlhF+2yOv/XfUazrIqiZFgnnOaObq02eZNkBt/Lk/ToqG6o
LWFbVp2jYEKfJyUfG4Au4Us4lRNAZ/CNE2TxX71RLVgIPPtvIyDOEDMj64q5HSCpygEJeXEEmaoq
oiC9zb4prIulvb1+E3584sSHXkx6W/FMKz23YSHYvxqFQpsY9ZNEGSzMJN1B5knRcXAcPTApFCRO
VQPTEjzUxJtU/9yw0g6B29r6JCZ3fbdnaudfVNbxEg/WOlbgTfViCO7SYYegZ2s2lEXg0XmIRzLv
2r4yCkZX/lAwW690FjeTtxrsuvkJb4ySuE1scKOpb+30yenVc0Mo5ranFrmkLV/UbJ/LP9v0Zftq
GoDUaxGUHkCG/ZDkGYwSYdEf2Y6HCK0HdggoAjg/9PSvF9B9aIvFkHBcD9s4w5YVXOPdYQuL75Vj
2icF0wu5hAC9viPpr3NI5FR5Lf4Ya0xjTpcYSSU10OuhZiwCM8Hnu3/Oq5uIxCH0HZsjkh8XxEcI
efmhYgDwjiauy8dTv2CwWm8Xv3eOBz0/mxM34/LyCXhwuhjufWnn+zGz15rgYcXVRCqq0EV5CC+0
IkQc6A0cXdVHx92sa+vCxX2rG5K/TMpdye0cPKbPwu6v0GZ5pC4X6A1BfrhooNbYcOkHwSgcoxqP
fMgH889QsUGnRZXMdwZqhjjiwV/46Q4mVIR2BYrBF3HkkYuPJpL9yb7ewyMnu//NBeOy5t97W/66
giCuIrsGx0JJGr0kkw2p4rzl04c/X9XjlyOVe1P5UW8Q12W9sKMUmLO6uEZVMEtC2b8tC7GugTnF
m1n8Xg1aSpgmjMhqLStV/UHMnAeQcNHiwpP1Jmb826Zy1Tg17wCxIgDSUzieEEoHJyIcp2r9q5Lb
Y7+qhcxxV4dEffLRWoJG9kMZG3CSnWVHPUlC2VzrUnSXseLhKUcFqlM1DYdJP7wr4cVR112rSDyl
irVBwlLM/bOWksorX6onRlmaxqqoaXvPyyyeljFVz6riL0jBnVuDRlP65Ks9imcRH4K8HKKC1qmq
cjFtmkx762jWa8Mk+qub6lBqyGZuCJNX56A8ti3rT4uNlaph10R0Q+Ckn5rGle1kpoAh4S0fan/M
lcyypYosoe5eYpJBLpC4WohpZqvdzJYAgExR4j43txsZAVdSMk+F31p4mP0u9nzyJ3UpJBY6e0jB
0EQoAnxpXD3lBsZ277y8V9pC1jIXceFiCGmYZeEicmsXfJyezZSM5nGb+JhS+tR92N9gx5MrKFD3
Z/1hsH+K54pxemzgZ3J5QAdXw+Gn0IKWoSIV/cH35CVqi2ZJEVgTrX2MW0f3vpQ0x7R1zfulQ2vQ
ntWy+//sj8D5b4LsjKhllfZ4tgu9JD6p7nsIMnAq0lYFJfAU/QRWdq3UU1aBDLRJ6r0dscxUUDsk
0/QnVmDxKoFcjHA0FH9u98xkvQNn7lUfJc6/rqTNQ5cg5riF8MA4vKm70SI3p2sbRxriPzCzXxPo
7NaJvRYtcc+BSd7drIEqEIOWx9lTJYURt2i8IasyQ0jUhtG48UeKpP3a1dbNEEk9crXYQvpAglnF
MigKQkFcmHJIHAVWRruBAg9fcuwPG3HcTiHkQ2HoUQzh7T0s/ysWMfihtgcxvM9dfCgNC1LoO4RW
5F5wOJY9ThL4cAttFfbcn1vrszgIxv0SuzNUGgxUp2s/RwYzgelqL9550fdMCVcBoZ9qeN/85vU8
aEbT4FxnXXPQ6DCF66zM4X2JomSlDP226ZNgtJmu+HRgj1e8WrPXxkA85ywCAQnlP5bQFm19H9WG
sXoYpfGMyYQA4h8po/And+S6X8BRT6TcuC/UQyOgdgI69rCk6dwUTXuIsJyJMvuJhBuDL/7I59PA
qXauLgwI4DpH6px2MNb1kQPF1X4G4vv+N3lzPaYuqxiqDvkLjVqJ0imZtor5SqncnJYYUTx/Axvf
FwBZ20rkI220reYzGxyUmn0378LtlASm7fuh0nUigj7gcszyEp0W4sNFNidaFkCmaqorAPBGElwd
dZm01AZJ6TM6aIQHeWxboGLU/6Juy/gMqM8UIDrBPVRNIy4Kbp6Gle3+ROuVfpwhin7g9u+i5zCb
ICwYkNFkDw0ADGl7nY36eiqweo1XgUJrAN7c20UKZZXR1ei01rvX7nUL1gQ+IJjbz3qPIlti4Dh5
Z5lu4Ijw1qv3Jq9I8zjgkTmqCbKuWASdP8hPhSMMqrp9CQe/NX1HEd0WMJp9mz60bbrsa01j+l7+
cPH118zX9oJOdNjPZZlK6+PnDv4cD6lW/ne2L75GeCVmVwwfmLA2GSLpkD6iYO1hoS+e0L9VDCMW
xq5uO7exW+AS5QtgEBu83a0tWmCAqGa1gvWoxnUxYhNkicgKW/Jorbehx9z1emPits9SFTuBrU0s
fJHGKV9/AeUWZXowsZIhocF0/RXBQkPoWrEMSFRhrFQ3ufD/hM+Tir4C8Mzz5olY7Avcn98hIvB+
1UKfewrXTtml66bBGgiBMG9sz2cqO47SSiwvGIvm1KEDVQlzi0U1Mq93BYsS0hNq7Uux+7InI8tb
O1I5VJ78C4zc1MyavnqjdDnZJztPzcWGeO/cbnl9G93v4cAQDH6iOKjMEQDz6bpyxcdvU7Dt1Czo
mwDq0rpaNDroK8q8NQCDr8wtzQ/e+ZZ5W05ZSVgwdRi+KO0yrtV14pO1QKhIYOHgdxUWqEKvHvmi
NpZcRXPKImkJwTG7qDyZVjQv0T0GlIlQxizWdfDcVfj7o0diXFIcc+ky8vgTFrfn9e3LjAh3I8MI
+KfJ2ldZw5clme1hFgOG7QcFV5k3L0ffQQIppKkXOxzVo29RaD66Cq6Cj7eOFsjdkb/KCvZl/Lab
CIHzlkVA+AbxOyQMS2VyHpCYAsowgLBZpug0wUIzsMH7/+dZP3Mnzxh18gYJ4Crqtq86t74SoDUO
Mb1BaLNYrJHlhKlncTn4+d+XFHzHLkWhxr7aDVHFM7IZ68Yilh8XDV3Wz+sRXa3+edoGn2i2u7fk
SfX0xa9CBzictjnk9Xta+zobQJ6DVNfiEcebRQFA+wiMj4ABweHqlJlPauIbo9eo3kCSnkJT3uxW
1GwEGk4apoGXL1+YoVEpkXAmGvsmqW+ZNHzx5jbaMjTSHK7dG2+J+FEsvtgwKV06ieA8Snc9T39c
esNe5qXZ8fJC65YHBwSkaxV6dsWhx5lfqaQgsenGIXGgJqPWgN4mxQ/UZSgNC0hTzqp6F5YmwL+D
mbHAEkuQ8b5Spvtby9iUmZxs8c4YXIdmQAX6okF9pdLFNGVKOXN0gfe6ABgtBWHUiIWxzySJpZ2h
1SWMtiFrtx/h6E1LFTnQw/Jqbfxv7SGk+Qs0T1vfXov1itmrdwk+5iyFkTGDAvo+u2cpcgtR002t
fQZvSRDsu9x8tE2Ub5FpyqRIad3pBfvumU0gOAS/b1UK2r/XGCMSQgZYhwoTDftgjbzjc+TvRGty
DSuyKuqYS1YBAJqWZIBI5dl3mtlGYoYpuiLasYeOfaMo81ObJN0J0dknPUs/2YV8cNjKQuxJmMix
Y7k7ClRildkk6j8GkSJwpEF8IICMTL995IVXrn7OkQ164FjJQxlx2KqULvd9ENK/Q9FwXQN+Bnjv
nB5gNsaAa0XK0OdhvVRfZ0CvNH0zj/9h6CaHr3Ag6jnUnLpDSRXicLQdIHHajXbIw+iTXZ2Hfne8
AOlNZZozXJR3wwBAihvpmFZEbKvGnI3yYaM+9wlqT4R+n2k5cCevz7Cs572fDMBYmzSe/gA+/F5V
YeaEsYgI66I3P3d1A3RxooGIb/jwpeldvyhcMjGi6eSwUG9IjXn7Q8aagxbBLKjYcADF1wp0YNnL
mwHcBCO8ML40ws6jwPjOKKdYZp5C3KzquBrPf2NlkTDmwMXeXuXQYb1jHqSvf8fVPTLCRbb8hfOP
caXTzvJiH6anS1y1g/0rEci8PicW+iJLkw6IrcX6XQ8L5d7Kd1Fud7L0m1M2lKQtN2PKLv3tGjBb
SXDkKs+5kOVc795IR3xx72OZl3RPwzGVhg0tzhBXIgb514yH+yaKMFs/tXeMAoZzfTx5Q8Ua7KyB
zHtfNyEq9lD7soTTgL0K2TwMYaYM0USucKg2N6bTrK1KA168+d/WNkenuIK5rg1zkqGQDtYk5Wx0
tGsMVYWrGJCn5YSwkOVZDySuWBDdmObCwy1PdGEVTPL/fili+iH1Ul/UdIcJYZxiJAqKm55Vyfm0
1MEbFXKn7ppmjJomW1W2KsCzge/wEu2zw2fzyHQKWqC7ZsdB5oU6yFdLqXGh5HYuf1N3pjqSwhAY
n8mqP9KBnh3EvTNWIhg1Wi4MuG1s+ZrzMAPPSIBtcL4yNYNkpluLeNWniLiaaoDsOWxY7cpxImat
oLVZjcxj/zZCgJ89jWc19vIZtEeoo8lmkDMEYxymsA7kOfmNFmr6RDbKaDArlCzxS/xqCeL7y3N2
crCd5710cascxHaYYgcDISxbCBo2zljB9aMyVmO0+aNTph969S6LCzWcBby5q9JeH38yz2UgctE+
TTlLDgK8Cfd0tuB6QVJNksXk1p9zLh+DA0FerqUJPIOQgDxBzOxVobL7HOdCFcIPwOvnxvmAqgtv
j+TJX3JCOwS+WnaaOEARFxAdaz2A1B6WbfwC1o8tu4R+3Mv2gWX7hd+ntRO2KRPsJQzkE7G/raMw
qrSk+wVbpEs1Sxod45y1UTU73PxchCv1kNyhcFglDPCEIq0QxfBgnhzRt0Y+F+lQ2+q9erpEHDh9
+2cgA0Z7Yi4a4pJkpYmj3lshGYymwBnXkYQ9Vr7BFvAO2Q/SdBrd+xZbLhQDry83UTKKHgZMxxnL
8grzKcQ8wAOiH/kuKNv5BFVWY6RojCyII/r2qIwS4GsK0pYcjjUZiwK89y6kXkCxzP7bhIhwvw86
bSA95wF8OuPNXUq0BImjITWQ/gkYGpY8+NB3AYVDeuDSWM+fZbb6y0gITICvKKY0Rns1VebDilB8
hldMDdxg2g30j60luJcHBscjbgm54u09jCw3p5/u7w3ikwdW+gx719NWyXzqGnVpDkQVW8TI/3uX
7ur8cOYuPcNmXtJ7PlsO4WizPtvaPXz6srLYe61Avz1NgyjiC6ytFn0lcJjL7nCTstXF/KAl9wsN
NOVwy1ZqAtFiLTnLezIGWMVjJMqed5tA7uDfhG4kXU/9ikwYReEeozAbe3V1iM3W0kUr67KQ+ceE
8RF7HB0XAdsOsBNVOe0rObdeE6IfHf//bZF9VJMlLVnuVRO/zuuWUpPyES2b/X3IRvysZ81m8+R9
bXgFdEKIt5jjfEmgjuwmVdHpY3pGGG9GlJZyNkq6KXYwuDZZCjTAX95CQ5+tVC9+iScqZUpj+E0N
46WACeqLyqNM/3G0S+yMAIHyr29AtTHc6mUnbO4ivFdrrhbvQYkGa2qFRIzFs0RdW+BGeJDnUwOw
QVBJnS9+3SdF9Yl7+bfHEOAK9REmo8OUGJ20k8UBsA3ukK7B3wi92Mw9Qi3fa3xO3aqO5nn61Au/
tinUnBD1htbDLbWiHE6xKV9FyAeAngkxCTTZAfP8hpVKdmvTT3/l+FHaiS0zozyzz31ihPxd/6l/
VPzVjX+YaGR7FA2Fp3PnBdDr65JpvrPbzXpXIkfKHD2VMhh28AJFULvxzrla6dBHxBw6+yRy+u5/
WsKfLlmUDSToGXukG8ReFzBpPgwgeabNL+Q4Pl3ks7VS1jDItgA5l4eQGdiRLRE1GknKKed8kfIU
JrygavPiE+0wl9lMxEsWCC1tMnB3ypbsPPimpyw2L5A0yrguDRztv28WMMrTaNhdlZJNMEgFER8x
QyzxAsCMDZSu64JWBh3xqy/IvIyQShUP2gjn0/BoZayUf9Sm7evKfQIU6/ZtR+HAk3emkGuruyTl
FVG8aYVzIrizsXaVIVaqMFcS2qt0WOBsJoT3+0Z8SSjqFWUCci5LniZizGKb/38RNeSxGugpHSGX
49oMR7aBsHXijtRYdYyILK2rjzWFSnRvlOQ9mYW+MrTw1yKZjTrXG8mPJjHmtcqEr3l70dsbF7Fj
s/jJRDzbpdbxmCpJJDyydQkxjrMNE2SJ+verm9JxltOVSk3dISvVUVKs14FGiLmZgUM82U9omYV4
BgB/tfQcxmZ917+aq35DwHseWOVUxewSxBUvww4SNc+ibhXwr6ZLbkzpYlrVzCl3rb1gbIPJylrW
ncPwFqaYSOqnTJqz9usq0DjKa9xV3Nqq/qLsxG84XmyGnT8S0L0woxZp3wLma5x04EPbXSh799E7
mSsH9yMO1eq7bpxwxqKp6vV5GPTybv7eoGifxDCt6XffrVNqqtH8MUWC45OBy041qVN6UcLX+DrQ
3FsQtnAgHowkpI5gPrxNvYyuUVk7z/W8i95NH/HzvFZA3M/HO0ei5yHY8xGxmRtSm63UcyiGGBZ5
Ls5gzcxZRHQIA1LzKPGsghOIcolk3rf9eccErO94toy4yU63G6AmvsULRW+44mc/7+Qkmdv/tmda
o5evJFoOZKU8HawUg7fGRpV2TJXXbsnsgcuODbxpL8pd5YztUBi/JVXyJjpYw3SgwwDapLn+UBP/
0foqEcWm57mxhauxUZNFxxVhjmyPF1I06DVLHEuvwcvhUQwpZb+ZVbtlJHuMZvNdF0X3D6kbmqbX
/jN1Ya0dmu5+ZS4xCKgKpuXsEUc1e3FyT/c13Ey6utmImmDq3W4xvZXXVoRmW5IOH8OPfxv5cFmO
1MchRnjx6Z8tSP8Lj4eSc9zuOO1yOFb1GDXOVdHkfz7rErNUiDMV8UcPCQxxu9CyUPOFPTmH2V0D
UwGSVRCwZiVdkwXddPzj2smWz2Eu6ZUvKMgklVvSRZLSzARQkA1FjygVrFG7GxLmfEwx8YaUyMMj
2LwGOp7hL/s7Cd5pmGYIZtDYBCGJkRVVWVR5+JyTrsu/fKCm7Gsg+WT8JTVliAJO8Yyf8dFJB2M5
q5a14kJkoyBUxww+alVWKo8vz18TLJ/PCdf7bgWcG6xMhDsYVhqsj9+2mAkjArkzPpHsfXEZkcHo
rviY/Z+TcJtCEDK6ejmREmVdEM4H8mUq6lK0/EoXxtJQMzcrJZ2Pr24U7T6AkbEhxK+MkC4OLu1k
g3ZNfIvKg/+Qa7IgUuCnCczpYktpbT96NCnsivHDpBzjV8eTohxGFf297Sau/3gEDtVj6px9Eh10
v4cJEJMiBBKGrN0Sa0cGOSjBhUiThsQWSFUCV4boGdnNbmmLwt90fVeMMX+fMySroXD+fOR++v6+
4TZ8/MX5DySm0eOHORJWOVKnOT7nm5A848eYJTpzbZO3mR9uuyw+124i84eOZUCVnX3BWHY5l9/M
mgpk0/2RIX10XN/klbd1Q/y4UUQeiDijm+m6CMSKlcpLHfhgVGJk/ZrbTGbObgzf8ynpkpqClfjr
QyC32KEyIkZS0NPczPgw33Y1CLi49acfK6vq//tsNGb9bf6klMW1aZZ+1GKb4Nyp8L41coF8sFjv
QCQmMsP6w8nd4l3hX6x9yT1IAeIX9/7LvoKQRj6bjJw+L+y6dJmp/7Cir3iY8hbk/bW4ITe7c1B/
F58/L7zqmvyvcJ5D5oMq14NKY/1qnCmPJ84Krejf1pVWHN4ooDyLX1DWG6Jrzv4ZXqOdCIZlIu3V
6DGHZorXQ/yaoVuYyodluaSKnwPgJlLCUpPRElqV1yazfauOTCwyVm7ihVJDE9xgdOZ9Ao7ZEuzW
Z6+v1IKhirf9uparPzjZxhYEaRLMWLqUHWRPlDx0G/YEZeukygPg9T6FQoy+gFEVa7HxzBmiqTay
XljylzT+a0wtLT4tPlo+D0Uu16SXn9tgAanYESLbiikj1WfasJtwL5S6OMpEczanUgC0K/nSLwRJ
zhW9Iti8f1X9oJlpauBM+7LWfikrtVKvvChRrBH2M+HaEW9nyO3/yk4oqY8Mdhzf3aJZ8OhI8GMK
CdnKg8AUcmSapqz4F5c0RKxJ8q3b5NB1vxvodPdYSoelVmdRo3lUndA3Lkl7bMO1ZvHaEVWQzzEg
Ifwy37gSfJAkLQ8U2sv9exfQiAWuwAD76fyQ/UkiQJdNchT4Ytz8zlZkVy4fUCYE2ZeMCOu5R+kD
wuMGzLj+3Pda0Ly/KFEyX01Co/Y9kSrneZLlnMPylOxtBsVdrmufALf1R/cZ2rQ9wDnYSHBjDqwi
ScpFB3fZ6zW8H/jULfSn/6InT7a6BJuWbuCok5tbq68yyfgwqvn9RxaDtbBgcxulBhNBF4fxn7RR
sh7BnHO+TVjHNgXdGr/vRRB78eVI6/4AcfTDhBxniSYgxpWQ9kYcGeao9GHQIHgtJ91T5+nzhC4l
NcC8a0qsLseMdJcPzzBuLBrsroj6c3skEWiW9iA+26kQR3yiDGFO3MW+fz1mS3oenzYZVotZT+Mb
jxyvNYD0725+wuGKXdNvxQGLG244DVr3cbRavySc6trNA0zo0mN5DKvNMuccH+Y4MamUPamfKrv+
hONQyth9U4c6rVUS+9Q2hWJuPYWjs8bE+qAD4m6jjjYiZXJ0tFTFuz80Z5R8X3GvLfhBUDGJli5T
+Cqz2siBWYnTNiYy0hQTtzK9V9P1Gzc0KajrW5HfFWbj+MN9MtSYwThWtiCnhbWSntJbvlm6T99T
H5ekrIQeiqwbeK/mhOgANg7dpCEUbMCfT5BRC+Jtxzleh3yY0fPexP3rNghj03b/mN+A7ccDLYED
dBk6LF53hPoHqyiuB6rwuzJUBD9r6EYlVliY1m0/ICkan9z2BrN/ulz2z0A5KRys4h1mVkmT8XGE
5UJiA2N4LKfM4NBoi7nr9zQtH7dceTDtgSRsWWzPBMLT9M/r0YQ9PxpANDCynjghVHz0nqvAoHFf
wOldyDbIaj21HnsKrbfRx87aYyHX5PvPiDCIqEi2RrrhqbHb6iqF/FsmCvfx5fYIs7bjrQsgaOdI
7Z3bABMEkpqcJCErGDAS6gJdaZVPPLsK+NlVAhGrdOK0067rhNNfFj+85aXcyxskSw7BKYjZO9ZQ
ADNWvBA88dJ5MAFRnePHTKFX+V2teu7/VhaYCeJQYxBHwWgawICdgps2/cx2NPSV+Wv+oKChO0tZ
5t+GLihWX6C+RgHB2iN5vmT1O4CJ+qY7CmyCS3krE2BPw+O09vVEZZj4rrIT4FSb+iyp3Zz8UJN7
q4WAWcnUMCJJVHLRXAGusPOFogM3gNr13sLdnH9hmPrU+ZdElMANGPrFQdc4Rb9RO9ei+iyESUj7
MZH5igORndY8sl61FFMGDzuKSTHrdaCehorTkkt0US/X7zDMedbCsgFmNUpbY8V9pMjCtYbStNm9
M6SUOsFnihgwHY6nA14qqY3znG8eQ+rfPvoLHxbYaNUVVXk+NMVIWWqRtRrprv8dNAo0DhPIg4m/
7TsYxsckzvGNJMLciPsfyK8t2Rww+Texag9pGL8m4emXe/XhrRazLLVIzVO4Z7r5l20b+SP0OJmR
zdPr1hIxDwqLWu3NfOJCBkespB3tV8/xuEf52ShEouh62yV6AOreWuepTGJLiUuRKUe5lXAC9ruW
54CIdKYZGaiPOS/lug4UjgpZKVcE3YHjjmXMp+8Q/5z0Ggk3h9+qwD6uSgj21jc7yvrIp6jZ70nc
h04meG2j5xllfz2lTacmDLbbdOWOd2StbzrJ5IlXaZ9zQkVBRq01/62erXKLroqTn4FQF8rTMSRA
fVAr19Khd6iD2Ormb2yEb2IlrTso4NMfmBotbFWrRXIFe0IjMIQxlBrmYcpDfRl5e/bwiMOasebZ
vGg+sitzBraChB55/6rlXBFkwhcngiq0wXFzj0Xf5q5vwWpuh68O0VJoHduqS5jyj4FD4monm1YF
Kgd8VtC3MbVECkS+I4Fmq/+DOHjoxpjbJirWr1Th/1rZU7jTa+CfJAO/JCaICHVH4W13QgXojyKX
UorNI4wkv5kQZeSwf4c2vcu1F5E9cVCocmegg6EuHPRd8qxw4lPbwvGvhOlqTmftY7urtU3ABch8
5csL14+Ux3J1Ts0DPok2n09TeYd6EpI6M0ZtFRz6ikHIDJr859c1QvI8t/aL+GJ6GX3amp+ZYbEH
rKEG2UXK9tMngMdMPxKF/tDcUckXyq5MwgoH2IaPW8pGigsQ7SwWK8caMzhDQLsSSTKTbVyHyK35
MVYGjwKIFkyQOn/qWvuPR02Pvqif/yzUmQf9YRqS892mxbZMuFen1zx3AYi2WAN/GmXknAtnFyiS
YoPDcBdKy5DwScYRNpzW149ieM0IcrY1G2zti5/cE9uSLxzvQzy+G97Y24xER7wKMjB5XNxFuiYp
M320FXxjtxMZac/EXwWq1/DwWIwtE+l2OQ0zIvdx10rUOwMGMEDn51f7Yq1JD4oa3UEDmsIN3JUH
5z+9MEjUWyeh13r7G2Aatj27pBMJWXwDcPQqDcjsSfBxT+8gv/nSqAvelV/cOFFs6G64LqmvjpRk
8/5k0JglSEcFTC9Be1bqj2Y/5LjBQG0Z5aatrHSwpGTkc1rvYrC39to0FiXajj2/HnbbHUGLFx+6
ddwZ2EAOO+ElacGVYVcCX3hrST2h1XbgvPSjA3puNiqdgxUThtPir/2oxkdJv1sl6wsKXeblIqbn
HtiGhTU1slF214Nl5wp858fODiMR81+VZ2q6EpogJFgEZZDeRQ2TompjJxFlPJlSzC4w1yM+D5TO
qW7lpdcGtr5k8kCJAI65v40r437O7paj9e1dxjj6A4Yw67MqJaiBSx6uhEBh1XNi7Du1Gj9cx50I
yk3unzcwvcg6oS8Rm5wuDks1SnqDtl/SoBv9btLbtPuS5UUM4x9a/I7ZC1iETcrdiMx440Od7+Xr
XC5dviVHanu81yQVKTSnI0iOho/hwfSDNy+zEAf2N3MKbRt5sZie4VmL2pKsMQpaa2apH8yy24zO
Vvuklt4KmyfkdK+YPWrFq0qBH9nbTgu2w7LzsFJhjc4cXW7mQmAa/bmMitl9MdZBnnqQZiflkD3X
+W8FNZz4paG9mJ3f2SCtkfMT9w+mbFI4ooCU7ZPs6ETnjbrIVCwbqpJNQl4iFv6yx+iAn77Aeg24
bPfu5HWGj2h1/ImNcVcuLOpL+ay8DJ9piKXuatXJev7kJP6Rnqj+SMSV5/1WgGHWBGaLmXacj6qw
/YFJiOzuaYLcsvrTKg6Zi8kkNXwhETEholT+q6sJShY8alfXSTHX9LJXSdQUxlMH+ziABU2p5Duk
mY1Rd+eBQpEuANgMHvZKxrEVnSCmgSOROjhpQom3gow4xRrU5jOrvCa3+9CWTaQRnZ7FpR/wi+J4
YVQ77rCzCEKPysUxLx0gBKmzFbVvIRszDhhesyKnl3I99Kr+WN6SQbXJfYsxdDA3lXK/wZXxiw0S
FSGPTrZHajYHaaqSFEc/QsL/dZck1Fg6mh2vhWsjfKvo0BeS4KJ1OTyXIZHrM98a2owCWV5FFvsf
yXlvQ+DyiG+mxG0z0o5lsODVoD94r464iO6bPUp2tUNlCtv1qZnXUskjUoeD2G+rE4BQrm/tphnn
BsruRZZ/ptVkDeXgJADrpCUJjb5H/A0IadUZTmOLaqwxmkqbgZLjHRQswdBDLdPNHiy5Fj8a5Y34
O7C23FkwLywfhUIz7SdVYSumltF45iN0Kk6LIAwQLclU0JFbWTSesQNzXVJhbMIyp+yZr03uT+EA
Yd0nTZ/8G19C8lN0QGTe3xQ7x1jHcX6aJS/4z55rGh2oyBXDUuIUhjtW6ibQ6WWBjG5Sopn2F6KY
L1hPSix/lR75VPNHpQh/XKP1mJC++YorScQCX+IiYyJHqf1Dooq7+wFr/bG41v4wsYg5juYcOsOi
ox1gttoNIjsv5qZMLBqP2FCs6A6LsBYr42r0dyu0J8ofVC0/hseHIPyycTL+H7Cq6hixw/SpCKKF
YZANa6oN5LSEn5iYe0vz2oNM+Zfk5ct3/V7i8qh/BK/N07vmzedaQQY+y1ABcXdgtzw9y0Clx6fg
f1UCZH5/eUPNp2/Su6JRcT96ugJMuHBvJas2Z9EdVXh4Uoc7HC4LviA/FvkGvyW6fTnlkXX0jvuV
lvoECdRKcGC/kIsUeBMk17LnPlm0lDB/DwD0+lBO9ugVkwro4hrKORg+hJLZLUrpYq9445Frlm55
nf9tbcKCUgwo5p36NQ0bLUCNdyg62u5PRM9rpvlDcQclyIGPCM4bKnf+/IsYUgGAk31kRz9XSy7z
wV6evwnMicU3KSuqj8xDeI4KGS3XBkFLyJ37TEJjuzNsrvu7CO8xd5ZFeBYPl7cvsHzeAyemkv6W
NPTbw3sy+gWDo75ge7uwxfaJhcsJYBQ/VdwCihyxxQZYldLmIdidBVF1WNG3Sse8tibeu7zitvyK
SusXUVlldzRkwLqyUzwVstwht8WRQ/kujmw7BnCnZx6pT69suOX+3YuYHhEizAwf+ld/EO7dVpvn
BtGsxFuhIjof4QbVGqtdVqKU+gZl4/rRjSlj/MwIcrq0VJ2DHhdX3BafU6s19+DCkukGGORohbY2
zfmPV0TIKk26ZkSz0iT2Uj3N5TDxrWVE1AonUnhodMqmjh2eNBCKp8kLfx0IewdUFvmZiTycPVzK
q8Ek4yfanbZQ1WrLjjfKVzMLOUKpjBD/4PuogCF+R6IC9Zjb3duwfLXmPA8eUMhYWrgoUTBYKsPc
4mpSy5k5mLD2z98SWpRJJI2f+oUcbjNHLG029rY31iYYLThHe05iQPHn+15b5ewCak/72jseLRWr
eyVP+gGT1A+AThn5sXj+J3+GjJmjhTOAq+2JHjD/tOmYzCjYz67O7MrVPjwYGTK2MCAmn4rWtbiC
WPSRJ5QOXXU4PLgheomBoYLdq+CFkD8uQ3wt80HbSDtHjnBB5lohKrzQj/xCK9MpYfQl3IGiSYFF
f+0QsJBZocW9Hguq1S/xcmzwaYLRcFsiyo3yNP2E5l3KPcHyH4QUICqOzSdw1QOxJ6ICExNSYjgs
H39D8tVG6tK1VYmYZuKUVyFBDqIpL6F6vyDt/HN85/+Q16XSY2aEJsxYMkw/9zfMI4uBB+OH5mqx
hRlM4Xqm7TYL+49rayVum/i5XHBeM91oTAkfmsgpxQ9+5xWQ0cvK2bj720u6xYES5Hv5VbzLUUuS
2woE+Zx4v7XiPCPu/FI8gkd1AOuyJXbLA72Y2+sQGRIt5JXHwkar2cWVhN7lP/XPJh3Cd/mgi3Wy
rZRdOFvkTE9vXFWQxdtbDSszebGqOnQBUjDqCvKH29WFe+Q1ZoogCph8eltenQ+Y65vSKmuGPIyV
c3JgERfvyBY1CTk9YCCtivc4ts3nCaErE/cxYw6ZtZJaO51vOnwF9qwUB2zTED19WvgKrqT8ir3F
xuja9OB7gNObY+bUTSbDWyEGTMl8ZNlb1LMEWAIX2kFKc5Ljb6UN9TzoDol4ccCrbQxFRf4k1D7O
llGM/5OmqsFlkDXnNWGO39WoOHkWEpwW0R7XXbEToVXVCHchrL+VKel7sX+INcbsNABc/N3o4EZx
wssWi/jn4AgDcaSsBtNyxLxZYqg495kg9ZglTv1POgn7hzOE/ny/PCqtZ6ioYvdRGZt07jP19tmV
o3TUnPHKwgxhsJH1ssDdfyZb284Y1onk7ZQRAFlhyfaJukLIvjJv/gPreTQdq65dy3WovYKu0Bj5
wyfD4kkD1jdu0WcQx5vO/5RsaNuaBmWZnbRTOW0C5FAlRKM2TXQmelwHS8Oh0m1mQzP/ehViD7mZ
wtGKrKKChSacRyM+k8CwN75GJ/zqncIsqX3qKE9n7YtNsT4jCa0VleiHlXS9kHEIjKFkIeqF40kG
CCH4PeeCSi2e5vFabXXQHOL0PEGoYP9703krc6WL39p4+w3QLhpS0Mohwd6gUrEHPbo7SUBdynsl
cUjDoqlXCFOCZFFJzb70FRibGkb6EpX0SI+3IcvdwdPejDLQ7AiinBZwf5ArhSTuuNkjDBUocVEq
zO8NQaMF2/63yNuTUwIESQjCC+sG9DRewrRuSS5XLL7MCQClBilGLmwlZSMYWmevsAUJcKkwekZk
Iz0VZ0A6zppsIJ28WhrGmy9mGpMpcUt5nJp/PjaRh/HpKr6Lyvm5JHB955PzHdsGBLkId6PkRF5w
gre5fSN8PXWyjfTf6rVBEby/QzQ6ctEgGG/Vq2c0lxuk2zWuiirCBP6yWyoYvPGTfURn+e2zodG+
qUOboLlVdxG438j0h0TOaOZPENg4vwK2nvCYpK0Tvt5/4zrzoZoUM4wdS1XoXnq73G9Jy2Cj82c6
7t5qdsUsbpR2Ghhom2sZtgVSAamVuYo8POkc8upV7VAeDA1o8Ad11uMuB9diXNcAAcNk/eAv61h/
VxjpalO2C+BLjwcjfUq6881SMxARlGBd8A5osGwmOvngsjPgWoq80NtMEE+jBOvOMyA/k3l5tkbS
xWLfbnuT5QaX8Eu+SgsyY/HX+PCSG2acnutQ/CeLukHAKV0HFyGjK3B07X3f8SajiNqXfA/hZ+KB
ADMZHZAKt1ip93cIX0xMNw6Vto8beFkoj5ABQF5Py8RqK2OU+wetKEwGWvji7wUQOdQoo31vKTYF
q8Xj/O5RTnmuSseojg5MMaLyXS0li5DGvjkOETaSc+R20FWqWssCsc6LCoDadOa0WlfU8y/jQ7u/
oX33fRZsek86+3K6tSaOzpViGFzxDvzgXFmyLI4JmyVDHszPoYYfb25tHI7eriXyd+0q7LNyHHa7
qHA8+Aodo8jRkLy6aeEhnmWfoYgeiexI9zz7CQgY9QrUNO8qN+NVKFAUVyEam1cB1ATF6eX9oUXD
rLv+z/SM8/W1+M3m4qwDXs3DUcGUcFQhjTcPbLZEr9I8ZJfltsim2pjlqq4jSVop6Dg0vvceKpZ6
S4wNEup0GXZ4PfSDTwxTsi/U7BdnnBUeL2IeTJNgrODTnBIeMsJySy7pAStwgTe80Zlo/fMYXYn8
kQsH62yNxxvS5LHH8IScNHObZ1a/LglXCQlXTfWTpEdoOL9III+TnwJ3ju+RcalIlAh9w+K8Kx9Z
yyPoBNfwu166VD7MlWpVc3Ki8WHVFpKtm180ZVBbOjCyNONGZOnM/yTofvHxBN+ruHN9d3AissvQ
HWxVRA/0Kfd38LJv99JQzDBcw57m8Mc+iqKyBbUIk4G30+LEZPqiFidgakdXWaQtr6D+y7HtH/zw
2fHz/6i+sZq5JvofuWvMjuUpo6+BZZFXKEGLmsRAjZt/c0f1rfIRK2uqpFL1+K8cvqp9QodB7H3o
R4X+pI3Bd2ZhqkCftH/gmvRHCq/1tL0In0qAaStxyM7CgTP9HRAbtAlIGNbpIwG/Ok6TFhGyfT3V
WZAACPJKHyQf8DhIOY1Ucc6F+RaoByLTML3jeC9G6rEyMOCZFTpa89irjVVhIimIiFqTjYKCAQco
5Vk8uK8EVE4uLIrRgtJHqLCefBzr+6NKNHrpG7QGTdmp4Gt8nLPF9ROWEJSkHzByn09CypGmVEwP
ACr1a9t2uzjWt8mbmWuZAQQidcvka7uqNg02JMYvVTMhKr4PRlNjak7E7tgyGl4Fflf2NFdAfc05
8msa7tivnaHf0TpB5KgMgMsh75CfOnRYKk5b0ql67TdeDJw6wR7X/4EmZYdQbLktku7Vtbjh3icS
RycVhWXGnRQDbZ6bsm4WAJjOqiBmG0fempqb/qciXSRRNFeamPeU/fvzD8S7W61NfJ/UU52CmrS7
N0tMktUSchjIMGP40+YGgW/hziwhoOX2DiCv/rhI5F2V7/iGDEVSUlNNwCxfP5QqplU7st1DYW1f
3tDawI+ISQi9goMqio1O6SVELZDgt5i3SEZz1O91xVLxlPHYiXEPRVY8SsP5DMNBM3m6EG1k9SzV
0eoiONJE0pg//ovvk1jbBq3WGMgC2xWdUnR/GxgrbjojVrr/fWEkZ/2AB2d4oZLDmez7ryyaB2H8
XbBoFjAjb9OuaMv+7h2AIU7yGT2oSkY38F5sxPnwv9Wukw4p1H1PbqXiK5SVbGKlzLw6Q92rPBVq
lHsxIBOdyav/JX/il/l9ku18cIdXfLHcRnoRy3qlJi1XCzkPS5NuTBkTfl3P6eLvd0v+MAzvyLXA
LcZSelTXnvfAlq0LCr6zjJiOpruyfQVkRH3h4DWLW9szRCt6jv8f9fbxtMCIRi9eS4LA7s6whaTe
ZFSlbVGRlm/ByzPX6fKqkujCWbWA5pbgz60dlYiTuqxABPUP/+01Cof5LHg5QzxUqmC4w4Jf3agh
jr5tQAeB8ng5J4K4Ms153SeEd8hqdt0g4lNkaWl92OHMmzSFykeHMWQ4Xwa9Ma2sTyZWAg1X1nmA
iC8f5ZiDriHmrcnhaXQWOFLgL6gYcOssNQv8fXIt5fpqtRUkpzPT/w6HYKpNax3vp85Ci5tvYhHL
SWCZgdyMgt66CokIATaCjE9HWA1qcSDOeRuDe7GmpGUEZ5sMU0ewy34Yb90OAec0Ivpor4BGydAF
A04siokuQGLMu0+ypH2Fc9z4l7n792iCLvNMec9CYaUmFJfbmFNnn3vyedGC4/qm7edbceYCVJNM
p++lk5LVBxFZGmW1HOmY7DNZvEoXCeRIxewa0o2I43os8EkBfTuHt/J3rl/b1FrE61kYF7s2XLtq
YdMxs2BYi71jgh7VAc85++X2oQlKxQ0ftCrgn26S83zozm4ciG7hQuiYwhecC+W6LTftmALvliXQ
ZJhSD74U80n4RvAtTwd5Db1NDR7kdbA/84suEr3ZC0LHKFAJMc5ZESWMRCJEvR/dtasObLVrB9iM
XVqmr1laQCIWlfjBuxuSVAqyHxoXxMfq7F1MGz7oIHNjApP8zpRe5CrMGKeX/2YjtKFmWxUpqVKH
8gHwOlVQyvrKg6kqXQxES2PoLMesGX8XaURxcwTpEmCMeCuxpAL+rdFwKDKU6GG7DVwUqLZKysJf
KZuY94Z3iDTrASzY9sEo2DPUAbNqqe48TaXtBboFkY/FnmTWw8a3zIdPILtGQsb0Qc/7NobK9oo2
jj8wDhOpt3D5lIIYdQVnLwTFdiLLYjQmsJrtesktXGrJFNj9ZWFTYh/xJzG14N1bsnAUMJ/AN3C+
USEbz4NPWVovjw0LGEB4YnOuIeetTCPVZwEaY/LkYfC3ioZhTSnRMgM2PLCKFxZ2tYPIbReb7lc8
LVxmiX8LSx83UVv8G3W8rRhy+KMCqOwni7e2xHG2HR3W3COBNRvXYOylkXPxLrSIGBTEuC2hjAz2
4IpHkmJegDmSDpxJuYlvarpiT3zp8BQenBsaKhQtD9HCj2BngFf0hSlfZ3y+w+znV/6r6LsXgLvn
/rCbDICLj3SOiZ/QKfYY7NrXDozVeR3lZ0bj4HEVTQH9feEh9W5RE12Q1Bxmwfv/vk+sy+ArTqap
1a0uxHG3TtEUy1vHjMgvmB5UUi4WnV2dZfPVCPVVNQMoGFZ5r8ltLdAu6Z/Fwm6PB6DMfgSbuKAU
QgTDgG5nPMkNKMevKhQtj2c29oMWd82MCs1qtmkmLXs4bm5VbGwniYby7vGMWrReG6CG5xmlSkDX
/Jdb3fleBnDdN2c/caOzmFpKx1yM8KPLK9v6nrPU8Rj+tYOSzOmR0Q7BqI4i5u6M2EU1StFPmRoa
K61eanmyvQ6oTRJ+TofAPhdtaV2Z1Vi8uCJBNdMsiG2agqvQ0K6Z8kQ1vLHUo4PO2Lxr2n/wgjSa
sBSy0SED3bkDwz/l+IDycE0iIbGCK8E+ssI8nzk0JRW15agRs8HlXBjPfBawQwHrOnnuI5rPYsmq
St/iolp88P7OjDIM+h4Wn0z6Bgoew/lSIYWyVKUsTpY99kl9ePUxRmc8it9ByKN51MYmwaTT08cm
zFaB7D/sue0IP92FtGrhRfMo3SPUhA9Aji2raXMaRjnqyqzjLsmo3GEK+bs2kFEQrXYCO4J66c/V
OvL1RRuLYxNqKwolMvGJCkUmkcOAPaGv90ulmQMwE8jKco72I5xCWzUClp5PBFvgMYGUi9bm7ICU
JyQG40Ixt/v/bz3n5NkZ5DakrcTjrhvcUFPe/sP2t34rkK4PKLpIxqEWrlJFGPaWBUcCXKUFmx9p
glYg0bXdIfEd+J7suPX2ugQbUY9I3+qonNadBQO//ZlGQc6zRQ8ucdVjmBd0XxrxQABH+9EuVQ26
JoZHGxQhcvBi3qi3a9R5jldlMyQpddtfkyMAQ29lNTSFGs2APG/wkOxjTfi6vaCHK8oXrr4nClUN
7j5X7DpE0tdGxRoYVg/nk3c4aJN2o4j/goxpCXdwYMiI0UeTkTx90j+Qquwi9QSfVtuOuAHLSKRn
YWVFoi/u5w9P2qDtUZZ/eB411fSchwWUOt2oR7a4/I5mm8n76ZSmxHjoijxsLn6Gs4ZnIKjyGs7L
hcXEa6jmPqv6hzzeEfLgevyuG1/cYOtgsvqfmTaOfkFzKyFLDpWUYv1u9em+fCgRyKCtX2fS1atP
3mFgF706MjlvPAYEtZMqECmTYqDBa2Tw//reC1IYouf07XPPFA5tkNbsKNt/j4MQywod1+kmZl0m
BHVHAvlCwkxJACrXfB+wfPqkLUg8gCti2xfKUbALMtEV4m4lOAQeCHgcyPM3d0GQc61ULiH6qKxq
H0MnRO82JZ58k38aaTG8aGpe3DhX/BXTNdoam2ah5KDwKcB/nbzpMYkMywraET+Mhk6AydW1xbpw
iYRPbtBgxFZhNRmxIMuLbKGEstaHOqOGcmEo3ggNJgYzBMG8YC1CzMx0pwk9Twcoy9AOVqn4ub4E
MolMNw0OtbTbZYWVlAi0ZjJn4JkZOu7HTLnU3xj9J549geNZwuc573Yp9jDKQLB3+jlhOwsUlCQ9
EHqpi0rjuybu7+oJH8me7UnlPUO5dFgT2DZK2N33m+3hOFUY9fMBXGh5XYtNlX393JZBhSdVQk+V
ZTPolSE5SDKW0tP9zvsEJkAAmaRLFeAtIlyYuFwQRb5uaYLMw1LQRLl5URFQ5yIxfq93RL1bcLn8
SnaoI6wrEhNF9pdC9oLairsucXlx57sL3FxSy1E1b1Yu8dzVe+zeo0i4KVxeo89OUIVGDcSAlGwg
O1dCjh7OPXDmxX0yv/5UU8vmg9CbD50XPGTji6hzq1817Ej7QTXj4m6XzQtP2416H94WcpZ+oefv
WQUctKa7YY5t6mjVUJivsngLDFh8lRHz1M4srdUUbWpJK8W6sG+swHnrzGd2Bn40yQTrBuOEPvWv
xnPbNpQLz8KFZnRQ2HYUpCQONcflkwOKSmUpxciEOK+8n4xTlSoEPBr+MScvr/sjT06F/mrQB6XK
f0On5kBmOH92Rn/igvuXbCPbArdkb65uo9kzS5KkIklCE1PRGt0g785w0QoHtg60CYuo6hlKXecd
sZKrXBipWOWD0KqAVooFBK3plntYauINZD67L93ITgmzGTYI4BBFYDb5AZSLtmt4njaGvNEjBKzd
bZactIYphP8J+U1WN6XOkMY208NW/0WxWLXq4Cz4JRXalZC+Hu/P6majNXh2ZyAimyNcBAwaNoFy
rBfOytC+C+RXLPhFadMjwXWbtyZWF871WT1lZDGIUubSxZ5z7rpE/Fp6pkd/AC8+k253CIq0Iu6e
HBViOBys31QIPEoqAKxJKxCdMw/FOrWBEzkkTKXwEoy7hYnAPxStaYiQXdpAR2Y/+uPZ78JtxwVS
ByRFQn+jfYGAnvjUZ2+Ap5u1qSJ9KoNis3RLS76pas7qVR2YFGpHiezgeL85VII4+SziRum/Lmt6
aTTfOqmEPSdUftepJQvpxAypp5oGf5jpRTHeo+d0OC0Ew6ALUbGTdzwqXTTFxUqhM77/lLq9g3Ox
7A6/pSQZQMR18kGMjyTEH27Nu/lngTpoejT3GqCQd3pIlqZxw82iLGzq4tp487yuBCGu0fowBjLc
NL7Dz84/zsYReIyJUM0azdUNT4lD90Bv7kuZ6wMry+ZwXU0hI+dopnJwxHs+LttU8DykPbmOqyJn
OVqUQgSAfPwzhyS6rCiIhY1fcRuwiRLtBlBsbImcO76YwOcRJ981cakxisebQJrxI+XibC99JbY2
HTfHy73HC2xQodV1OtEASjSpz9TW3bEJ385ECVoMkbvfSL252+iTVkbEVlJotS7LdLZDbYK2i75N
mzL9OOawhUGCKk8lHM69tJMOsXSqmbXrfLy09pZ6XiWBEC8hKuWMTIqKtjm2Tf3jvgbPIedmoiSp
LvTECguDfgDzm33JvxI5YnR6Y9F7fMCKlSkiOxiNplsFhopmyCo0kNWtl5uP6Ns9O27z/VvbrV2a
lekzFjNU4JMO85g5DhL8Cnv7FxjIIQfjM6leOPz0Er9UGzJKE/paVNTm1/DamW1K+vmR8ZNHs6ri
PeFUMCUacVYmCJF5V87shCqGi2yId/G8M8Fo0wN82v8czqgX+qn3OdDqGUvu2K0jK+Xy/K5+5tyt
YqvWCGm2J8q3SvCqpXmxxyzATZDj2ShC5WDBSqzMVK7jktUIIS9FjzOKjqiJlzfdPEoh1NTjQLJv
fptxuutTBvNr8CyQjZ8rCjZWS17FVAWlA4/k+oVdGFc9V7bFQYhoY12T00+k/ECNglPVHvECG5o6
TOPW+UodpRapElCXSQ4pAovHR9wnZFcpbY3eHWBa/nZoasbo4yey6w9tjydBsbnSHpWmmfVToH+y
De948fe7urYyOx+JaUwfznJhAq/Nakg5WqodsyBzQinp7DbgPwO/RKYUJ76KmT9gIrN+ujDSdCCB
PT0Gw3crXXstHIGXR7OFihI/bODkKdmxNO31L85jqRf8K2/G2aLFptzqmCT6aSOvOxwBy9dIVXzI
jpVtQryJ9P68TYs4MbueqyE1toTRayWBhYrk23SiUEiHmA+OioP89IH5uWbcikInfl1HOsRtnzdy
UqaEFz3Cu0BgS6TtAtu+zQl+QMc4fZAmub776pQRxhcaqjZYOIuhCfFcZOVzRAlIeVjLU8gCCoav
wUQWUzFwDuhZr9btkm3/sEkUqFtlzHGt+5vofibv9f+AaCyt/ARuarItwq2y5htqTYau3hRL72HY
QerY8Oa9mzKMvHWXsNbteSe0Ez94G49CMvvRuuj/tY0855TXI4tFEuF3qD9CCG8WVE8DTvgVvkcQ
0Lqzr7s/UpSKjHZOZuMcYf3LOyroouxoUJuDDZzoUQGE/PkwH7jZq3SoowrmlwtB1jF0yXuhcFcS
bP09Se76a4ANMxZBdbFFHPLCY4O4ctpPtUkml75h5mHyGuKkre1xYraybzz/10a3gUtZHyIx4v3r
6hZ4mtsaGtIbVBcW1vrwz+g42lFJbCGacm12GwkaSOtGzAtPVWKBvbuLKfTj+/bDs+olGiRihj+2
4aXGQu7OQhOqmdCq9KUtc5hDYmZIf2RJp3HjN60NthFQNa5zuniPO4n7FyBzjOjPQbJ1f1mdCygn
nQL1QzNMbggyzanewl8G9btO/StQWxoUVwfOBYXmOEUJiRXaFZ+SxRsUIFzr+ZLnw3xzOk9uFQcV
1zyD57o5OHlSsMkxyYnf4K6SQbVcsSousIGYvsHaNR1AEIdg7IMeL4lu1H5FWsxdVgBRB1ptu7ia
4uaWI3dd5DVmPNjAZN9p/aOrjAE4q0HPASwfdR7t2Kz6OyjkoIeJAIG3rB6YXzdOIrUP1IVlsQAX
ZmfFovUdHxysZ656jvMRkttXkY6JKYvrpZqE2x2hIjc1FH/GCRy9wFfryPjOMhoxK1hOZiZqBVvP
HhtIrZWFQGIobz1xfDptofqSub2dw3v9K+5/XJWN+C1dvWxdgBe4gV3nzEJrFDQAICdjIv5OvHfv
Jj/ITR/CSbZsFhasUQK0f7V61M2kigZrTAbEmbWaEySY1psJbwCfiwyIJxiPwt4EET60X1dYA+x8
G4qV267nzsURXwl5s2CJtdwCRXZ2WcHmZ07Q6ttFX0JFmiCjn7YHrZSQeZcjcn4StF1vV1RAbW8i
l9WGT520ZGY8ubhp1tXUcnsehxi7eqtNbm0ATGsc4tkCEfyHvKX1X+EAJBEJiOtqx9az3dbombEH
DavbZQR9w4xTfkILjgS74WKtNdhMZ9AiYO6dN8FvcL6vf5orroqMfKlDR1SY7Q5e+Aza/xOT2ocH
k0kvlZ1Cj1f+INd6NhY7INsavYPqHlGJyXxhtC0ph1VOokm2OAdjwznQ0pCW4QUjsa8oECNCVyIy
h/csaGRkJy0/gPtEtknnGoAedEAKc5aGFoDyzXQ3jy53v51yYfoGEejXr3pDorROeDK+Zj3sHRtJ
mlgq9LlWazp+0MNJ/x1ZzTKFA4N7P5JibWthpCn+DKawOwz/pjcwdQs1Ri39bdRBdFgvxIJeQypy
wypc1b7Efz02FAPjnExP5L1ftLyqduLIsLf1ZEJcyW5L6QdfZ7MfDWgiSYfpBhiE/URNFAyqtslH
2AIALATUB1UBtk5otKex62yb8VGrE2K6E4RdWBC1yhVpbZD00WL6waoM0HU9+RCmV8qHhFjYtCgR
1iEqyaaRrwLvxx6NZYs/HPlYnTiNVl4wgNb4LQZulEL3I3mYRAkLcvQ5Y+Z5hxp/zpRHGS7ZJFpP
x6ijnRs0qPtfMHkYZEBEo6oNS+U5+LUaRv7ZB60GbCiKCIP5qaYBpuoFURfAH205mzah9gCYBPyT
NMlaj1+kM/9wHQvFE2BaKWbX5DbG65WRoTCOX+R9uWLE/MSHqzHBRrLH9eRdZNpmz8B+SxaRslPH
d4B5g4VoAk6lSXCe6QniSi8Bmmrc4isf+sVA+9IzJNFtUV0JNcmjvNH7D1wo/9kdm6IWey177LLp
MzPdlftD2uXy1Zm3ZTzVi2suzVwyO9ORFQ/U2qBdp+/Y21QgjoYaP8P4VaGaMXRSqdeb1DiHBHpL
ATvzK4T/3WF5+dV18UYCUv4rxgx1u6IzDCZP8T8TbMYCAXaOCsOaAhfPdyr+J5UUwETVUT86d8Rh
H9hWwVQ+SS+wkZ+ZgqOJ+ftcaRlmoNhCOZvYJJ+rowfx8xFpT3DL/fsjOSnZUDT1eI/y3bC4gVFM
J/y/AJc4lJ++hzT1H/cNgJBRHuN+h4/H0AnaV+S9twVVZCZwNyw8YhHEG2b+m4ZGm4nDdSK4C+2r
ltvIpchB6DEfETzxUCabE+sDfqoozQ+bgcPqq2I407gJOBnP8I2nh4HZ1wq37yC0tYwtNP/5yYDD
oNAX/vbvdBal6b+EJFVbUMz3s2zN7AaL6b68Edt+liaTKQ+LmpgqkIf5ifLL63XANF9c1BPbK5cQ
/BGfVlJQLATQe/bjPBMAVDu33UC8zARR3OeWVKiAtCSLy0XUS+Vr19HJ6BUeYr+xdzuCHlrgc/Z1
dtJD6+dEunahefe2dJg5Cz/JiywJDwRee7F1trVoe1YkFe/Ds7p3A5pCt5XpdyVXsVh9r/adAnHl
wW5/8KROyET1iit6xG9LSKPtXOSKZDbE2cL9pYhH6xO6hDh7lVU34GEoyI7yusFzrvxCDRzlvhEY
3iXum7UTrxaswESIaEyhKYYut2laRqJ7XkvPn0Pc5MwMPkt0dVV9V7XiFhhvUHTM8iMIz465qtwA
BUrha1qa0Zsoo9BqDtiimob8zJ7X7JdyVai/ZVEaOhtQrnYAsUOzd8QgiyhXe18BVa7nKv8tpthO
My7KOyGBQylO4lkmfHOe29RTpE/yYgjFEt3enYoy3C4lULhcA5oM7x1Mnoeutj0IzGgaoMwRLdUJ
a5jSRR7Gp0BHTOHmBcRimeMKl2qh/sdEwf+AJ9a3tZNcoWcaZQ7sahMa84xcEDsy8ueWNjaIXU2c
RHb15gw0ufWo6uqMhjCGkW4V2XHobNNo1E1FmTrlpLAVFFgOv4YTDIe8hpkUqq2rROJvcCJZfyGK
B6x1hCukfrsoQxfxMcMS5Edljo4f16unKNNMOZo5IMAFf76K4MpMpQ9e5RYuAFRrAOil34zFiI+N
LwlIyPowQLBlYGOFh4rl+4oNL+yG6mVHzk+WuzTAQx0fCJJMP86kCEUB39UWFFvLOdDtEXFDGMvo
WJBwuRxp6+RsPu4VWKOzOvmYQLxAnXVjEtInhPLc1EeSoCj7N61EEmHqF98v4A1mdjduRXErwdPC
wkFq4uit1oGUzQAsANvMO8fBpDIGT0AnsNVNkZexHTCfA8SatqNAodbvo9qXzicW+Y6frMBl/VmW
lZcpJRdHJEUBwehKlkmqm8Se1mHryNFiAFp3bjXUSx9OqzubKmweYpvbkpjoRL9cznvQBbY8zpVL
/vxuAxg32Wn0zcxST9zAzZQ7EtgJRqNZUcGA2yHloooN7xJrzXvxPI6yGvpC/HHiC2gr8FQnR1tS
QvfB7zTKIbOey9GNhqtPGEUPT3/3Z5GSmnXWQVXN5Q1Drau7dz5GJ53QI/Ee+nlhabac0vLAJOnJ
5aNljRmzHApDCxchwp9k/spVA62Q87FCg6lo6lYJn0sG6h0Mym0s68rMig8Mdr4rCfWa+F5fCO7Y
+gT1aKk/hMT63PSsdVW2NUogzcdGPakRa9if58IP4g4HdQD36v32vuToL+R/jvVN0fAJNapK272b
pZ3igJ8pxpqUVt1fUu5IvVlqeywTJieJFOwBRGwDlBGhypQa2OZKlm2UoRIcjwV5YStHT8PVx5MX
ErG+WhPHyEhHGtr9WmsMZCQi+9yV8SRSnpalvpeDRqau7w8IiFkqed1WCKox39AOXWTab5mU/sdD
O/Ksv3vkR2rTHtXaQHb8mViIQDvNR+hFFS4Jd5yBPDv2pa0SQMRYrvAlGh2rI8tHmmqhvbAfMl56
IJPcIksf6sUokiTQ9qFjGOmtQD6/5mskuzXNss0SPA6uZC4hD10R3dRJCv/+KQQeD7TRwMecil4q
OIbbxXYEqGA00Y8blfKsQBfobsQz1giWjxapW5ohlhICjOJemSpJS1psdcO5ZP5DiJyxSf0Ik3Ui
Mms4Zt9NFQG2IAibXF1dptkN7pxZTsVmizlsMwGX4wnYvSq+clv1Kpw/lh8+wljzWHSyEFw+Z8JE
h76lCsK9k9hLUWwZ4GL52zf/whfYDOFNjeqkW+1HoI+PgH7vbCdFNOxDUW1baZuXniYYV98lReLV
xTWXwj29CMNhyExL6ZNtjdW1qoUoTrpLJ/mQT2El9+HHsRbEQXwdbxoOIsfAoDpsFTWaVf2cZR8V
EX0+aIA5Mfe3iGRl7psZGeYjyATz2uLgqj0gnh9NbjFn+E5NJaa2QZW5vtvogzHl4yAfpd9OyB6x
BY/QxHjgWc7ckv+IpZ/2pdcIw84hleqvbnc0q4KnBZoeCjUv9pxi0TFDtEEPgp4Q37gMGb1q8hUz
sRyChriuzMRQQEFRTJI/2vmRDyWd1XWnQDHYlRJ26buZSsRPpZc18JisFkVa6EC666b5fTMVuMgU
CqKP9Qz+XdVTA0a3DrgBhy1Gp6GARvFq1fZWNQX0+TOiFftuTufq0Zn4uYcxmkv4OdfsvvgpLGPz
YXGtu2ttx5JP3oGF7qHfLvrke4KP4W+1W4gUk0RH1z1wibqVeclueyMAcAFli+cKYE9IBm78ZOGj
Mt2hKUqi4X7uFbd7UCDqryAi8YzbV8zYl01/40DeVX5OIcF+R0zlOQoiwY/dcPL8rid+HE20VnWm
2KiF1H/paJTaXbK9OSELbmKTdjqLWdon6vm1OG19aT2Fd9koSY7Hdgwjddg+JlrEMOVK/u5cYdde
Vwn6ueV06ZvWow3lzJ85IkRliD6dYamkdeAnoy3mwKRMkTNVVnGpLtwd91zTwEjb/sofFGVcJ00m
MSNQEL52CJgslXCojYbZyQ3Og3tqkFMJQAri/lmLaFVk1IleT6yazJjZu2I/O4uB7qt66ApuGcpY
/vYHUmn4T7djma5xPjGpOixhT6cCfu8KcFqGBBn0x/cddqALcOdC3w4Ue/F4xh4AIEX8QnoV7dNF
mxHiisrM8EdpQCLjv7m6y8z7VOZcKNbRPlT6ianY35T1bU6pmIKO4J996NqSbhi+JlxWuTxc39do
JMj9/evj9LE3yDZ77jT9OEgdcs2lX2+o2BQHiJFkG5hCj3bmxVbuZ5ffFki5x/LfQ5Iq/vOCvI31
p25jvXt9OxM+np2c3xsWF8/ac2vhRrwKvj4iAI+mLblgSkw/qbIsa7oIOrnNIqGyq+BqgPvKk4dI
Pc0r+IcfSoT4WuT1P603Gx/BpKflXMtAjA0AeHIcglUb5Wu2fp3cgEl2yFjx6zrdSAKmYte5akJY
JBeI4XOAIxOgavIExjNXaH33HKi3DN4sW5KCVpxWCNmoeRroafoNC4pclq0sVgjIqa6nMIIYirCO
/KLnhEjU0GFGwo6Vwo2k49l/50Blodd1y9smggIOoSb0iAdtRxTIU0sx0TU4rC+qWVNH6vgQbROq
Eag5J7QIQURszjwG/1gcVbr25tHndl+FDB9lafYQW336PS3ZhiQDI1AlxggastG/Lorp7yt+tPGs
yVPZSXAv/ipcPzENwSN9UdguTFjGIcI00vw19F448dpJKUoOonmdPOcRa3SOGt4PLyvmfs0T3qow
dJ8F5yfMMEn6pDfc4yByMhw2mIaJJxpLE0mk/V8ING3+cNGMKojrGODqhJwY3PRVB6WnjZjDh6io
MGACplgDYdI3qfsM1qpEkNE01sdzlup0dQ/8UgqL6Z+a2CcrKPfZVmkOZFvOoyHcQBxeukHdurZu
9OkUBTCRVlis2eh3WR+4l2ITqTmhf40+z3Mp0xM0AycZ3HqRprWni+iov1DhjwzDNAoXJqqAn1Dv
LcrqjsNRk+jGt5MtG8AWPVUdasGPmX497gUxdJ30yznAAg3/orah8O99Sy75i53XOY4L19skPNSd
aWoqWWX2ynPu4ogkJTKKtNeYarPzdaPyIFrTM6libXHYr6AwjZtb9bcS28y/ucKjKftKYRYLToF4
6AYIzfAixLKpiqzjTDfjlVqrwA8StJX0VM16PzdiXJXaeqz5qQbcj2FDptDOCdt+kbDOAHHGBcLQ
JwKF7bwKd3HhW/RGsACnfVQw/ZlJvg7hO99U7tKa6KKXbBhNWzgy0SX5lw8NW4jXg/fiKObSMQfE
C2LpZMAvwlZAfwCT770U8eQKE8jJxDvxjPoi6/uajRaAeWpq/dglrTexOxBR9mhXszTpzKvA/S5R
hWHJcAxbmy+ZjyFBNTug+xn1CzyOJSb31d9uRjkv+vro8l+oTRmhMTkJcRQIIFPNgw/V4ECNnJUv
kaB4l2zQU0chUkNYtus4xqeQdfi2/zJRexF9VI+taH7WM4oENZX4ZNVCmO5QXhQXTVrtbODB5VNb
axJynkj73ly2v4UKCo/O60yLdzqSLAo0TnrPL7hvwErGc/53gLrIAcYVQtD5GmP9/JC3U3H2AztD
OZcmuW5CrEUvGyHKwKYptABgcCfBeqU4pk9Kxr9IIDvW3HVEXXQGzGowJ1cFMCHMa63LBoNPMzML
ocddblqtdu6PoU728GnlOOaMx3v4H7enm6trG2ekD+ECCWwvN3jikB1GZIs7gmdTYQcM7NyU1rLJ
NyKuwg/DhupuO7Tj6T50OAtzOshDBgss4Tn0MzoCvfVVogq31j4VHw3kUWCh8xR4+cpRj+7poR5g
Z4UDuGBji+/fclPLVZNRwiJ9+gfXn8P4AYUwXX/FIoqKMAjsq3gaeH2qNsHO2ApAfk8QqTcFRFR8
WNHAJlf1PlccSnQx2D5tuWqqauVIvTD+nsZHq14eadw/MXXbysloFixnrCVfBcS+jIs1x4Ihe0tq
mgxCYYRTA0vaqSQpM6uQwno7vK2q2/oDqDPHGN9KnCFmSCzG+mxrQTINtahZEdIVzsoeAKQSXwwp
2Q23ddvAUlNP7C9Ninti+kUu5lN+/bHpCxgjZtlIxeyyQd0v5sVVYUVoKQS7u1loISKwCiUYvse6
pFTihmdK2O5yGNIpViKmF9DoWfBUR+AZHwW59CtTVCg7mWfX9nDk9sAtWZGsCzq9VNLtjXhKw6re
4OHTmk9hRmYKMsxVuUEks5jvgCK94KKgIDAnqYr/i2FzCIy/NBYBbSZ9lwAB94mcXTj0DyUPROKy
GfbKWzGngBWfBmNwnZLQ/ms+HNXN2LdCuGFZmvtvh9ZaPTLXl6nyMCZAyow2B1lS+A/Ug++MiLaE
UxGNKkm+SpkJwR4+l1ykR4hFhHniAx34SB02cLdnSMZrIxuEtMzSNvDsHpNUTrJoay0y5mjQ7/u8
A4Y68Qir2S8yvAh90t+hqEW5KcRN8XvsI6nA922ZgDEOc9o0CnBkN6T4z2yecyhPIdkZmiPiW+d5
9wc0RkEGI9Nnx/QdtVKp5joADp2qLMaUA7ADi2L3TlXMQ5c2VVnD/CtpTrWkFJrdlhd+JtA8jNcb
kzRibz868whFLXSvdJIFzzzLaWzS3PDFR6Xw5UkhYZbbD7FT27mFzvoWDZ6Im0Fns67g8jNB4WU+
ZboFsghsrlODi4IEHfdaU406Xw1T9DujG7EHcL4+PNo7tNxTBT4F/ZmVZPtXg60mWJ4LQ9CUrD1e
T8ETqLuOPZTU0OMyUFHsi0PwLuhn24KOitbXEOwf+fkww9N/pWEadoG14PBItYHh8HdLTU6XMwfN
FpHjP4yVjAN9pJQRvGpoNhWAwILw2LjRupKz95czyZa55R2cre2yiYCOcFDS0sO8nmoUx+mV+nnG
SoVrPmtNBBRGeads6/CHlk/t0zexobaDCdIjCDP178/PYPsr0O/j5KaPnsB69yh5kVKEbvUEtKXL
m745CQ7HiDiIYgKMaMSLGJovCpzbXTwoDHtrihBlR88FHOqbv9UmPeXqco/23mjFJFInU0x1cot6
poKrxIZV9Zido9fJrkv0QU0HfOYdXyoMlEcWefRtCPwjpxvEdpmVhU9CvPiN3ia3wVRdmdXO3qgn
Sfhy4eJQJb5MtqNxKrY5NeyGqXcUWTiFEs8N6yuEGZOvCu5evjNUgmGmj32j3unY8ES8RxpzXLDC
G5cUQWZmZkCqLQJ6VScV4jTt97BwE657PPKyL0KyD6gKbVA2DTSd5GV9/6PyJa6ME1bElbzQG2wH
RYbr37eboN2k+YiN03V70bQ4bAyJ3BDlsatw5uGyoFvujBD1h05qzEe3/5N7twdZrgS1ZJlBFesC
2iY/WCzOX09r5lfMPNYsf+qoiM5yn7ZWApBLRnsVdFzSRAb9QilMT2cl2AXf0zQveSGJA9rSzaXc
x4UMC9R9Y2nq+RNLg2XENxG3Holf0o6YsRefVSGWnErSXjJVA7m7fVW28F26Dr8BtMH0kU5DJfOK
mRNLlJ9XrlmUstNt9ar9/OIZvKrSgOMI8BmLoE4mF2a7SOfByw6uJ1IrpwS3ZI5JQC0gaRgY/x6B
2+OFLUmYPy7A6s0Da2euDaVRMZ4vtkhVvYm8zCHX3TyPU101qDWz7IB+o89tySQ1FV85IwYCuYev
VIt6uoNviAlRR3y8pMV1N7srOO6If5Zn7yqELGSAMnIM5B9k9gP7xl24wOw7LPc6AURYoJKUPPxU
TEopWNX+7J9KXZD3r6jse/D3Dwtl55mjgtPselbt8vSDx8HfJ/qZgLve+oJ4HKS3QGX/QLJE/haJ
aaxPSvDXfQ3VIRY7L5niT7qel14YybkZLNsl9qQJkWetNKXGLEY9sHUYZNupYUA0ZnM+xLcLHtz7
2JTaatQog3WzxuwqRGanjqLqd4uyGeq466/rmvbyH/xLq7vsTtX2Kh096lNNa5L0X11J7Tb2MGCc
SmhENMv1lJY68BORNBH3byBYYcN8Ho36CDYBVm+2zR3bwvconWwYQb6mIJzYSmRRuS4CaGOit6PC
BNhF1s21Tajzdaep0A81Xs5wbYDq9Jocu1GNBWJZnvuj2gX1KQoldrbnFNl/0KbiGZyfkc2QMj8S
VPwDJBGIEfUu5fujMKNyj5FS02tCrgkqTPs8NhPclMRpllRHCVm5YsrF6/kbtTRb/R4bQmVoTwsO
KUBWsE376KgmJ9cxSAq1KWxN1QX/YqvBoBkBc5lBlSebE2Em/jnyZopRxrIygghgexe9g1PHGqFZ
0/QmcIX8fU1d3ri/aiITBVdFib5qv8xqeX4lwpccUIkUTI+FBcmZjnPMALiKKNAg2GEYnYEr9IH0
6qcu/U7QKsBxCVojd8CnpzzmlLJfgO75RFjzPKNBSnRmffGWMed9AqhCM2S6u1voGDJZM8uxktpK
JOs96Z6tgUVMtUG4K9MUT+bGhL2+h9XLZJ6x5eOuYgRTq6aXVba+bM8hnjmdbmHlPIt+oW4YUBYj
xt+PrTpGE9yN3XuHMtLrgwf8ML9i+Od10a2c6D1o/CInWXmUYgquvpiCSkrxYg68SwoOZWJwPlR0
6G/orVrkHkND/4rW7V5/a1otcwg9uyBMuqDWPYizMFZ4QWqL65/FXdkR3D6oLFfTvlM81e9tVTOM
aJ5crj8A47wUiUrkSOziuS5LwuZGVgcORlguGRuE4IeTf+Y59vOsYg9OUcT381Gyvi2BBcgsKy5s
oOguBHgYjy4HBIrEaphhlfwJkiAojJHIywiINsLuLlGAe9GOroyEGF+FDUl7wmy6SvYOJzHmzyVe
auwbYR6ALctaRHoPYFvBRkEMH6AZo0ZACZhgXxWsBCwcPxlTTonheuc7w0Dei2n7qcNUPI43JoNo
Y9gokSIT0oHBRR9hGlkOaOKTHBqvmxf708XNW9oYdAWteA0OlNCOHdpx9Z/TUCUQBRm3OYF+5uyA
GdwqSnySIgXPCcEYcGFuMTce2IINqBhCdACYObRZPRKp2otBAlZGXgdsJbxKmjTDDxDI9br3d5//
NaLixoH6sGC2tJeKaoryUchwYyI+VqXq/Pr3kVpxQf0O/w5EScp9aml9og1b7PUQeljOjpT+CcL+
8jMmeWniPA0MgFMvwGm22hJlU2D5LYgAA4uPBYjf/EVnDnAZ/wTo8d7A5ng49ZxvRuplIcnLm0c8
+6q6isSWXxwodlxL5jSNFNJ3NibkKRlK3e4fk3mwZN0MXjKcmC3S/SE48BkyXoqbxiVOkpddCoNV
JOsy7sBJqXF8Kb7rJ56pQqlWV1XwRBZcblL6feLFMw4pllfJwKN996OdViEj0/xdXj3Sih6/Qi+s
2MYJVzLtmAvFnOYR1/3mHvXGWp1AIMDqBTkMavsQZTRjUos/GybYKbMQvPUjifLYVhVabP3BTCGu
aBeRHOqworuZub5TpFuwwNmDiyGZmcoBFO1Yp9gGhHCVCosFrdIv9FHX9A+gktZ31cJDfcTjTcrA
iCzQtOYD77FIslDTxmUNtjr5fxhdkwjwCm4uiu5iZZsizm8maPwC/P64tmYFvqqQw088M3VolYfl
xKHEP2/L1BdDd/TSIuo4Y/QcGzplC67xfRp9jcZ7xPqjaOhzkQS5zGep/XuIroRYnuza6arHomhV
R5lWEz5XHF2/1bneDAgrBGUmZrCrRIz7UaF48UriiPczW7gJrA9PIekNuWFNaEJGcRWRnmJ/v+A4
s2gKwilnflvs6Nx7rd+s4IllsLdzkjcl0d+X0YLND5GMtvme+k6pW/VivH+wgs0DY/TbVtP9MnAa
WiljZihocTqVdv/pmZ8jFpdeuhAfPtT3IXL42GQMJykSgZq+xO2ErvNey+F4jhRNJBKjkCaEs9/M
B1sbn2EFgLFMITR7+LX5YAdFr68BlhqYrY2tdNWGY2qW0MaN+bma249skTNhYkzBqOPl44+gyOjo
tXIsV42L+rp/09Gks7e+Pxfjhl1hby3ycDLox/aQl4t3eEBk8Duucvq1FTuvA3Q31/xMikRX6Hx/
EFn8lgAsXQRVJ0yZBx388vp3c7BK0eCEhQYkWqm2A9vFdzMVIRXWzBJ0YdjvC/JUIQgE74fAnlQG
h5Dz+ipflof9pDYIwe4mUkrXNArd4G2FSF4sAKGzynvSsIOX/1JCWAS38xZmHHEw2YkLIPb5XQtx
4VVhYnnr7eWMfyG14VSP9D3tuMz9aCh0HLYXU/bxgMA4KmNnRLYR2aVN9JfKe9WoPeF4+5+n8PMQ
FQJ5rB2uiSHSEvNc2XRAvGU1Z8QtdFIqmiRewGVUarOn0DdnIzcc9BJf7Q/qiCWl8ZJ3qPS+49Zo
6ANYSPSettVnpuofd2ZoGIQWbWTKfYJV5vupateuxnvR/79GCXQdVQkJW/CQWlZPqp9SuAEHGaqJ
U2z/PT2mGIqTQE0Egk3EGoz5kJgG53xo0iH7rwYN+f6+8QqyihHpkNYlCl1QGtDJIwrJV9ITrmma
NZ7Q5j7UXiuU+1LWr8GCZ5Z+YGg41GjCzDnLLgkqyIt3N4rXhD35SgHmEAIjJ/eAaM1dsF0tZ8ab
J09LUlFV97u5r/H8TRLe9LJZJv1uSHEBvAjlsiUrbu9eGuqN65SPx5bdTPb/SE2DYNFVZmP6LYD8
ieevDJeZ2i73O+hf+DJdy+HmXjKGWpk3lk/ECqv7gGT/xiNC7KCkiL/QVwIrNXsIeZ5kgIF7rNre
7908gijSt+ZYQsOdkUS6jI3al02ZbMideiVFdUCG6pByUhC7Mf+GQWHdF8ylVrb4WRH3UhdJ1tun
+/LDMgepDMpBv0HC4ydi0feaCfnHxv1hrPC7WaBVCdqbEBUIU/g1vlhJoNZapftoWQtMeW77Tsat
kW6DZc9Pet5fMXMU4MVJFX5nTglZ96EpSiYd6CL/egktIJNqUsZO4AN2QuJi1CvjTq0uu+7c2Rx4
Z9Kkv29cQ6XoJY9JFnCy6UJBgIvLuQyzPWj19HPcVF57PH+xSrH2dIWWERPp7bZ8PZ5g4qLQA3WH
zd5LtN5fz/DzEitStSnUB3tJW+CKNjOKvCMWHW5sC4wxdiTmNa/8SaZZrt++t6IQqSwJ5BNRZdcI
AAyJct6xWEGMU6nXpack3a/pxw10WybRz7ead7GG8/q7s5uQ2KHbd400lg/fsjakchtj9AcprKJs
2Q5t2hT+cSYAG3K+CVgf4MJrOGKmQ+WUwb+w9obDKoZaVbDyi8jfnO6cX8r+SEr3HdOOmDRkAmhA
534dcFPbWI0UXRICLm+LxBATnH2hHK/AlgE6opijI5fE0nx5rW0T4dx8R/N0Hz/aflGVnFkI7pU9
EPoGVXyd6yQc2pzqEvdFaov94KSGVE8aNvj7vbPsoxfmJj1zgv+a6YF5yR4OEjJSVr35T39928Mq
bDz4BrfXI4pbwYYQvxvVmXapTAtYb1Lzjvto553J4zKBbFNrdZSPVjIV117qtvrlZhlwTusSKu5s
CN8zx6u77zYbE2pokTeZEkoG4RqskQ0VxXFifZ728Q1H7Lof2KVcpkaCgUO7mubkQgE405lcHLY6
QttgpOYsv8WnJ1AuwG5QDAdgYp+YafC9RysoyR8qzyOJI0jaOigHsebtADdttl1W2nbTe5TfqOQv
oLune3FvSklQWd+J2bpjcAACxDSt4AJGA1bSeniur8NPqsePYo1bG88uDyZETcavldX+Ersn7J1z
OpeVh/M8nozQUX96xeSlFjghi9BdBV6ZJ09Txy+fRUXJZtsMMavOy0covlP607DZnSRyIlxM8dHI
8F/CyY2iAac1FZS3EYBRdYSIP19uoxi8YNaMMCV76bIyZ7lEZOZretRTVFA/TeBdoynXidzdvqwe
Ed3afkCBSavYqAFLqWKnGEm6YzL0BxGzfTzbzqy4pszp3srD2oT0N7emLM80fbs43ribgvJw/ClL
eupENAiRspEjkifjEbtYNwIFvsxr42e11gjUZ5WRHh1PLT7hACKluJELxY896oJMAZdPKz2JqCTO
KShMx/oY4qNXz340bd0aHLzhLjsD+FArC2LodlDV9dTrRRUjUB3RuOoOZ7dSH/Dk7Lxn/EO1mafu
olDseKnLgxL/rE8fCTGMjCRCnnKLJi39xFGfbRkn4NQnZZ0zOYO1PyzzTK+muFfQ4eUX9LN7u+Jy
Yi1E4VZwW0DPBwZNcUWb9eqqHeGvy/mKa66IftiQNElhfA9AwNM/Gf9p4QjaqdLu8ngrO3nvas3F
GlZ+M+/dVJqxXR33H9jtVrZ1T08Jw+NQNWoWfk416/eU0dSJdlBEJeMjGW1U9yrWKqKXs9614kNa
n+2+ue1kpuNiaGoJ3qY7KMjh3zUcPhAz9f472wwjbNwrk+l2jAv7+NzkKz8GZq8/98g+qtMZPEEb
PSxsQ7R1p6+ok260R6f/1QHz7a0CnmpD37UBYUWVnDHD2gBDvG+XDd+PB+wbn6TKQXlEvQKAIzto
t3yDrMSuQDUWfEDqEzOilwYwfB5Yw+RHzHW+B9z228MvurC7e2CKesfFMJ/zArySDk3Ku11WJENK
UqOgXbzCpngE6ZdXHZ8MEJgeKSv93p9VGetMQhsdd+ByqipIjvPTElhXcx5Klo7N0hWPaiX9jHp8
+TmKbyQZwi7YVHogumuhNrSGrKIkl3kaJ43A4PO72Shysy6nSShZdGjmDN5kPITPceb051UAJY/v
7EIhvnP6vN5+pBrYr+7o6GNeXPaoAe2aB56y7DaGMrndgCxE2J/C70zmoSQ0xDg8A5a8q1w6s5Fl
LUh32nEOPhit6ibYWEfH2PyWUKsvZji0Tq+f58sJ/KKg9cQ3pTxDhVw0Eb7Y9vIM/sa7Ver+MvnZ
gUZgHlH16M32aNFSXA2ZR9GDXvEuR+z67+yVLpumX498/y9r/WpQhp5rmliKlxfydWYNg893ewCL
taXYvmiXC4Ls0uwFdbT22ieGeHNOYRPrhB64HlLKnum2PyzOHMB5DaVkRrAM16Js3yfs2ZVK+/I7
CUpws/XmsEVv+hfyG4IWAGhR7ge+dCElMFf3j2GHePwovT02+5VOUB36kMJEdcSifqo3OnAFQs2L
YCAifO67uQzw45Li0ftYAWEvWaWXIcR0c1iGug04yZWzmOgdTldC5XZZJwQV+TzvTF9bgFOKoNcN
uc544zuxqfBwJtgA7FNA/TPR8ixVxPhB+hLgYyRqLQcW1TdOIIYFgXCQGGlrg4Q9HHuD14nJn6GA
oaomaMzw67Nsf0bW3YBqH8c0yzf7m6r+jKOMs27GrlXtD+dAjpi6AuTBAmqob/+F3ijm7n94w6oY
TkKM/8AohQpg517YwX2wQy8JYHSQp014I/Eol9uBdCDNfhTkEvyX5UzLRIeiOKyrK7ioZTKt+qp6
Y7OE/WOpMdRLXH51kqHv7q4ayBHPEiA2jLrMA3+5SiJmmLURBd029VuSI4l6HD4MnxXziCoP0uTx
ANboPOevj6cf9T0hL3ozIlEtAVtWJLujbxJajtiWMm4u1Ykb9i7eAj4m9LXJQDdynRkl1lXwXemn
fUEwyQal7O/D1J32+t8YD5UHAIy4PQ1rR5RJs/3bWE8xoqoH5Jniz+Drx7XhJyxozIptbUc6OHsY
IsaiqTBPF60NK4l/v4phsGFS1YGJ2GlsgqkJD8l4r/mCu6XLgqUKqhsw4ii/U81wr9XD9pXjin6u
bm1viNKHSeJm4H8MKTXB0oNSHHnC0EZ2HFsDDhVbVkdNs0kQxugkhQjVyFiMo9gTIKj9INWr/t04
r9dbnTZgYVerbp6+TVEZ172wQu2NhDKEY6BK08TCZYVXy5aqxi4WtIknn7cFOJjygNjsJoDX96GX
m2a1Kk6oEtkChOwsZ991dWF+QnXThFybSujUtnDpsmoHtP3hNTYHi0FF8cJ2kePu9p2sy8dbJgIf
r4dphCxe7O/OZEqlGc5WzXaHwLehsxPsEyWxYN7ad7oHIo2ghjNoQlM5PirV6BU5bbnpBIXxY/g/
Z8JdkcrgaQdyJIGQo0qFN7TbjHYyuU7kc7XWLua3VkN7xgyFSmjoLlL0kewRCDLPAbV3OTE01IVC
tMvN+gunzUUxzaxMHIzxMrNKGeyP+LnEl9ixArcSiG0ZTorPiW9S9LlGWIKI4NzLlmkhQ4LNtGrb
errK0fJrjtvI2F1MSB+ywD4kVyx8ruCn/ZsLDVqBXDQCEEIWCI/N3Ir0G+vpR89/lhdwrqyzK18/
NypQ8jNY6kw+Z0c9CSbzDH85fIWpb9rqKjtg9Zjdtn4NIgKqsDgzIjdkRCKHk1oXTEbFiegieXdz
dKkiicmWK8c+cCQTWSfJW/2+G9N9n0lAzrdTNRucm0zTa5hiB45Y8LUCdXWMzFWGHkJlitAozTy5
cPs8E6QNzblEeU/LfO/Cnj2+HmC5vSPgAvaosmHNCGS8K7gIjSCBvp4P6YVe2+qsJhSCa1GVDMB5
P//XR9YX5LFThOS4NNwVcHSJhownFDUsZ7pczSDj079WtYixqC45JC7ofW70aeZAQEC0wTgwWUvi
yg8GBvvDeqesXTSqOMyqKUniXS7/qQTrVbii6s9I/exjO/cBh8BIIk8jXxWFvxo+onWQwfjPZB5a
JDW57L9nXIzr5vZtbzTdo6kz93eTL5WgLoycadxMxf0zZtZUZIrSboG0ATxpbhG5vQ1R+K5k2bNK
pYMStw1uqIJUp72xtsDB389kN0l2kiC5Hcp6iXKpbuzCOWBa4u2qY1mav/ZgaAPybtuvyy24L2ds
wAGmqCWMjjWCFKb2zkZJeIquI+WjkYcAnBPwI1dI4b9WzD5lvtjv6IrT0kftylWVXU3r8eYA7me5
ixGPBvWIxe2wGNIJmzSZn+5rSLRMRErtPJwSrme0lrGqD1cn3+s35vI15frEo1dvpoTOz6eCqJvL
MuxBP9F1U67U9h+oI7udMo/VnrqUQEWevfEu5ykrd92CGZFcu692enpNi3gb8Gft+4Z71FfEUC86
VP35nipOJaJgpGpsZRJMp4wmqmRNPZLVSp7ew/ENGjrw7uNcdsHklrc2sTudUTAB+zAnyPhnrBnH
WZ2yTwECKYTyoP883GJLpx1wF7IO6jXUCZlqr8l51hPALx/ibM/wrkbwYelBuUFR0P5YRvsXQ29J
BM370+0hzpToZ1WulqE6Zdgi849wS4ZA11vjdDy9TMPM6+UdU8BYpwOkNo2K9AV9/uEUJb0Y59jG
BQ8zsErsjgGLnfTI5vu8PlPe9p+7+qCVk2vzp3zovDDNAwgbuRDVA++6LdFF4VHp3cRDBNNz6+hi
YoZbQPm6zt9g0tyao0TaSHqFycr6smZUoNQ23rMrfq/3lWhP9lxExbcquFcjnGKF24GDccfojrCW
toU5BK2ZrOwbC3XBiJMSA39EhGKwq4kyJwOtUdQfTXsT4AkjpL5BMaPvwCwKXiqJgdFXvyTYuQ3v
o5/oJ3dkQPMmN3B71Bv2Mk4zyiXBb37xgrXEHR5Sp4BSbZjV5auLq8WEVNJOZAG15fzzS4kZRKaE
9QSijlhbALqcdMAaDc+zf8ioHCi2Ia92abLa+nqu8cnI87ZjUy8XIBI/tHY3kPgg5sIfSV4ry6so
w5R+Z0nbsGCSnYS59hD6krj+yyWLF0lVpUKcAEo+KM5nzYoL5fhoYv8U97GlmimSYqWnBIJSZaIK
Jqb9i7jrJtWkiZ1RP5O/jBZn9ZvJzIlnF6xM5Cx7ypvjPyqmTBprpCj1p4P5yt39jZsyDBH02qDb
J4ix7SA4IxQmKQGJjiCWdYnH0C5NFAvUg3OEGblA/Ht/hy+hBSSK1gRg0qA/8pOrYCy5jUzJAofa
D2V//NjIjqT6EVbu6nLpfLdBC7ymACIR0RJignwoA/tdT6gYDqZYUrSRrCDofHWFcIUP2dL1L0Xp
TNqoDdCQSrENaLAIwqjnc820M0zUiZ4+EIFjrNbEDOaJ+pm6+7i9OVRyRBOTUyIjqh8keHn/90nR
avCoUZE3hBvIMcCHPwlKJDuAkgdrb7IEWdLqGs9+QXGnf0JmOIp7p6vHjWb5ghcx1J0XwK6Vm/BV
0W3x7JZkfsS3AoDOiFkzczKy9XNlPAms6W3ZahwgvPs8xssLPRm7RMKSl9InKeT+xUCUPdEAR3Ap
8AlISfTMkT1thvtsQxt1wV62SNb85sR408Kbwa6qimXPh+Izcd6CMgXbbM/lnbeGQKSNYcwO5qpC
AyKlT7DyAVdwyd7vMTC+RPpqyMHtBqSd37CBt4/ZtuC8xs7QLn0NOTbWVWISgBqWMRbpA0VTIWix
MEJQjfL8YAtJUqYEVGzH+QSPuuiPKB034eQgGDQ0kBldVRRThU/LEGb/OjBRrImP5xXTf37JfkG6
td9yDz163tEdiHLDp3y+tZ5lD6w5hq+yNEDQ4T2UHGi34SZ0cauj2Yg0nmU3wpAHXF0gX89mmYjN
P+eZSMxefdwyCIJzzlfPcvzBTOdEJItv8zhxTw4BKUuO8nhbCY680gWbLCWoz+LjqiL4uEy1DP6Y
GdvBYTOTfM5PXBlwpr1v6oAlrz00RBdGqQsg2F2pKUrz/Nzs+Zz8VR5443cdyqwhyvuSwzbiKZvE
xgk6cInuWp6RBTRu683WQ7j2oSCiksobdXpAQuh/8nDGu8a9VhRPS77+YbuJgoHY7VSn9B/bVJyR
WwGe1j7m0BLTkQtCZgWcLPp/RM4dzsfvp/9LVRHAxqXzPRG7otP21GjI8wjodQ8p750tsdrNudmu
GjOnF8/E2O6pu+TADrlR4gG+fEik33RtcwDkayncrKYNVcmoLfrAVd4Aovp9FGJdWUHJYjK1BFxC
nHAyHHZ6oxcQyjUYSQjsGLEbtQdZczC3p8VTVhkW1ISWWfgrXPsEBEyHHDC7Sm4GwPMI16irx7Zz
Wcf7S82s8/G6npGYnoNDfxqZ9UNsNRFlFxz5zh/AQsCxZ3EjqbRhFT+Yh9MHcR5kNuWhDa8ZpuDO
xgJmm2aGSRVYFGcZCjZp1WnUK2xkSJCUiAf9G9jVaFoenWabd6oquDiyfonoZ1TAXzlw/5N9rV3v
BS+c9SkZxZC+pMvixXVilkV6ZuLPauk37IJ/6eUQcFT4zmNjm2sjKRRxpMYScEogtizw5goGOCb6
Jc7hDw++ohGuUOVaKUlAEuWpALviUj6DpZBJbTvEW5jD21qym0L0jeN+PsVB3r3Cvx4hGj2uKp8B
AfNTzCiy6cjce/xwyLM/5QRoXgzRiYK6hFDUjjbjapoU1EdDfceq2h6S06uutsJWhbHaVRIQDsPq
a02c5t+8ZzfVmOS5KFRtwrBFKyg9/0DoqgZM+ziSsZl/VY0RLfnRIC6fl2kzbPRgiLwfYb//VgfG
+Hz6TIYVloD97rI83NbndJy32FwaXiM4vtqSqJSfpgsfCUNQ1zNS6mS9yxe7j52Qj/Jx70W6tZXY
meYm28pqGpBh/tkLJx+L+d99PzGnG4QsR4F2b45cj98ANnLWEXecbQr/oKBa9NqC049sdEnIMnIE
W18JnYSu5Bs42d5NZlMuOgySHtiRIuE3ziFqA399K3HwpefhfXWEe7iutk38zRYMXkvW31Rr4Irc
khFYDvjuNhGsZ+YAcqq/VBDQ8bhNl9waMjZgwIYkmnnr6gSNHoVCrvXLj0+zuXfYCMJ6QO+PV0NW
zJyzoZTy6ocxkzNFc0BmmJGPat5VLHQnN9GbP9kTGe9Jgwghi628VniCWvd3r7I37mnQrizvOoY6
XxlNKOiLuzDjymTK8j3Wl2hecOdrQAOt5Zg5p1oUFMeaJ2Ul11on1vYb0L5ZanB2Uo40jxeRyPWq
XgAKXNgUgomIPXF6hWWTbgefcZKyGzj2kIHAg+g7rJhv1kCU68o6Qu4GyT0xYk2poFKHBV8Cw1IP
pXdmLJ0p8TAw/FR5UGmLu9bQmg6kHzzT5aKlZU9MgxIHpFH9FOQvthnJyYszLcJ7W1VWeM3Ce6ln
p7UZxEmrlnc9zXo8/4sEcI9xdvoJJREGTh3EYhRjMnQtzd1bE/2voaRxDnIFcUGAiTPaA8evHIlS
9DBbFAY1N5gYHh7UTbMZREiNO/1oe0ADXCMdtftVd5xpPoUfXazvZbcXfsPmaMUOcsBXOr76KlZQ
00mKNzU4FACI/Ylnx4d/1XEykiFiGccaFWCTExV6tkR3U5bc79u20u16AU3sNDa+F3OXgcvslXKf
CfxepPA2YdK/7bCE89vAMzzpJmiDgeDUtU+rKQnRZaeF9lvzAxaN3glLrz1D/z4Lvy5hiSmT+BXB
Bu/Ncq8Y2EQZv2ds4kf1hIVoVhPt1lIYjctFgQNoImGy6rC3KzI8aYCIgEiuIu8NeksGpG5QRdgz
6PdKrqwrdMm3h3NAmgJ3kXDGLu1lg+BQTS5plVY9RYqvpOOUCRPbFyHK2CZX0GjM+i5/aeJdmUCU
oUXZHMD+vOktsjHZkf00vbYAQQsN5iGCqTcMZZh22v/pNPMg6w8/dbp5GXESkCrpHFPGi7Q/43ZK
q1CGGkubU2kLr1tyZHaEyvsm2Q0op5+hwF8BmnGZfXGXL4Q3tdDx3/UbyJjhYlQgeO+GFTJY6Og7
igzgYBSf/t+7BCUuKgnObHoEmh4IKOvmla1luEz/2FYmXP/pJ53Hni0j31/X6H9bZ1Vku5+d9A70
WqCkK91nAY4F5dgSuPWei54F9AWAUiHQAjYr8e7f96JN88zJWJgdvtFO4hl9hJ4M9qYO0mTbXf2Q
ZrED/A3ii670OoF5FupwnGlVc/cg6Hc9J+vhZcY26Vu+u9yElreIpB4/fEeJ8ycUd5NgT9mwxf68
OpFUGidPSu4RDUULIT/tsCUYvUH2Jwp2vR/A48HyVODTi7PhUP4gFBimNta1zWKxP+OeN9Oj6t9i
quHPefHdM9VaglwsFvpYFUoE7q2PhQep1pSpOgO/HuKCCQGOzw3vXsvc1CDlqi4df6oBCpBLczZF
XweLr912lua7NwgAfeCI8fISKPTKgF7XiXgil0JN+lF2BtgS95wnOCwCSwve28FtC+YKzdY6uS4u
9erEGwOBnmAySqlpyRNVWYtZXciOqEaqSDcV4CsGh0+zKNuSj8zpbXb+NjrFbfmC22qEnf3oZUxg
YUc3AOCBHZHFqJH251p4ECmtyGxopWtoAmlr3JSFy3NfBN4sEezmFpXTDjz79z2bsdeX6ie5pUuk
p3pfIpTn7P55h76iWXlDzULPDdhJcJ4QSYPpGPmVT3iXyx6O2EUp2AUyLmEZONYzUhhT9B6RK8v6
B+WnySp+Y//2QZXQ3tef/Mm+8z/duPcA0z4IvuEycXvgAOPHD7zXU2eMY4Y+2wRTe14N2yqBgkhT
upwfFuADPXNNu23/DZvSM4yL607nfXVKLYlah8jpcyArWbpniPknz7f7T0OJ7zYpIt040vILRkVb
xi+AZfC7WiCcMl8Smwmnll8fpIBtKUt9w/eCi7kgLaqFPZM7Phg+Rf/TVGV67xQ0kHEISsPE2tte
LP1+/LlZqLtn01iV9z+h/AqOq13prJdMdXErDNIrWzETbHT0eNAW3IvdVSn2ziyfI/HPvAHvdlQY
mdWFTzsZySvsyCxc95VNuSxakECfeosycN7jN/tblSHz7/8ppk78ekNQV58GHvkIs9qDHnaMYEnk
ouZIL5e9SA41zS/f+RI+Gjrp+mP41WwbEapw8I3Q0ls19MggMbg60HoW75uTlhwA4kc9VJFjnjB+
4gdAP7VdevoQ/cSvhcJ9evur7jjzErqARUVAVTHzrsnHwF81qjsMuQ47Ok3wqrHU7Geg/PA5mTPI
2Ei+Ig+shy8WkUZTBDnFGvnp2XpYC7ySuBqW39BridfnGhih2ntWaJWK+mc7RG/mtA7vM14FPFeD
pxySayMQsfUGimfCuoAAg4LjXZ6XNmJTHP54BZT8lOa1n+mioiY2vPl8EwPmUPPiKI9a4AvzbkhF
6viTE10p2XuE6muYVSsJEb6BP6vNnhh2c8aY+O8+3X0PIQn8WHRoSA8bhsG1yWvUS+3yb001PzMp
VcXFP29/KVsH2+vhyJ8eJku/QscInYajIaYSM/2mQZw4z0DLwfbwKMWuyTDaaK/iB2JrWYNVyev9
fCIMpNVyYIbXlnsgCfCt5YLQOe2rdxtH1ewL7YMvAGskapKu7XjU/jtpmE1Xx9UBuLdJyFGMqS7r
6+NcDyuBZ9FjUTDGcrSiqZcbbPgUV1P67VpQqngCFPkK5qDQNQ4tBaZ9kaA0d6i4aiLiYFph2DRZ
bLR1zuhuFD3d7/XSQoaPE0jZpzA9UZGkufQMFAvlW1HSuZD4ArEjWC72Uf5hzudNW9QCT7ywNicr
83wUJO4u3Fskx8dUyKIOY2W8SxgekVy/NDInFCx7CZkc1sbxFUTXDGR/22cW3OxErTlC9ySxDMwv
677y+PcFYYrOr8XHZdSL4Ka0ZFPUAF+syyeOKcJGAqolaTbMNww+ZDibnOPW+rXNaE1M3Pn8ByWf
tS0ElWSZJah7tmVCy/7d1YkfovKVVCpFAhyN1A4UBVf/lc22ACJ7uBA3Qj8tukYfvst5TtLxSBbH
t9Msxf7YyG69PfzrkDAaLYD8KSr86V22iuPKO7lcoXyDP1L2Gp61izVk8PWmjWw3nO7hVPicLyOf
5A5uEpDoU6bXq7TQkiMeANeb1qDVkTgK2zr7EI4N5JrMbKDbfMSrHlVywHKfjOSEaD/kkTC7vvdw
wNUa7z4wRafxmSA5oMASbzlkZhdvEdtG88Vb44omb65ipEdvs9jvLZYDUNw8mmrT/75gZImdh+aF
a4AQYb5WfKFGTzZecx5fQXawq3N3ogEOP18lbC9XOmMYjJOPmhL9+OBz3qlUj4uc/7nNRj2P6RVF
NjLIruzRZZMfIdNyrbxBcSRf/80ZPPQMVM/mh3pYhKyIFm2HS6iQHhCTEUr+xrjrJUP2Ok60GtS1
DxIYVrCjUKouMQQ4dipuS8DRbOPKT4hLed7rPDz0tT4kXThFPtkZaB58h0+XG18D+e2+FdiLAuY9
QRakTC65+y1J4a4oJA+/zBAwKF60Py195XYLSMrzceUxw2hrLgo7SRMySwS87xk4EPl58JQ2Rlzv
BQLEiYjWznQxHBkTgYGqIlFFYtYvIDY6+djraDbj2yi6pGcnywrO3S06i46Gqcwgi3VkNI6t4+z8
M2rrPL//CpdYeU5UVOIpU+YznSd7LfxEp7k5tV3TDyqf2f2bdXklqpGRg/3F6bguXUDdb828O8BE
fcYp6MCqQ1ty7RvML3PQogX/0ILq/dgFE3+JAJPF2OxusIrx9j8jnhTRK0lmAEo+wiyCqL92QMeY
9F50m8BvWnyt7hJJ273KTPuK/6CddJduhIGEjtx/rBd5JF8mVjotu1nrL07loJNwf0sKWZYD6vxv
ytBsejeU3KHMaM4o28Ho3n7EsckL6T4jgiAQtaJ/4QCGwaZnHNpBim9CFX5+1o8z593fOBNe4KFg
4XcM8i8AS4H6nuQWM8jw0J/riKLhvtrQwRtGhWcX5OCuuEld3E0Et5wMWrwm/BzWgehj64d2d7Xp
AEhyMc6svNjqL5nFvZLJRj3S2UytIgh+lUWLI90SJjjoH0Ze4aRFLogUighTCsNCjQcVpGcxN2Y6
LJnWtk92kU+nu8K2xVaP5NOB/duHiI+0sggF7QpIXIUxEccTj7t/xTTtvmpxABMy3yaBrnE8OKzX
VinuDy+R6JtlVKexnQ+TigXehmt3jJbu0CYM9T4ANH3CPTRmEvjO/mKpF08iCmLMTMd+0HDWCD8j
rUIHaYMnnAgYb2n2Ei0dqjvFjWWxBPIYJcfzV5p1PKR/rO1FHeZepwqibgxn7YI+eTMub+uTcTpQ
dUkL1BJGxAG1pPsW+ekHN81tzCecmgI1RGtw3yWvBwfZOndiRl6gZ8KOpuQTStHJFBKk2TKYqLu5
RmsuFYQ6eZyC9mcWWSRNjbBgGf5HfgNlGWNhIAe8BHUzxF/6SpnzdHraNJpwGBnDRU/M0LNrS2zW
dTv1voN69UxCCvz3YpkKGUGU/PbZ65Hcred+4nlrR9m//aB/hkuEGXnXJJ5247H/ID4jT8WvGBKD
nniVNXGSNbdNVyI0Q+ig5P0WHFaGerUgLUU+bZS29bwSSFm4ymdnQ+xNtjc/fLMGb16T4HiqOm7S
72Mv4j/DOYFq6hVkIVw1XfOdLrCRh5ih8BtGZzGURZ+SACzXUvXHdctWjm9+jmdpXYg8L5gX3+2o
xB46DpnuKWhjcOqddUeM/3HygnhCCQSpckKcMJj2if09NE6WpCnpTltdgGAMjkD9Iu8iREuq32Rf
YBUVOOWUmszNUxNhQ5OidjZlrO8JHFqCLYWEEDO44MeT26J8qKYiL6fVRsaY3gfb3IdYMSQAe3P2
fpl7Lp7C3FqMqsxamZK4EisEQIDOMj9w5rpBxlBAK+CFbwjbwzotYsVhI/dg46N0dl7ALMctMb8a
Q23VD7U8nd9ZCWYfzEI20ogiVuXAss7/R8KtJydqMLzrgr/UayMRtlcfZkrwzsYrpHaagYUJuVyQ
laUuRh88/FuJpWa7sFCGlm/VeIoEcIpkjW2wzkJ7zsdbR1gO6Rn+XOQaP+vR2I71jh31DO+lFmOT
qLZCv5rwHxr5b3nhlgoG/lLuEZvDxifCte/8zu0rNmLK/96zBekn4S6ordNZURyBZFblvde57Eeu
bWtCbjsWSi74clxAcnPLWTkTZyxQsQst6cA6zig+2RTJVFqv1BKb1dDn8K8iq//aKc1cH/f9Y3ps
mDDqz/rvN0YZuwlVpETBdAMgU9yk2Z0+S3rBMTHDdIbeXFaUhk57xjyyCymdUkKH3fR2twDCJMg7
lLUsoBopdJmVqg9526y/9tlF+/flL29462TFdYzGfu+76nh3doMXnPp8zm7RA0yYVdVxq9yAEPiZ
D9DnWqZlbZgIk0vbEg5PFjUbwwW6vdCHLC8aCQoizY47ZPiVzPQJQSGCtnPuVGixxIvIAABDRpBP
Gei1mjfkiPys98ZY3Z25CtjpP3FUIgMXk4jMJ4PI++kUQTqNhNhuYRvzfJ9HxLeVS1oN81KvkAvQ
8ByCSdnVyVQ8r5I2xzDHLGKMzOOdLlEHihttj6ynLlX4+ClYOcQWfHZsTrlKbh6JJP61m5SleznK
PBzeBInFRaZ0eNALwULwajjfbhkTlcqqqJGzNLQVhUcsg44IB4voktFP3B4RsTl9FoRmHkvCvFT6
wVPaP/6AtVVVw/6lir2PDwHF/WMw9ezLr2cMNId5cw9llnfK7lzt0KD9iV739DAPO6TZ6FJtRN5H
RqUyZqU3vz5I4udD7xAYfZkG236bWDovPaVOnNVVZfihq7q8GO/974AhwU35O0YvN0ClQ8B6Kex/
5zt3w7p1Wi3sExRgmsUwRsF2M5FmrrGpkiWhSIztyO5qA6MEgpvjOb+4YDD2YjR3rjT0dSlJUs4G
SU9U9Xg3Zz6Iq1G1rQR2R2nMeL+Tot0nS+jY/zcWOGqEnOo4XG4YXC3RPkhkgIejOkuL5Maxrt3P
2HA21rUSZR+pqz7xVHhS2WH7DK3JXo5p97jUdAcnzQduDNV5/5kzuq7Nh+AKqKZkDwMh69xjSrpz
mG2LylW/J/niIKBfRzIfG6A8hD6YzSkBgEFxZuLAi2YL76OFssVMaH1z07Smobuh2+bGa/hpL41l
yfP/DJsdqtYXdcFfxUxJz4HIkTkoOL/TtS397UknwscnxeGabpUakVWT5gj/7Wxj6klnnSNdvfsI
tzOpw5EIpTB/lIgNMZbdm02Eh2IJszRsCueaIsdDNDSvnpEI43iWQZy9PVPHQCLhs2me/BMozNgb
ZTtJbNI7fb3cfkOq6EYCxBxSyQjb3rW2MIj+sMv2NoKGWrdRpLVsGVZoLkjgFNij6IQxfpfUwzi6
e5N5sEiz8FiNW2tKCWmHLFZcOdqnr15hePHmk9EoTDroA9aIZMi51EzLgURE/SY23SlRQ3WfkbSC
Dh2C9wZitWlc516Mixo6aUXg+SjLTPTf6RwpmUkwQCZh7iPoV3oHjT5hDTOO42lU31TZ4f11fZts
B5t61kzby+zRMuTc4zvw6xyX4m1C99qeN5uQwbVP6OsPVgH5Im0+NwkpVLK9aB2eTmLvhl5EUs1G
P4lInohU0DLGAnl1xFjYb4HyLtrEt1Xq9MkSesQ2F+hDzVql8kpCQ8DFdHs5ZhXhpAQ9ytZZSLYZ
gL5SjvSsApV9LIHjmeobV4G9kLbJbgcegB0+VGv+4QH+eXChe2KucgAQvb/w1B6f0rJI+Rg6wzvP
CKhdCUNwwpufMNtPmFWc+GfeH9s8WxdzQzts+Osx/sqGXZ4dHRzqDRPqltJu+bRgtqnJXEh02TsK
A4M20lkfZjq4eJgd9fBNok7jfKXpNIP4Wh2To4g8aBkcxUqqRclxlkFN8EXmGK2EIM+lZoFZTn49
gUquPgbuUBdZO6En2S8B2NZyKn2F5BO3wnkWhcmAv23Ulg4kHtMNwDBA5H4L1xKhqydTQyHHvR8s
3Pm6g1p5aGzm10FhPTJiu50wR8R/63h1vJrpziAv+wIRCCbhOZvntKcCKEDpa1NVstNUG2Pp6FlR
p0EnSY/5KQX1tZBUg5rj15MhMc3I73iZKmLsV0oklgeNMQHLhUsBEldYMgExj8/Z6qFZ8aSeStMr
NfC1g4WYKQzrXxfvX9lNriM6zt5RT4vkbsgTBosYdrkH7uRGzNlIwmetCVIKFd8puTSg1AY+Y9F3
SQdERPZoX7pqeWc+ft3yPzxKh3OfMqacUBVJy09tgqdHxhjZ8nQ1kYex6mE7YjjM1gBTmDsEZ1pZ
WgTpI/4RBkZdui8iK8x9PyyxsEAOJAnKiNJJHVqamvDY5uuUyeaAVm+2q655KTE+IkGSKbVGL7yr
KoRUnmNHiK1+DElzI5LLm0VTvxsydbmRPXF0YOMgkL5UUkD/UWG5R+q4qD2YIf0x1ZX7aQingbzN
R6SOqtibvTDQHEU2lCzSmKugPsbXkAFzINRdXe3pIN6SDWMY68SOhKFHHt5bRgAHi0PVYWFygX+g
dijH9Eq4Wm70g8EgVP7YNzjVKKJns/9B8qrn4HTYH/X0r2kE1OKYRBD3/WNvP2xFxIdP2sjflxAQ
412Qu96kuVWGLcH8+2YbtJFcz5CEgp9HrtAQUo33TTv8tW0aN3A8siLa0aZMiXa5s0bZdjM20fKb
66urY8rC0Z2UOicMTBk15Tr9Ql9WO4DaxePw8sV280i8TC+Y5oWN6Z1OQ6BZr8lN25gogyIxAWcH
Qe8rF69sGkezcWOX4iS7hmycrXTHpwMYvuOLpYtUhRLzvTLuJKTL24OcAxTwwAW/f7HElaMDWraq
Umw+y9BEo1Hz3cerMgmMSwu4iGGZz9vQHzR86U2KBBbi5uQanGxzKady3WXOhXiFlsUSKUq0Lrjw
/O7P+Qmj+rBWg6bTRRzTCa+hNy9CFetIjECvfcoqOwAaQmDX5Py10iyGAElwEHO6OqVJgQjr1xrF
6o7O9jjphwqGkS992ap6iWPWr5V+TYB0Bq83E3As03aGUDHyy6osCEoZKJ25Ke6mtqhltMLDyRJF
nfuUkQ1fiTL1bsqDL3uy9QL6AAyHMlKUOu6ok/kpSOnW+LBIzzwxCUuCgKQ+f04Pk5dD3Y+XRI8G
+gj2hs0m+a9lUR34HrhDWQtojbtsmFWV3Cws0Dz0MFTgDqqBPyNgYoY7ZVwPJblDDrDvOUq7cv4B
AhI9KjyEA2irlJOy3hAqWNT8ug5J19SUYHyNmDiW1n3++YGMDmgiyigp3fWShsx5VtQkIl4rn2wa
M1cIlJ7Y1Mn1amRhenDYuBVJAOghkTNaR5csQCJnWavjFgaW2HoZRYTLfDrjXWNAEE2o206K70Ly
qO3SPO39MYY83WpiKqcRhQANTxIQUHAgTvDX4xu4TqqcT5I56omcCM7h7BLueO3vdW1xX4puZQMj
yHQqWk5jxzxFMhns9xwX4dg8vvOEc8X5XnGCgzgrWkZ8iiQogFwkbYHda8VoMtiKETsuCC+z6J1C
B2CUQWMEp9bxAT9V7tEQFCralhrFQHxbD7WDxrXAxkF0qv3RGPansWd0WIFCsP5a5FQvDuezchkS
cDCXlFNbBiejpg+fxCSdYAT3HfD4pMoz826ohU9W0QTOkFWeyC/oValFIYMwB01mXq3fxQ/oDtu9
+gWUXhw57eGYJblfrCafPDySBWw+q21shlLv4vpPt9+G1AtYpfvPw886zl4uNupgcTOc8/oEZf0B
1PEfA25K66Vd1yyoXE/ARPLbPSi1tQmzWsbkP56YNsGhOffePGbptXzDRwTeb2x88UjhoOTuC5pQ
Txrmhc5ek99Is76bA672KZLdt5YC5Y7CK20Hh3g7EGstNFpDJ5ruCvz37/MgnO11t+t0cotM/uzU
eAiI014Gz0HpjsL+Dt+6zAEj9d/pDTDFAfMPoY81J0Shui42B/A8vnCyHt+xd8fYxY5ebTbDIkWm
CyzyJQ12bkQMI2hhGpfFJOAjP3OAChO/LxnALb/Z6w/M87988hvuyGFQs7B6VyS6ItEUoBVLAY1S
K05nBJotNf47Vsq3H/fSdSVp4H55eWCV1OwMuZ1WeukXe6xNA+NBJEGyWlg6Zef81N3sieSyuMub
pzqP502EM7krXFoWxLWv+ixiV8k4Dr1++om6nutRFRtFyZjPmj5FBJaTLQc3SjGRQ20L6vy3jemU
mwyVcqoJAd3vptrzYC4TC4QEzfMfIoj+kaEnkkwA7O4fTnUL8srQA4FD6i9Qu/n4SJtTToQxjIAZ
pCs+9mqXz9ukVxY7ZH7M3Ambp2yaQ9gqJMVIg4rxzRnBCWjSbWqdGDUEdOYJ4PBFKh/GzAivRfd/
E2D7MCFilbL2Mq1/E3v7PVNSmzUA88WFQRZ0iqKRvU8lS+I9glRp2T7+UpDYo7d76jR30+7hnyz8
cbqnCH/vVzBjDYcv6DxYMPFj+rNHKNh6z7g2260mUto+UvKifK6BehrJxtFndgHqEWWWe+34Z5Lo
dGB2uCEH50ImXpnwjeE9a6TZv/KV8//55dFNwglz3MPb7fHVOolmoD6xmMi/1DJnm0dfrQYfG4eQ
u+qbfzHHGDMnLw1c4PBG7y/aGXc04kmpwvr72t3pwKNSCgzobXkAwbxBen4kmerO/xqi6RHvDg/K
F3Xg2oQ0dOF9mFuEJmfGDFd9ckmpGonTreJJCrNzZLZBrt6y70W/koxqUNqO3+P0OmaZ0LnjZO3d
9IqLrybjcABJZ/LbJNBjra3u8FzrsfPyOny/KMqHJkXUCoPy2aZi1fyabW5cloCYMW89EqR+7MYT
D1iJaDbChxHfsYW4sLuCeSZxD4AAcfitF+CX19pIId7iNNtc+IFroCGrr5QTF9M5LXRiqI9n6qLS
WMoD1/maAmwmPmu4trZYmylAWhrD9RJ2VtHn45u47glDsnCw9hwqlgfChnTiUnXaTaQsm/9Po3Hq
9iTetE7XdYy8ZQWSCGHS9nuT7r0ntmeNTIrSEsHfk2wqCzRJ7+lLHdWXaL1IiTAfD42K4O7zoNYp
JLp9Tb2K1wT5QteW92zRYZb5mhQA65Vbhnu5WtKCNNVcqv8w1FdRc7kCnLPexfFM5NmSbqrhUdpG
mB+zo498xNytA/H8aH7bOOvbZCOmFroP31VmjLt0Tj73ERQwgNp6Ekt+aNDS5DokXmnw8NxldCPn
c3rKH3w/pJ5H8OSxz9oc42jdu2aIm89eq+S0MiQtjm25tBydW6eL4dLllUCYKoa+dBnHXyBUfW3Y
mGzgXQIzeLo2vlgtv0ojlwcEfZAmwKS982gk/V4Wk3s742Q7AlJ0lYxLiA8fPql+hj+qgf3PBL3m
u19fJzEw+9iOCFB4NNsC7a/sMr25fEI8vAvkXI4ItTgYlH7/T4355yQUvFwcXT7tAz67hV8GpIpe
pYB0xu081qribOfV1pcU7lPxuCZpvbqdB0VTjSm7EZFFfA8eULx6U1K17VqkQfFP3iRF9+0RSxEN
pJ86aBPfSN2k7r7l6ROWAAVb/SzABAfICRj+iVBhy3UQ3bcx9y+tPxtow7xkcaGTZNTA7SQYuu5y
y+x03ugG1IisfPKFGAL708/wb/zfFBTUknkOGs6mc5TWLFXTrhNSxTde80DFqgYEmP7Fxrm2SP6C
l+3CEhNd1QBnrWxWFOk8uLGdBKWXfm0rUmLIr9l4oqFNnKVDgB1sKz0+ecw4s5rWd+3ORN6GAwGi
4FRvD3cK7XOgN6U876ibnfSaPuSfEdMG7hKj+hFwLr3eNjj5WkBCRraCtMWpu6fSzW7mzMLd2Ibh
PSqWaRBp1a67jnkEsce0NtohbNQSkOWjiL3Fzxbe3omDKGdZh9i7ExI7jaVvp3fLbIWiDJ0ui5Hf
Ck60FBJMDcau4yissjI0U56vFunAl5O91iD3vWGd3vIg8H0M0MWrfw3lPKorZ77qwkM7iis9ONZh
bTc1TFo70tA6Lc7eRToxZelWmmvO7mn68pzAobUu4AMDsk6w4L6HXtZehzNoPDTH5LKkV4jtJfCj
5KbT3iulMAc5ai9mH7tkENyaQyHZLnlvRUIqMT8KSRjoaPs+SBj677p2hhlpvjtlipyTECWkcM2M
XgOq7MIbcjUS1DhCVtTBMBNBqtIXevKpcCsacDfXpFQFM3tHCaGb5m+c6Are/V2LpUTqu2LYQWHd
7GJqCJONHCHkVY+IaH25vgz89j2qJ6cD2z/RY3sbA9Xvd+chPGIul6feOuslpIkC+9ZoqEc8j7zn
hfpR95Le5dAw4OGADcvmTfefHiYj2l4hfUkzmwDeom3w+Aoi2h5Zz2JuBbzWvBpg8OYdpeUvtDve
q4+m3poT5D8nMsoVgXAzlamHTXPT+SVVsTULEy3VrsP3OFAsDDZz80e1fX1rmvoGJCPcuUoM8JpD
G7Vkqgq7iDIlV3gn9Cj9jzpI+W1hr6haSAcVhvRz0bE9mSJ4pnXb1ia5+tyUc6Hl8/TjItHmaZFu
Y9uQ8516Z99zxkdwgxPuRlhFxUI3u1MrdrhE6upLukULEpYZ2E6oPxPlUU7d0/DXLnfsJiJ0N+gD
FYrRyS4KBi7vj9RBU+fJX7KrIYjfEP6T9aP9RY0gP790RkKclWFvHRUSwEQjJh0O6GSyGPF9N+zi
9TsjV3o/TQujj8OlFdp++Mu1Xq3onzvTeqFElPzsaZ+VH5qYzExJmBNu1r17Hwy9CdDs939vU8BP
FvWVGjVLjKcUAOw+eJdyirfNLfOiXsQ1WIeho9kG4tYFhpgJ88CuiB4BnkdEWfjgfRPyjTR8JnAl
Ni1rU5LZFLEqyd1nK5vDpFQSfNnRN1CaqdRyAEJMPWG4pVWYrTREuRDnZhqF/Ju3SefpARFRD/q0
GAXTLIgOuSft8p/V7yvbnO0HJIIyXetZ0VF2QoBaW33tRC6jhrAKga3iGzTwGDw7Rn4W3Ggadzxk
16NmsvU4Gi2O2PAI1iB5/79gTTDIhBdPveJjeGi4edvs3qedxalGC/MmZtiVZ6v/AC8LJP7wbI+F
PvRuDT06bKHYKEpMmHUvM9jAbjoLZ0GSJCP24leKRosFszmwipLz6B57HZjhRTnM2pMhSG+6BunC
XpuHwVw3RAU4Mm4YHQ4ER2OQ7cTuTj+wTHzXDwclXfHCVJEyLKeD6BekxAElL3t7vI/kGpxCN9vN
x6Glo58umyrz4cHq3kBwaLv+0c01IDkZPg42DjxEwFuFVgLvKnqX+ilLdS5Wf/MNbH1feu24RuTm
fEjW9K9bXHuwwFINeXxfyZOL+3ONcI1fcMnJ2O9fUSzfT8WqKu+kDP53yz42l9W/q/+Sc5MRyhog
mOUr2BgfyKR0w6VA0Wz0SSXhgRiBX7TtDRl/2xMFbjRME2Ob2z0i9PLYxcGoofRfgjUJEfAcHker
/iBj6UV1Apb2cDsYDSw02RKTdrH5Q115SvFPFLaRnzLLi2YPtvR+tP5pe2CFc9/gMPBEbxh9lUUn
cfK690C9ZU0mIWjb4fN6/3ROtjBQ7dMgVnNUlUp1BVNZ4ENYHsx+dLggFNFG7xxgEG+CyIWjAjt7
xV8GE8U9wTvDjk66ROefgJXlb8nTEdyONbwwC/Dk8BeNIegUqQrWu4cWV4ivn3jJ628i50Yi91lY
N+g29iWP2tqkxyG9IJL6q+M/gqk+Uvxc2PNk+49ISdjCYdkIaEXLxNVyck02yq9fR4kSE4rn8jmt
5uMCvs2yXFk6/ooIaWX9OrYsxjLcPGKgzmtnxvQlyQV6C8b0qiCMIBFI7SHREWtZjkBuoY+X5osf
6ZB+RVGhcxev/LpwkJcEm94AFZ4qhAvOgtYIMzc/S2dE3S9tf+mCAlWqQpwUkB9pW9fdWIFy7akK
CTbNuR79mmi8gItV6cUcNU97RzW7lnR5gQkQgBFfGtISPqC6UE//eHQBONk5gOhyhps+aYmIfArl
ypZ79nuwCFwMwhmlOIfX73mZIz5fbB7FF3BFPRuQTSJ12L9ygflaL7SAiWZqf42ILD+0G7gTQZKE
ogXPi7j1E08hJyv8/g18+g+ODwJIsT+7u7eIAgw3szXq1zojI9C/mj+b00Dgr0GN/6sSgM6uh+k8
M9hVlvemSXlZVzTRvSBiYA4XR3tb2IvH0IcXa7i6MYplJjFUExk3Zl4o7PaPSbYeleBVwRYLWG0z
9a6r9K83ktqbG/s4q4VWvxKw1Lc94WLnBcCIMM+8Kow/NLqPCAJjoJIwb46o33lm1+uQViMzlYEe
M3zoJMPELvJ8qGfmivQOAQptJWFeKHaeDDDJM/B0H3szsumK5q4DguyMZAGy+vCH8GTseYaAnQFD
D+7BbUZkCW5jjtqOZBo/zCFqXOf2MFXCicNOjz44ewJy8OUulGHgfOTMXdf9fi4hlRaZF3Q2jvZj
4nElc2elqYt5S2ux3TYtVt3tbvfYta3feqgQogBli66LcGY43tiln23aBDL/IDAhFXojGyzF96kA
ZKir3oRTbHVh+dkeVHBhGdpaBPS1ivpWs+ok51MLSc0T2rp9i12r9Tgy6ikLuKdE1rkApbBElQ5K
T3GyDI1BbvRnJIdv9GMHjYLA9x38AIVAgDC1sIZiMrqVFJHfeFvYD817wfTt/xMa3/PHeGJWmqGw
K+O7ZZHA2yQMtGfkpI1hJ3fJf6D6vs27Ka+icrUtm53IE06H/Fm7y7irC/imUaeqqUfqGOlbIGiZ
apUhOUnW8rj4udoNDIF9q+bTlsQtWf02cOfsMLy8x497xfKCV2u9a67LRQUvnMDyvFWRYwmFs8KW
OQiR+3MIBXc8zkhRS9b/77nMkc7PTfXlJDNwTESunPU6COIX674Udup8wIIaif4WzwzvuJ3WXjd2
Z7Tp7kqRfjwHhUfFeQox382GOvNHZa3kpby1jVjdVO8gYMwqgczBzjh8r3B+wo71thXvsvlYE30e
jujOTxoh42jhYXuUTzuMDdPeBBh5p5uCy+VPrW/Q5bcxS/RtpXK96R49oXVOgEdmM+GjB2r79rcv
vIUsnLxlKeOXatHwh7vUqMdLd3/3gZpCm6gxfGNNlFYNF7IouVJYBO1VBXsxAuLiklky3Ie0uNZh
EK2+ll9Q3F9sHibRHM9S44Toxd+/pDuSiG5pc9LyhMUtdXYxLoB+McsWLgH8xnWXuRBAQ0U28ka+
kluWDrDSj+Kf4tglIWrbHBfmWvb1Sb6YzB38lKGk+EfufeFPKMuZisWny+/Bg7G8a6p/NBAqw0MT
38SXHnvxECKs81Hh35LNY4ToOZ/oxV/XEDhyu4MTT+ev3BoOAVBBcDg9L4YPjf6UPqbh/UOqC7TB
sbsQug1FnliCwRRrK8J+b10n+NNgshEPD9X96FK5Bx2Y9QnzcO8kzO44yyD5KgLHNUrU+qzOTMDs
H0pvA06mnIDeKSK4Tmwh37uAcQhD2Mi435sNh44y1IXZeaqLP4w05qYKdGJogFTCGQaIj5YNOTwl
9NwpvR0mvnpiYByVZB/N4wWp3LQsJp/259tE/IChsQGf1xuWGita9SdI9/TCj4VnSTYTeQafWi7v
x/+i3B409WvCWILKCFb4h0+OXe4ACJHgJxF8L1iYcOD78u0vJG6VumB5mih57EgUKZaD1QVt+Q1a
ld6U+pNaDgM2BfVHWVCuQm8/t4PKy/8UjrK0gkbfcO+9/+mJu2/XGFsH+3wpDD3bIQYMCWFIgRwz
/NXKRtbkveLTaIsGU6LkXcJkLJd1Vt7gIPqLbAwgW3iNTCkJ5LwreVdMhwzxFdvCB747MpTG31Pe
mbM5f6GDmJwjpbqj1qygbX6AeWc0pmH0el/FWRUcqKAJJ//R8/R8+6cBjzg8v6lP1ru4GECvEtrR
IYU5Djl1mk5XjgcrBaNBuJs1qsExPgCJZ0RoGgDAB6iTkE+6OGSq9Y+hovHp0JXRagFeNftGo2PJ
Ld8v6iFn0+m504chdKE8eEdwQFwVUws6DnA8FnXB55eAHB/G4Cgtw5UnJYORhgJpIIgYC/baTyU0
vWVU8QdCEZHP4IDijO4QFI+qmhDBmcqV3vkk1XteCiZY2s5uNU2YHH2a0eZtiIt2CLwooBtP10ZT
Kixr4wmXx7OMRvXGYP/+lfnnHNqzO0aZYRKpnjpsO8knhdJ7KVRYzNf+9pD3AGtoKq99CpJAgbml
ZNJUfGm0XSBPlhXZnkOHEEIVXsTwelzSt21a9qlljtao528V07yp7eklcGesUe9+R4CkzHmIibxN
iqKrNAt1pViB9BnK3TaXXjN38NEyLXq5kL5t7l19FTW3K5iIHB8kRUWA3MbX80Gtfb5rhzAeKaYy
tWDWR80hBP7QwZcmUxBPueT4oxUkkEaqdIOJpR2WP3i9tsVvV2Ur7TfLYWdriCpUuy2Sup0l9HfA
+qDlPKKtWjiqQ8GwAchKbgrrizyRaFJFn9gyuoD9ncz2/IjdLjHea84cXr8h+R6+3qbPvhTBrWeO
rc/QC49XxtUImj6+A5rBE7jHtqmZb87bqTBm7enjTnzEv7nYfST3Uc9Vvhz9Y2hNt8wKjTOPv/17
bU+xXxUvvFjmhubDEwRYAvi8ap0tOzA0BlULznjVfok3CXGjzGp7g7ZVhv2x4bmE0V4B07VJxwMH
QZALx8htgo61kGVWrX/aBoX7gvJ7PWX3JHr3rZ0+/Ezx4ZOJc139msPIYVz3bSKyyCgV/tIZcgoc
+g+89AZw50AcVqZtY/vN0rwx3KKNYUSN8LvGssdngbJjZZRl5VnDxiWnoVfRK2bu8bZ+M77ObDOw
gI8hJe7Zv86FMi2o92KaZmbnPrDdHDe8w7lC01azYDOs9eVxGnxxtFocko4Q2MwBjQdPAPVT/ZzQ
mhADfmNG+VeYipISMtyeXSegmekmIbgEPdK58EUtcQYdv8E3BEYKaoJK96rJ0H+N/Ko32ID4itOb
zOC2ypeK0d/Mtt6vt1ovewoyRvm2zjUeHCYiWiF/EiSO8RA+wc5fGEIpeM62I6zemxeCidC7DaBp
SCjNikaJy1s0Riks1RgoSPPwz5PTAeYzbONlzkekV90W//n4mrY35bpoxGuaOGV2Eweaw3JNpD27
+UysGTedZyB9UIEJeLq6PnPfSpwvd5Ir460pZhyHJiXiDCScZLWlcE67Jo+uGaQtchOBvPS5I/d+
d0HTn5qgHziox1gyjoEmgzdL0qsCBcy8E7NRbs4+sY6BFZt2r8Nn1WY/8olwD62+RkUviUIGqgQF
8+XdayVnox3vD6YXT7Ge026/M3hktj7J+VsqnLa1ffzxorgXhKA4IbwmDbs8oruEi3TwSaTUHFgy
QCNqAn7KZbEgX0k6C20yfSe0Vbu+LblJD8x6TMBMKhSMlhrAq4KQA4IUbdAhLhVPewqCzi2f0MSH
/BbybZXE3HsIYyK2H13fqyrw5VxpM+p4PwzSMHPg8J1+2k2JaX9qkxUEwGdIIdRc7mGosr6CSWMl
lDawxGNP5NEWb9YiANmrp3jQrKEK8Z6PlUS9waub+GKtW3zuOV7MHJIORr7ltTlabr7t8OhwnYV0
d4SOe1jeRzBymcUHjodw5mjFJFOk3ALd+Xi+JfIdS1L95kYYvYPPFak5JVIUhY0ohYp9iz7TylEJ
oM89yMQaVXsBoQAiUA3EjCprJsFEbY/0s0halO/cWuVe++CoOt//WVU1fS9+s+KF1oFVt2i3KOU4
Qml/erMOsFd1nZ9dIsYjQHXaFZY3aRkifemPfMpsTGN12KVSrANsVnYdSWWk6q92sV1iqByctmLw
ZGwOo2sBMzWaNYoVnztKn8qHnUCKXcjk22oaNLy4ClXnI2BOn1N6lu6iFQapXcJCZ4LFdZSWjN65
4sZqze/omy5ewmjpom/NRefckHZAc1FDshb0KRX+gofdKsC/MNG2vLs9fAMzvfBn49+Ayqt9TMgg
QSU5nJIpXKdyeAg5rBbnwNmmfU2OoCzncQ2Ad6z8brYNqna1LY47VzZm+tWtrUOsYd0++8fGKlRD
R+IMf1repLr1xYcDa7tOBBFnpftp1XP6kpy3uGT1BINVKlCFtUoubP9y7ceGe8733fYBIA3xm/Ie
85NZpT7QMzF6F3+FPU4hqjW46luQUnBIcO+GnaaWy70g73GJ9ZvEd3Q8qIyH9X5FGTtH1QnCQfRe
DBh4W2gqYGe4DGxV59Hk92QcdI7hnlcTGd1BC7faVfAJUtm3A7wVIW6/pEfyFdxhWQvwW1o2zp38
RxE2QTYeBotBURTFy2b21dy0gMQF9KWQ8z30gPGWoJ1UDg6jOE6GopfrDfvKGb1cNciLIt5y3aNu
uZ0QPJ/3t0CHSUG2w766Wq/Ty7vcQM20ExGrGZN0/sVJzyeUYlOlImxAcd+dP2Yyv8/TVMUzLNLL
RPeCP234wb1SqGRb2hQ3DbTfr1s3hrOX3TdcVxgkfhQqqlbK+30pKmOeMAOHdvSS4NY0mtybOGjm
I6jYKUbWvAAibYZjUMoeq0FQ+NI71I/djnGopM4Vv7Nt9b8PT51iAOBPV2yORQHBnfvIW5xF/g84
c1GwhYyOcm0DbV+/SX1M7YlmqUb30N+cQyU0DdYFL6jv/L7KDfgBzqheG/zkvQ+YYEcPf/IyuJGB
MlSx/Bjjx8NI2G0vapkkjJzN0xSuWdBgB2yoYuAA7QgOGDoBnS106om1kch1UjiJrbCrLqD0gpbR
MJIVzg6vc5EWZGyl9xrjg279kz8tcD9N+m+ThjOLvj3JHM4Jj5Nc5PQlrIL8I7hDteBcitQjen8Y
hqrO8Z6DBSoIgxfywza2bf5FazAiMLN2KodBwTA+uFQbP4EdzBXE8P6j/wfk8f73+P40oXAic3IF
u8Z3k8Fyl3t/OnLiqASYs6mC06syPQCrmd/X6eHuLNKotgJt7xfsSEdtsnh07sUI57JFz3Wb1hhY
Sa1pyH3ASOrXPOmFYQJwDtUCIz5ursNvGPsnZezFtEvUWurPB9KaB0+9dSM2C92v+fCWFpCJTZbA
wsEXA1wz4DFfNw7+w+CXeIeHm7TGJh+XK4+GexcP6x6NLEpLVqSemYygXJGcaaNgdxrJ0ySK7Okn
5w8GM5r2al1pMq2rMApB7G2KpsKAvbBWjHzINYLwsS8PATx+SqkVpda203COf36wqKMEHUDy9YUA
LR51SZfu6zGLfCVCPKh2pk1I+UslcuYstze4xPODau4ib1do3u8QPlHvPn7GnbwjpGdqjxYGarU0
U9WKURwsLRn5k950YaTptUIrxRmkeYJVY8xMlhZ67b9z+E5A2jk+lZyLC0NiQ97BE8+1Avz9N+wV
ctIkdU/mX/6thf3lIFD0iKugl4ZY8QYqVzuA6lbrxQDZeZrWLCObbcNCc7uo2oioJMn1h3VPvnFy
btMPmrTTn2QL/8M/kaA7eJMV4N7BR5N0Dw4ujCmFdCTGZ+OKKmCz004xt7vyemN0QY1IJ2YLoziS
Pyg6uWoeVqDM9aBUGdAuXjd/APHNHVT7WB5E4gEn/czgDsfXnx+fzXh/WBSLvcbHvoqBlCWBkzvy
QCOcmYbyoc+RQPlIsNmfcPKAocRU5oSFOkjnDDK0GW8zZYjjjPckJlKML4U3bH3eLCAg2Tjn2L4o
asQe29HhRQmaYw3/2K4SqGxdcwC2GtDjFrihOSZRqvxnUaevJ49mYM4Gr0ui9e/iHNpDi4aP70g8
pJ6ccby/AAyIHhxUsOoMaibtOr/I7jzmJ8xTlBc7pWUmkM+wwwRH8JsTeEraCToTdLFWGMuwHy6z
wSBUYqdihHbCiQ2tb75gMNDuwCJA7ZaHkHPODrqvgVMy+VGctMm66hw+JnLE5FHsezRFl41PVh/G
nGcDFSIZuYh1kdhWr/MaurV/U07s/pYlp+l1565PabrBsZ9yE/gJFG4G/hNgwLItI+5EFyloVoxT
8tVZmv3sELMo8B2G0J/Vox3xtkvuCCsHKcO3fiFTksIaL4Bh2rFfI3jM0+60GScMlX3xEC+o6L1C
A54exLZN94jBqITQ9d3Ja7PsYvYbQ+w6AC7wFG7eD9P0igzQk27gGUn4rhfA9+zeEM94PgTy85uA
sfYAItYBHh8r5Ur9I2s45uztnasfYtyCwqb0OVIoYFvMgFS2kvzk4DJJFF3vVMKa6Y+hRbyH6jOl
/2VFy7WZ9VrgXF2gdx5QfCx11wE7gJ4Kmq3P+z5yxdow2cX55fTiDIe1iSlw4HZl5hi4ND3wJBka
Y5U5IgdLqFmMg1//4oUNG9LaPPzxLUCB/q9sVZ/wlecGphedGuTQ1X61VZqj7Ajv9ukXVt2bc/1Q
LthzOG2ObBsOrAKGb3XhidSiIcMjx5KI2GU9E+uGGtsPE3tX2xMlCTYjvI+mqOzOGTrDrQ5mpkde
i1hQBrXiu1TTq2996zM6ih5k6961fqJfRsNUp58X/kiCMtv0qnH/wPOhlD4WNO8QerNJgXBGdPfr
PI804oX+lVq52wuoJRFm/8nEp8VbCCVkVpi0qpy7YNTbzXjpOrm82aol7bHIPht812cz7a3u7rFr
whV7NQOuW59wymS7qAJ6Mmv2mcFFu5gTaoRgl1w8RgZTyKoKIpySAJ3F/c3xpCHnLJ4l0cO7v80f
cWa0Iglm+D6W6cwqJvkiobSpDVQ6uRfEc1HDPPmediV0PNdgVFUEe0LKzC58aT7EgfLq+v/KxlLq
YoC4eB44wuWVje1SMkjxSUKCaVssA+Zg+QtbzW0k51DL4MCTFQlu6XXRtwoXTsg5mv6TMVfnlgNF
pOBC/TMz5YgYSlFpcMkFrf/LWPQ+9MazN6lTkiKlgYZvnwbFv/L7AR7nPuy3uKxb91leaoGwI4bR
RDNBBarXttPiTwod/9PspIlHj8rep2WchgaSE9LuWJQ2tzCYBXxBBHoCRmpBM9kqkX/5RO0DnhQK
0LD3GjV2TJn3Wa6+J8TuMpztqOXUgob2SFL1oTZSwfzTGwCe0ZsodqNJkqYoTloZS8yM31QPw55z
x4P6Ns72oLjgMeaWxTBYxTFowe7swzYwIEfo2PM9O5RlpFk7iwMi7KM6Ilut3QGE0RFJdtKYZn92
GHpMPOLxFD3PPYwNfCV02zJslRXN9Gvb/F8jh+mEbjNzu55i7iiUw/btejgef81jTX39P8u8DAhn
nOhhTgz5fPy7139c1A+ZElmuIETTrdcVxNMtghsie2kzztZdNsr17c6rUIIOFpoSk5ReTfuBOq/u
/k+57/Kk5AH5lZRypgGrTTfdskcRfID+nD16aCy1fAYNXO43JoB9Nuwyd/MglrFiv60viA4/4VTt
zX0GVazpbcpRvMRovSGx7ArWoAlx5tHeiUd0lMKviStx/ATcrNt5rBw0aQUhk/yE6ZE7x2tblXkc
5a+8RUjP3jTSyR/9294trNdWyaG3QFx7uA/bTq91w3byfWIRtIXVKn1znKP7+whNC8DtjmIFr/zo
jd/v1kFBbPIADd6OTPs6+K6xy6dnFeRL5ORRzSy727ueklKh3NkkAkNn/6yc+l8xfqATiFn7mPV5
tEFexWcxzCfB+L7+jvjH8lpdt6+1Uw+F1ouuudInYAKmSwepNDcHgLk7Kr6VdqVoqcbtIj3tqIAe
CQTmSWJaQQPoQYpjmjWUxlVCv8WYJMFBPi3/4oLurunqT1npxe35nMoOgTHSbwPVPZE8NuH8ZeVq
QvHORcw9xiCyYHIqhoLoGpwsU/EnXCOvoZQi+SgYyZlohbdh9p8SjxuiA7U8AYBRO79kRNlvpJor
euYYMtYS+eCYPkoaF2SyNaiBPPE9z5bFoyHcuzjh4ysB0cpPCC4XAZsO5CwcG7jQjX/EpgYl+Dfw
+oiTx+9l96IyFbvMy/eMadqRToOTyUZUPuGEfHKw8YT6HEKZa+zsJi/be/fR1RiUSh64ChjAY0NE
M/Js2vMwi9jXLTpxGRWH6vm1Mn4D6O8407TkI2Jgwfm1wjhdKHI5cwvgGlH7VVFTspkOuBC7x+tp
VnfP3b1KKdJkt/x1RW5LOMoYIZM9CSKNe2VTtGa4He0znSbm9ne8tmsStBmJGwrhsVH2SdP13YAU
V++kUSkmu82Xc69RlZK9BsgWVn0KgWK9Bzr/fzYsZeYAKAwchQpYh3qdEopczT1r60guiPmSMXlS
p2PnT5HnhWAXBX1JkfzdBJ7I6MmXDADIIXm4HOPLMHVI2GHYmueN8GHU5yvGBEOllSmIVs6c7+Qp
srX5PjH2fpLJJDUC7nkrX7pESc5h4BvBtVNIN9aKc9OAg/RlKq7g8qpOmslCLt2c+qr/wWWRST80
0FHoAtct+HSbE2FVM8/vSOj9nn6Tt2Bp9rUotJin8UsivId33+qW0frw68BXhD1XDAQMBRL0fvvr
qEt10EhZyfDYtmyHjuY7/+7MTtJ7H5YqRz/FivWWhOQ4OJWJEsgDZOyEojBlmSBDYwgqHTPe3uG+
DNoeK0DeHDQdFmfPL9p6Ybvhc1PU/Jmc63Ufrbg2eM4YOYbov+STfQi7rY87TiQNldjR2uXGmdK5
Gz8T2z4W4AfcdSON6IWyT+GJSisVyEIJkXdTfVjbq9/i12Vy8LYf0iilHUt5jAbaRTnxtWFne0CT
nvxWH87ruasw7bvv8tG/zJ+2zYKvrrGDPE8qrKAuEeF/z9XwJt9lKyFL/Nm1A/6q+hM5tDaho4uu
pJ0e8Hh3BEVwRV7CNCo61psjswQFQT8LqGHey64tjKiMgj42dqiynKTE5VAskfzc+Md7/1ancfqo
d+AP1OAeYrkCiJ+OXv4gBxwpBvMdaYhwpcAdRtJGCspL21WmkqA6lq0ePAiKMjxcuqvhpL6kNikX
t/dLfcFz4XvpiwBE5PYaehpeWf0nE+bxuauytj0Qvv17tbaSWXO0RzGraC1/tPmyekuRqJfDY2Fu
FwfCvzCEhZf5iDr+YY3kjPCe0tk2ktCIORjjYrX63uZBn4UVxk7OmMamYuQAhqEvfv5BtRVx9gLC
FzoeimaY8DqunO8gFCU4CFeIowlbQWkfwm2AlCfiCUnlXNaklk+wimuGdwJw2xGNESidJvtW47Jh
OpjceucT/VWBfocnLra8rVq28us3JNNLXuV7Z2BQttH/GoXdfSrQ9BXXRpqPJ751W/5e8FpxmaPT
bSHBGZx4iPlwxmbWseu5Mhg0VVRRXyYV4M2zF38o9R4Bx4Y4SH5VE34N8Lqxk+4BZBWH7Vwq3k/R
SSp3C3/WXTdOG+gQmdfaSxCAxuAIB+CskOGlRsPz/QJ6Of8iz79BEJc3mtrkzYiYc/X7gQwGcdQJ
79NtoO9eVPGrs6N/y6m3PPxL25mF0WHT4Y4F5dRaEwFhYUPrdYXvI3SPpANc2bt4910EFM56Gz6t
ZQapPNSvj6Ph5oSI/NlptXehL/3vbvNVYjmxznXqO6h+Kg66QnQv/UQIfnFBrIMjtMwoBy9kQPcP
vDcXbZZYm/93rgQ6LxLv/FNzxKTHOwG7aGn3xEkt+icq7HZXBG5NLFgABztbVuMeW0wd4X3Nv0+v
HVBvM0VZKdmks24FUKQNoLNPejQD6jCKr+cYTj8JlzVoQBRZcEomulypxdmqS5yaQnHg79yft0+M
iD4WkIP7n0eOAEc5ZWLKs+lvrmGWLDslJb5bU3sM8jDgraUT4ArqGdME/JJatw9953ZTbADKtlOt
o7F/AZlxYs5Y/HK9N1co8yx0CLULKi/I18yLTfumjKwTWB2HSshwREhN3QmFQacrr07QUF/RIVOK
YJA5Yar+XIZUcOmZZd+Avp+YSLsn6fyArV7kW4GNomXXdTvfNTMpZrRUHYR625g6HP8BYY85//BR
gTwMnff64JDq4jD0UCUUwg8QbtBlGjCnsuZjVkN8K3PG0uLbRl2Ze1IB7KIdRenuag3/TDNTvM9x
oyo4CiP9T1wcqnG3+dlc3z2e4sCPFT0tOnEQp88c5sluSPIc5NOVAUUnA17AskdiKkGRud3W58Ly
Z6pcWUMJYu7lB6JDxfb7XT2q0Z5GSyLSQigOYIVOcg5FJXrPRzrMSk7wCJsMeaPO8yNDXgvSe6B8
+lUCXSSjhJ6OhVkgKhM8wxqf57Fl9br4Ofsqaas0oBUoyv0i6dZGONWhZga8kNIBIrW+ZdXLPxyf
Mf5JN2MZGNpCpSvilZ2ESdr8IyGKKiBfrKfzUPZsdJLfprPLUVUlUkvc8w5sr9hoRXXu7bEnqOp6
rLnVummJFKwyXRBO1UgFzGMox451WlMAlxukrMjtac7kJChjob4nmf1n8ZLCgC8NIJIvFpCt+9b2
41tr5xAgUchmCZMdqxzupaSec1jiBr/pwQFfgK1YFcArmwzs/U3qDGPLSOHGxUSxoO/fzl1eLAR5
ALTceZOCRicHu87vIplEtcftgqAj7IKC1jvh3SRSTGPEsW7KMcOJ6w+YXnlwLHgDuCsDOI72MPzG
Q4ek7AvRpgdJgflscZZ6Tu12E9U+JEP/iXD+pd4S2lCRCs1GqHlXos3Vxwx5qMLVIePJ2Kn/PoZM
oCisan1+nD+12NjXw6/R9yeBcBChTiFdp929u6UcD6E2iO19YK1kEUlOZYh+izJOgwX4Iv/zSeGC
mR/5WiWp00NrlXGREf/CxXxV4OQliiq4jtB6QL3eoomO9VDrcPBqTHt6UeTMVWQtRjYHBaTktV05
GQ4NCjpM4Pd5p+pn7WBZQpTzfTI56NQT3mGQDc2i4Q3H+o+NPo7kMovQQR2UGKDWaYHjxSNsgmP7
uUfJArvk5rBY9lxoW0OyXKbmxKkUn5299o5rJhX6wAhldng0IrhpYW5zDXGx1/qBzO5zFTiJ5uHu
P/3s5etBRjwdk/YxQZ/E5siMcCnlLTAF05+HsZqaeekHcYmM9k8g8ZZmWOcqorC/3bWGq5kwU12+
k8no/wjOTKRd6rtMLR89GU7nJ57GJkTA2F4OPnuVIllfohar3j3veigfWWf03OnSpnWHtSnE6q7q
cKKVxUfNtTHflnU4B7vRdhjOC5Fol8dz/c72ZzvWvYtJjADa5dvCG6S3D8ti1pb6OJrmtgba63eu
M9nZ/D2kMcU2T5xea978yjklEDd7tJmwqRMzxdZ27tMA2Qff3FD9rjIwPelPlbGr93rEk2q4h3go
hZrvClyAi3umf8w+xhZTmn2CZqlp6JG7T6f3BCrKB5AiX3cBdM1DXoBdJrhnuwupkNiwq53pSqpO
XlM1iMbGDoF2bAerv4BEm9JHNJWon8UIvE6y6K9uSmY2CKlhg5wKNW/nQ0AhCMcMJitnMDGVpCq0
Qg/2E2nI2OsrLMFpYanrizIJb2NtQH0/fqvOdpZ8sIDa4jy5t+hah8KxfMmxwxN6IA+Jtp0fM/z7
PWbUfeL9yPS/jwR4HSgmYbwPxepkuza8j5BcWQlc+cQiSN59poGMU8GW/NrZGe/H+idKDzzwmRFL
LdHsmRP2YZK8mTLH8Av/pV37mwcP/KMSwcK1yLPkqr6Hzmg5+0CavBWqYZ57Y2cX62K2uxJtPlW3
BW5ODtrUnoUFikpOkkjDcSr1yFSekk/FNeYJwQ5sKPgPW2Nse+FJYi//d4IJDBqjeGecoXxPE/pn
Wi8GlOQdHZz3OYMQF6yHsTGevAqOHgDT/eOTC6HwG/XLDaKCUcZqbk4PZOt5Kd8zr4Uqp2Nh9yil
CH3N6T5whmRBu/3PNOzkqjxL+IlM0Jqc4TN0wSNNSECW1ToTlKM5mwHUrPqyYAFQtQV6Fhu0XaHe
DR2Muo/k1gNcrid4goNCmyL8Bv8Rkr/joRvwF4MV/x8oupwmD7ZNa+UWV3lZnH55TULH+JRXAaHg
+gkY8Qo8rvk40AOYOGjfnAP8lEw7HFZDNotpT/7yVr7POxP61rPNrF+YVtWF1YBO0dY+Wumibvi+
u4c9gTOI+gPyeg7sOGSKk/ieGz8HmUdw+muTowxoE+i/V7mwnexO6tnmWTcutmJSg16TzV3o1qLB
4bYdt6D3WiB49DGaIeUHS04yeEaNT/SmuGFG4JFsDNx+qMpSYU2S91PEHnUNQYmyYi/83Ls2Hr+U
DkiX1HTR6wTwGBlTLEClYi2mpOa/5gMjCtX7UiABzHyBWeF6jaqGv+fE/irybqywCwQRbqNXzbzY
Er0rxJw5sazRNZfvQ1PKJXCAP8pHopu9fqNHCf1G6BSM09D5LHPvmHydPFVfQMNxpzE9BPwVdOV0
8XlHKsGbrhb+Z2vysoqjNmvkIuZc/RpSCWxhSRG7dSbPLcmZkwY4k3C8QIxjTwxKaZ6wxqD4GULo
eNbJALg2iJsK+MLcCbc110Nxsjd4aliNGDwVntAQ/sU+JsL0xXYA3DnM/c51ZcY1im0oFM5u2WXU
x32PSVTrnuoyb/ey4U9fXfax8oSb7j13RPQAvAAtpLHV4c/z2NFYdGsDjekQzXUuepF9CalskpNj
thCezHX1+7PYhEPLPwX+YzxV7r+YgOXpc9lqFKPr5mFsGaqMUGz4IzpnMHnLhHTx5mlYTGXbsBEc
zb7ibcizEGyDsmfGVNi78gXAFT/avLPu0mGLOO2YDPW98BkmG3ZWkajMl3Jj85WQwCr+3y2KpI9i
Kq6m/EsK05dv1n700P18MXu5wke2DVzF/GM1B0bb9/V63TY3CLuOXXw2qG2riaah7bCCKIzjaeVU
RT9gjn6l4HdCT5qRJ6VsI7Aj0PkCZaVqlXGfeEvsNzSOPpHlYnGYujBRQldEH9n5zh/z1NIJanr3
4gwDbyGwsVSgOF7CiVwabdx5p3nwUKtl49UdlOYC8dIX9Vyntm5xOqExZVCW8qK7xiAFrUcG1B7d
Z8X/jEy5TCLme4uQ5Xx1MBEoBmGZlcCackhYhpo6q1DxiSQ26BOw62GZ+Ty0UmugWV6cJErIVN7t
diHq56rXsdgiD0kH/8JwlpEL1PY9SNAQQKOdXg1zeFvS6lotOzSXupz1ebhTLz/ONBXWKfNqTpba
Ixp3EzI14pGpyK7nPCQitaKNGGVMhK+DItXujFkUHcYfLaF27hdz/vfnDBKw4LoN/Ixx/suCQ6S2
MR9+1MxeTZSbBQm3YZnlE0QP+PbvLbATjO/NadcMIkJkjtaOlDpn1fTb1CW/IKzA+pQU4cmPSKIo
YRwoNlnJSbIKMRVVzsUvVV9ccun7i+l3SkyMbncLnB+3tZDJPpsGrQDz49tG87G+ML83QkEcSnrf
r1IcZ1aTTQ/qeV8Z+KOQygfpL8H1D4p9AFaLTvxGpeI/TxLJmrof/CdY4q5FG5Q7B5RbCaO19tGh
hEEYFPTvxuITTg05XWznAQ3D9dafLpGNIqOowgkYA2+usi6t5xwwcbhf/9njbVYxSSqAYW5m+S3u
L8pWkRpbmkjhTb3ZUVlaN6RMbf1ftNN7koE4iqhbANu/YQDzmNvlTv+N6PE+OdPdjnjcI+ea3UVM
TGNHN3dcoCgx4azjoLca+VlRAyzuXMaDnkzagDnXcz/R76TdRG80o1d+vl5gGwVHZ/s3W3h8blMm
FFPwwyM6llycIWXDaqauM34MHmGDvUpyhpS5Yqaff3bQrLun2tY6SYBLDjLCAzhQC988CSjyav3X
B2JyZaq5CvUTV5nr4DzUtlhkOfF38tT4qoG2EAOsJOFLVnzfRMDRm2Z+ajlRfD3YLJ+1jj1sUgUM
OMIbsUwWnIYFWWmtvz1c93cR++qe6hEH0pLnWnhLqKclou4b5WP/CetPTlYCq2sQbbRUVVwEHz0E
MJtFX67Ti5SiOIsS/vNceVlafpPKSG6AEc+Wge4KcP2VQNxqLjQgP15C0lMlTEfgI8qxQE1FjXiw
tAAoY2BErSxWFrS3P/rrInjW7nx8LKPaqgzz/yrldrkX5j47l32joKiKzFnaerw56iGDojY4K9TS
Y8Es3g99PxVvVBnx3L0z2xPOHf4j8BxTXOoebRoLyP2iSD/b4tT9Xae6hGxEaEGGAwbMXLv2ALiY
YA41tZJ/82y921TdisMG5af+vfPE7d5lwGdpBJpWdO12PQez0NBB8aqMSmN1mIwzFyIEmAL9Sblp
m6Ir5fo5ruJQelJ+rtUcOW2DR+1Q1PcAe8gjX6mned9szcyDSFEz/sB9pwxlbEiDBC87EreP1EKs
G7uYdEO1H4Y7rfsu+jiu0VMRmS2VEUt0IJgQKea6iy5qXhXHw4HNgOAbFnmqyRsc5LI9IKXNjoUk
2tYRmTN/nLO7GzI0rChusczAgMyIYv8iUjKV1u4X+io9L2afUflXqwI+QXQEfQu9/iUqJORU4M/u
erPSr4CBeSakWQLdKqLs/RpV73Wfb3En995/xjquXbsJp7zm1zYIbJWsVx5hvkNiZmFrCUEoWUEL
8dqFDdhqfoEu2GeiA5S3/aZShi8JH7pNVY7txjm/jzh8VnXaX67azF/04xiAYe4d8ORydsUr5Dqd
AEpba9Zxm544sjAQW16eVynKseJ1RW3hrdYEJbruJM++0N95Rh9/WrA/GK1ZRZIeaKx6VXffbMgS
CeaWdtoZhl+mtFYtErn+WALm+P6paSpUsFK3HxG4TCtCzUYfpPdHF9nPrWHW1O5DWQnWXUtYej5m
OidSRG6vQzXYKmgCfFzmNGcj741WYGCzEk1ESQP1ACfGCp1eIsVwKIigjVmGaXuVYp9IC/B84LbV
9+hqe4mXcjE25Cn80U4pmOKQMmfFNRXeupl2FtGG4e3eORaWyuS0xLbCUfAaXerK80DD1LO/KmmF
rdKgFvxilLMIKrNsIDGg+j5wH+d3Y+VEUB/cIUoajS4i14e6PrNUdU9LwEYgHFU5FlMGlbmDp9ti
mHy/xJKPZybYN4EzSUoLCj9oZWuVwfe0wbivJgOLupbFwjldvoW7AfIs3/LZlx1Z1mDnagfEy8OI
SiszFSNxnnxv3MDiwl+e2kGMCeTOd8jj/GZWRF84jpVVygTwqiAVPWXf0x9Zce7YkpIFbm5p4dDA
bK/299+0leJGe914is5sNQ4gNpQo30jJ23oqoaTmYmpCq2cBka2F4imZEsRtGEq24OAYCcJSgPiE
+Qq9OLtN3JoOF1AEVhH0v8VzDXpjOUTJodcjnr3lwb5rMMh4/YcOT7faO7jpumGghyCIndRm/IY0
eI5IeJi3DlZ7RXhHKlMUo1wY4jNsCleHlL6DxmO/KyXU7QzBeqvBS2ovZam10OveTpRtBiKUZmbb
HK4VzBTQpftjtbwDFiE5WIL9RkDVz1ECYNGbNwbOW/cFKgYfqtHMupYDs0CGFI0v3/gKZnZ5Y2uk
cGAVapCaNxkjJh0SnF2Iri6ZRfBpEZnStEzfojdMc5GsUyVNY6QZXMS//TZDHCZJBS1wlGwENRl3
pF0XUxXuoMdjAnwieBDd2xsiteQV1PEEiwnf6Xd4O21F780yYjJN7YaaSpZPudQ0N0/0I3mFc2E4
5lAxLdAGWmOe5v277SdQBeYb/+Mmsxw3r6SCY3b9uwFWbByicfYPj0oW5ehJkV08KrfeQQ1z4QiZ
MCKGJSDtViIEszFq4Mvg+3obZt2ty4MGtm7BDhKc4aUIGcyS99HAVBQ90YhsxVvBS0DQb40tqqLt
zDPL7+nXoYbdqPKAsfEFJpOe5W2ipxsaWRiA/HgWuU8ut/kYhmUiLAvJ2agQDrZRCG8hr2cE0+43
4U1/kYeT35Fxe74d4HdDYH4p4YSWtgyCI0qcb60xVs2srqtSgrwjqrIGuAehSRBIeEL2lkboiuB0
hJb+XvQkd7tc6hHV+7ovSyUlpMGLrKvzU2+n1hMQU506Z+12R6arMIkYER9R0dFRKOrvpdPzIC3o
445FV0e3qSgjF1uXmzHQk4COgndQOKY7TCuPkA1dJrQJQOs6Rvca1t+CrC0vbhKkY3Z9ra02jnw9
fglDZsEoQY+kqRpJ2UbNXcwO0H71wa5SmvpMMhgFOJF1qv4CKNIlsULRlriOSR2glZQoQ6WrN3f+
BvxJpx580uJkVFJ7pFLLVcLxTQT16256qgS0kf6f24eKNrnyCZgzn1ycrpYofBqOl9jIA8GFReLt
VPcmZevTjWuLlZr6SkRupaouEdtYuj7msYQybqA3ujYvZabOgUhXqFa8XkmSUEi0sQEvwL+MGx0C
B26Q1fTYywvzB6UTz257R9gUuDFIKz1zrvYMDDCviZXWSDO+1R5T/rDapH3FporFc0OEBQpK1LF8
weDXUKLQk19Qs4NB/jGLysCXW5h1qT3YDJKW4i0f5jzVItOiS0Ue1+lxDYYzlbL2WkPT+pLinvrB
vz9PEAROIGKbZNP1hzgf7+bAyqFw0x32Qf1gbdYLPuszVloCLfXMC4xUbjSsbRyWNX2T3r7mKmml
DE1FOjo5aRxJ6Qgc1KOt1b8Aikw/YuaI9KpnreqZiyfTQfMKx/oMpy9fHKCqqMKY2UYwuSzdlhjS
5KKV7+TxA1tgoS79HYnNvnstgmvMAr2woILJLilgWfS+qveM6OOQiSs+5V7MEjrTi165toB3+jYi
FW8/hPgN6vMFfUiGQF6/v52mboBlV5vZIddCatY7KmwoZioAcN9hb2e853Royx74YYNH53spzIsF
bEU1eaSe4FN/C2Kax0RlLZruYYgTob4nZSu7NnMa8VebWFDOHW2c3zxH+x299gdOmKrEvB3YQYQv
n8FkVOvY8Ec4P+w8uuw8D0lV1XN5Jzb/PTGewSqaM9SC7hJwdl3MHluqJoSbqeRIQ6mvB4a/bS0m
rr9Uytc9DbUZx4cKgNn79k3nKhEdKNjv5oHYG5eAtIKz9bI/Ugbf1RH4xoc2/CSbxz74ySL29fH6
072G66i4D+Bd8jk7U+vUElmeZgiv/rQ8Tqic86mmcv5wtOvPOB8Vpqx9TjiYkd65yPz7jDyVwfea
muygWsupsyxKimReFO2uliK9iyJQ3Jkyot1uD17We0Vc2ACgIruFpx5U+It1fofFArbY+560TfSn
djeVqwFISPagwCzVT5qX3pXJVJt/GhsiMOt0vHAGwKRzp3Zba2TsAIxO5J7dC1RT3yUBL2qhD6s6
b8jt8WZ31pI9NnstWtx8R19jRLVxBlOt0XY67/xidXvNbhkUpvUviYs2r+peGVGLBsTQH1+Fr0JX
G2EWqewH7ZP3//UOryWKXgmkROh8oKXGNUsRbkRXjyYOFe4/RCvJMQ4Zf/3UQ32qNcnxNVzcqOON
Yq4OLxglEVhrZGvRu1ah0qwsvE7Jta7OMCj7hPkHOgJHFko2C9ncYPqCQPjQG1KWS6JB1yC5EMBj
QRQbS6K/BQ2qA7u7VX8zemEzE5JYF4gzrllgdHy693yeB0ahe7ZKqgcaEtfk7Zh2ngHwIhZyebKo
+77VyHRWxp6jjbVmVbm0TgWGmPuG59nes/EnVCy9UIPwoxltuMovE7TvUsSGE44DWoVixjH6VkDn
BeigD9zcrmPz1le68nEmnmI9YCFB9/nBCnKb2ViXtajNoTbyzbtBUASe0hyifi5MsL+m8EpBv+3s
sEYzDMPgcpfFo+rXvr1rurk+iqGjjYMJ8Jg0R49eCVtudAO6A1OwFEYCiAZEQZOs5vBNfjW579yK
OBTWckyA6Sf0NYP5iu6J1/h+jfkLrqrxFHDXJhmqqZC42Jo/pKcsqFmIuu6NQ4gaAIvvAhjuM5wI
35rFwFY1hQhiSLAh1yzOwAHt06JwkTbTcFsi13ueCpnBDmNBJjy68rEO76+gHDQJBrN0pBr8DI37
+c/2xBO2jbsJZKkO/nfo+vfdh7um94zlWQnSMs6BXEUKgS6BhmQwwdUfQUlVYvS5fKawrCD/b+42
lJz1+I7bFHMJHK0oPzWxLrGNQfmvn/C9b/AftTVaQRaWCo64hHMAqjIiEeJW0DQj0cmWl3eFIE9W
JHLBXltf/JkGfnOEeS6MmhPBxJkoMo+7n9H74y5k6Z4aXycbKzxBrVIVQhYUOY1w0FbI349UoX5H
kIK7Vh0YQ2P8s59HUGP8KmEhl9sskvC5zeGa/TG+LmI8+tpzfNyGsXeN4VCPvr1enLns8BW15iyp
4e3rZ7tsBE6l0GNC93iOsovSK1c9oSoONgwoRjmsB+k3xwj2A+R7V2uWZeNMme5IP7dV/75NP6+N
zw8sgq/WPzlsxdL40AC2VKFqM602yrqd1tsyvytokyHoHdtpzRBRIK1VzR4coIsuw22n0IoGNlHz
S8p7SmH3a2li2SrRNkHwynGH4rbh3MJt0wt58/iDLkfkAIBVkIHIPk+8cOyH4FCmV+cMxmXR2M6y
zGMAm43s92lhBHn7X7iK/PHEXIk8e5x1AJpIMUgLA3MD96vWK74uEgTuQRotTDLYYGUAYE1RYdPs
e6eYj3YBA0KlH45BTH6RjwMSV66Qr/G/rn2A1vK+onl0oMB/q3XCAOhGJTZu1oknnaq2dHsTGoIF
oCpxX4A01fXlgLdTCyCX4vRyJ4NlR8vNN0dRXVv7t9qfjy30zuKuiCzF5M3PI+PvtGqFUY4phyJA
tPN+3tv0RVgEmVyflNy8rqqUTiJw53JvmK89g3wxVlKa3IbsgXKXLmiEua1eRdv/zJPtRWzesux4
agJ6PvEVVaZsqJPBdLz1SogwWUM0HEHm/sXssHBCh/C/9utjhDZLwUIj/JXyqVeyIl+EwFPlU4tq
3H8SA4ZaAS/UFXoB8zJBdGOEVy3grDNkhO7QwwLm66IbGf17mrNaIPnN3t/qbKpHiWvy8rXIO/+9
v/PWVAbfdwMjdx6o1ZJ8icxL194V2LL0n3LbOGK+gS40CJWIUnH6SINburt2hfl4j+j+hMphdImi
lEV+JteJQC1e0x/G5nc55Erqrp9NnPl2JHByWmJz1ZpPORT4fRgQNM+miw2Z2WP4YN2zSbFoH01c
ZV5UosoUxqijgORasy/Rzx1k5Z8VU7J8dmCg31Ck3CDB6EeFZVCEg1F0Nwu0mwX1x3M/JvoYr6Uj
sadONkjLLSOSWvcIIDGHMg7thyl6UutQ53Hw7Mi0po0fPk8C/qiImOW6hcIOLxpmElD6vsuxBFQm
PuWzQE3Pij3HtbfFJQlbozbMBMjey98xJfLSTHfZmJoZKwvOZNlGKgrqOEfYn4S4pTeuvoRieMlz
f1P6UnS3pmoIQQHHMoAWpgGALD7eNN2USDcH/7TQVZ+emHgNHzpNSH5wNtwvCyRqVUrQ+x0NB0Bu
9GYb0CI91Xtraovyv732gUXRfOtIYKrp4LOhAKSEe1cbXoHfQAs/NFvYIYLqQGe6WDSW4Xwx59+0
J39hiPfcH/0gtmCASbnvtA9I4lNVziTfl8wv6lYR1ep2zX18WMay2t+nyetGfkVowaET0KEDU8G+
p5IgKX5MNbBlhIM0/vljdwmQqJj+YYcrx8gskEPzhqQBzWrjjC4klaQSmOh17+bWW9VzWMWD+ay3
L/Tb8M1fTRtNkPutahN0+De3Svrr8Qz3g+dMnLURKGJq9E0QyJmA19a+zEflU+a+i63wRBf300d8
xp2evgBOJuOqnC40ALUtUB8XHeXJyWzylzfqOoAMXNBUOeb1b/i7WcbgkXsjLNHkUMyOsCEIjVIb
CX3Uc+Lrc/oXgPAOdR0Nl5ADCglnRNx53i/0MM1S2tByeVAUBvdbWLYKeVteruYhThh/1VNUO5t7
KpjKaNUzuUgCfis5rBZgB6xoOJF8gpr6VqQTMF9a5SpYEDmN+7gSI9hj1sHiobDtykNterU3f2aL
JWh1hLT+4E0iyzelPzBAkoDJ4GaWSdBbB74FAKBrmF+hdjS8hMgowgI6yO1K92A5owY1MQ/U/LiK
T0Fr/4rzE74fnSW8UpJKTb/XZ1cNPL9AVVBgBDQA4M9acAN7ytx+0HoIZPcFmpmimyPRzcNPoH0i
UoNOyKY56GCwgNDA+Sa5dGxlXMCjguPh4bSlcwNjwOfjkCE22uQnpfpg0Sb8EyF+017VJLkFaQZm
zmizSNKlY9NrmT1vFOOuAVYH1daXqKT1ont7rwt9ihhpsJaLXlm6AILmkeHJWzGvbZs5vD7ycRw5
kn1XxKMRAmCN/TfUVYzdEHw/mgoAFgmvo44oVHg7lZnqephGsdj2ODghAOzzBV6Cul0L1KmNSgat
Yh42KYAKc1Yeb6GasOOFASl8h+sb9lXmx6LyOLcRoPr3adxKGvHLyXhavI04YftCTn5FOMNPws5M
plJ8DmvZ1IW57DNrY8T8+m/WD/t3/ymVZXrNZ6UO3VfKymdiw2oQctzPhxpqcsBpr68B68ddQHdE
rA65iDDC1llaBTjtM68qB+rsw1/AQKtaaiDZM+0/H0dGecLHK1DNdJqk8fUUnlng8aZCkodzt7+6
nng1n2Jnma1nEehmb7IjjQiu6BC8Qdt01n+C73aYor3eD7rl6niB05xHV/BQmjOq6FjRxmlNzh6o
LPlvyuRLcY6gcOT3m4yLpElFP2kcZDONMpVKFxGpzIJ8SlZlKuiJ4GWzZ1iHjPWxCmIpie45U2Nb
MrzPsKXD3kGX1s3916AgywAKK3PgHO6R3WwLDL9ix6UlKjTISNx9o+qKBDyECa5szd0I1rSBKaS+
9KjbXg0yXirxnfS5aFuuoq0yG1l23lMHJt2JuiJwNNmLParDaiEFbdfXEFTQteMW7Rqb8GZJ+P2N
KiqF6lDD/prTcdh+Xf8b/7eOUt0usojjqDT8uHRqHgSsuYsQf7tCWn5L18GD2XNzF+cRraYVwTjU
U/O0VTIYlEMiYFHNd7g+v08kYuxhTcBzQBg6l9wVCKXiV6fa1+jUmMv5te3CTIRz7+/MS4diIKGB
O0SQ/YPR9qD3S3CeXTx6KaVA8cygp22eDib6Yrv+ePuZjqLWNzrA6Pdi7fd/07pVTcx9y4QP4o23
3J8GY6QiznE6XszpQXw8NelV305qQGlh3dFus6LEsPvOru6VWbp+byCBaQUPuD6wumEo1jvY2XvD
Q9fEDQ5pBecZRYibJGNnU9S+TZZbm1AnwC2c2BdUdGcibxVueC7UJJKIvi+MejhvplLR7T9XRrGA
yvEFf8smRFRA7dLxj4aou7nm86GexhXwV2JSJd0m7jHZN/OXc+/swQTYL1BwbVD2qIrRkVTsSYd5
irtc8aCgtzwm3YeeeEPsmuX78E6FeztQhfxdDiIGckJB8jXbd6mUxrtdyzFAf9QNzQ1q52Ew2pWd
KmOKQzI5ghl0x3RykiDCNFF66lvwfQewELi0tzLp9cwYjF9N0S3hKCxDhTczcdGR/6dV4Tz88Qx1
pL9aPOnsUl2KndJXXhmEV41Cwwzsdjt2PYIB1+4nsrvsZT6VAK4CA2S+LLLF+qvWqfIAq+mGkEIN
GLgJ71fCt7T5aKwkMPntfqt5seIkpsP8s62kW1+JaaHEBihtBVNOgXgeS2BuGF1Y4oQWqAsbKEEK
lMvMT7BYPfjEXPF0GAQPmxepm1o8PltV7vqzpy2zj2rlteD/l6hSEjSMCvyoEQ34tL0SXu81WIfX
jzqRgKqryoNvmq/4TW67TOP2Y8rwFTe2kUAMz4iYj2iS9/pDUFK8bclH3VLqyFRY8S0QUgSh+JPT
SYn8O4+sRG13ZF5PFBUqe6nKA9k2eAvEXkZtCdA52pWUAWdnU7tEyxfyaBMFyThzYnnNkWfiLL3z
RTxPAujkGsjnRy6j8z7LWjjMIs7O04PDFAwpNgmzEcfRU07nwKMYLni1vbaUIhfYScxUY6dhpssA
iwLg+HV/JHuUG++6O2BP0aKklh1R9xqjjTknL6JME7f0n9X8TZwiqxhh218rukUm3Vi8e19Umr1F
hO00QZC5Q54wqU5kzLno0n1vC0o9bLJUZQJWO2QsEulEomQzHe4Z1omz/O6DxnjPYr5A4miQDUmz
W8QsiV1rIv7WrmiHs+nYFdXjGcHikIHnlviJ9BOT6MQM53su1QjR1yv+mW8CyUe7kSRt4cHEsW51
7cBIGchDigHfhr2UTqsbPZD0HHzYajYJV7bIvxzriIiaUwNkHpdpxIgtZjOF/BziyTzoulro6SNN
G3M6d0t/n5IcuYaOde8r68jpZpciivcPZmkNjzsR/ws7h627Z+JZ9h6EUU473YbkeksPEelTGi5+
1UHdylDVCsR5q49Vw3vh6Y9IXmg6G12xmIBLFND1wl8lr/to077Vl5K4LgyYixdoK4qCPqCNERpC
q16zQp5c9YKPphYpwumX6OIn1DMhHxdreZm08Qoq9skliEK5PAx3NEZtMgFmVX6dWQLYN4XFB8ts
bLf0po/6lnBDpVWANbn3mWvfpwLniIdkeP22tMh5POnu+7YDm0NNCGMqCziua7pkYWhhqe6uyAHD
HOd+Pu3n0tPyQId/v2j40WvoGIPwZ1X8HvR1qm2PO9B8bOh4zbDrR192qRIoFGxpzqurP10G7A6g
gVjB3sqC2s+4LJFQrrCfoaqy9mPk08N5YqVu+QwbvW4opb3uzfTef63knz3U18Y1gWftt4+oLL+1
09fLFHlhPgxT8MiAOBkU/j/yJ7aFBEfR7aNgu7lNEKvXZv11nFX9TCZs5M4jVwSvbJLRKFN/mnLD
X6gbPO78ekkBHt/U/M/KWG8I3hG3IjieYKrtUicIHiWg4gg0Iqb2buOBdmKZ1Nyyjucd3Gp3x8L5
JBh1iXyvou9CEaScdxg+nx+GNoLKe4EBrCYy1FoKadwMlJ3RM5eaEB1oyTB707F9/PkigffCCoI7
4oNW+NFuytZqVDoOd8RuQa0B67Njug9OGV6A9flPMpreCA+OG+p923x6zZZHO1VOLhTy6dgsAmdi
yB7X+lUvQNyaKCqZHRxmFi/1cWPOv18oNam0kDRFXDpvWipLjWSjU54YFFpk/1ZKIMesJ4inQYOq
uK0gphHtStfo6vUXxxZZY3qXe/Fi1VO3cew8s9Pop1TCh1Avf4f0Oh1k3Ll66V2oTUHZai3ExFJQ
3rRJjD+Ysv10eNke7TM2uswWlXQuvzPNY/GZKzmsyOpw0FzweAdenIuwbbvSkd8VezNJwJRg4jph
CdoTYXJ7bGO3goTsJ62i1I6GcPYIAl4XvMqywug8/0psDnVLiuWm6LnDq9Xrze3vmhr+G6RgoZ5o
v3mJzTWfehN2Uzkh2GgsXjfG2MV71FROuAt1wq/uERNpVYw4YmnlHQUVLu+zC4e9eliq6vFhHHVg
8r8vpH8Dy75nBwulDtBazao4Eby0rz3Kav/futjmCXGQvJ6yOPfIGX0YrgeYajIIyfc5/F6PWXhx
/+WEQ3kxLDInnPxDrC+g1E5uJ082sA2ZFfOkIxb1HdPQqf+QFsZWRIQndZR+kYZMuZOjD/X3KNoh
6NTqXfQ1RgJV0CAj64aYtdw6GbUiaIbTriDvX0paHhbz45jU56bilrOcW4soaoNH8xy1jH6mNIyK
sFvrEg5+xq2IWDTU/L98bxviArxnQ7pRM76XTVbFytUCfLKhS/WzP7jJRGwkcCoorfan5ugD4O30
kpjzTzsj9M3+3eoqwOutHPeD5TH9JcIKLynt4O/BOhsBvPL/CMoiZeYXGg5HnSAIxgYiu5os8Juv
NHbujHA6Rro3BXoYRPKYQoWz7hFZHYpoPorEArlwFwlExPNjgIjigzpny/JRUT1fVmf6Awj+6OUR
wvRCaZoxR18S7yq1kTUOema6NDTKQrUk5wC9hnVsSwHD4bWGL2LF0i72vNVLnJfjLpBEuoQznOmR
QyHbj5Ji95LdsOXZxThLYpM1wrS+oTBIInDK5Eoz6/TIOgp6c05GDVb3q3+7ohkMLChB81oXcq5f
sQegpQ8lVLXE71S1bRbcjFwgd+WCOu/GK76QIaaMCNKozHiYrCihA4JghyfNwad1E51Uk/zXMJxQ
9njXu9vuAU4F8xi9N6XQ7w9WiR6VOuSNnPCaIfYBxXRO7nCFRLojLT6kl0ATyuF1x3uiamhK1TC6
SIjnGlffma5T4Bit36xz4O9HCaozmrNeirqEmLJKw14Bo8VYNh9E17VH+U1VGa3j+q5XblZ3DdN7
oBGW5In3e1WTKNOimCJRH3UKB/9/6HdqMxZMlTAJbgHDwVwUjDSqnKYXCaW+qqJhwKejG9zCGJdN
CZBe3FzYM3KhwFegXRgMYUSp6fV7/ogjbTGgnKsMzbguSh62+YcAAn+c1IW633pipLnmfKqz7kUy
Q9FIdQdEfNPamImRdRH4Mo8ww3Czlu8zRdOVPdttcjw9hiTYULf6R3JMT5kRVnYA9+ItQQjdHmsq
2CVHKWc/Nrw7zYG4M2vuT60StJmQ8uV1R+cJjUkGqRS6SKCy3gHM9qMHHbd0e69OtcpWktjqycyy
SP9hgRrPtisJ2+jSE470oXE8bYKKdiKtP+XWtiTlKTALVM8kW5z82V8OwQbuBJSJnJ4A+o+cPimA
+QaGBvRmVWEMymNAjU6IYu4psZE5kNAof9xNYzGMPfqo1WiBHiKh6l0G9pBfA9SEgA+rgzUrQaNW
KODopb0lc+CHmyDV3MYhhmQyu2l3AsOtdy+PL0Bw6xFD+lM0jxQ21yNVcAg9CiUg24Km4t8Pweyb
gD34saKo2Zx/OthCkOgyHDmrPEt1/7HKYDnziygVWUQTR/xW1LymqtCamrkVBN4c3OJi0cBZxTe5
vhJnTOEUYM4vaTldE8PHb2dzIbbGpyrZvyduzABWJymOSenjjWTkGiSO0oSCPHAzU8jmGKJ25zPO
M8wcxkWRJd4nsO2MOz57g9+lqn2g6CCWNTtQT7Ps8lYg2WgzPJIIyB973uHNH7CIhqte+RDRb/r6
wnZfGArMp5f1FH1AalwOxNlnofX8JcGQbzv3SVm+xfWgiwpnTv25G6bjIGxYreYGUUvSjxcUCoFM
Uw7olBVgwgiX+3OFdBL0UJyRHkTJ/ssoQee+dRt6QEwT5u5MAaM9m2N7y2W7kz2yZfXW63elvT7A
//zrrAclxz+NksfOSu7opu9ZoSby9W34OTT9PlMX5kxZkd5bCWkpnTitJYh1v/H22qsa2nWmQoWq
/zaq6OuZ451pL4H1zZVSYKuKjxAtxKwgyupeermNlPKAdsrDOmXvOBkA27NQzSLSAKO/fKvrq1FA
rjSbbZJQ2tq9Ezo+EDPw20bqHXjmcExYXYsc2fgDm9RJNysUtA7k8jA+5Gaeq+/cWXinAWtiSX+k
rON22QoXtbsk70ogIbpH+4XINRriCoepVs+i7SfMgC18MSQaAbuGfCacACRMbP6/FVXrg1t4Y4ry
atHB4O2FUtEp/l4n8rLngTRbgen6hmIWF5YL+6Q1megNlx6DVEAMKZO/VEG1y/h9Kxz0S1xDxeNq
vLbZaA+t+QcNLsbZkD7qBdjQNRw3asqIUIzQSV3spCdEVC/G6JTT6Y5aWTNqVR/p1B+/S6sOFvyQ
dP5wWyQlanmOW4eqqoh6idJpxXwJQ5gwfIIRtO+ZEwp+r/QZ8QJtOk5OnkEjjlfB52ANH+72xMXb
n240hBETUZksDkES9WgK5EkDpGEtg6DV++YOT4hBramgGVWgzt3x1frVu63RUf1pjgi2UNBgPLCp
EBzZe7ohpOLWqS+i49uaMGc7hVZDdVKLpPp9vI0UwT1BMRNa/2YIuE6SviJnRZE1SaPuhvZxRK+h
XV/QBGrTSgn9r/75YonrcuNa4/pLcUBDB/OzuVCseIsZQ1twXw8d7Kea9IjLkJhP+pnQVedVt0Fe
q5h1SfNqbNDxREU+pvRBe5pINvDEERVWJhpLLhTS0A8FtwrPx35jm21P07jM3xexBBNmhZxSZSZy
VUAlH2kTvhg1nhmhw0Rs10VwgTHTDnfCp+8Unrgg5cJinWXbUd53USRm1wwCUbxhJnD8Kow6XxP0
MzC4pakf/s7Na6aY1eJGVQygn3W0l1RzbD66xiEJXUx9l1O6QaDbiawmspIWtpkXhiKFc/pNz33+
lDSTrZOP8eokEb9816pqDp0WeUYyPCGtG2Be1jJTu2PrW5eGPRHCdZxd+8DlKJ/iEQEgSPe5Pl5d
I+e0xhVh80csvDLRsFaSBhoB2BIvz4NC4RqAEevxbI8RqFxFsBywambGHgcZfvuRVGGZOB329uXc
GlnU1t/FuG7vxSIqp+bpcTmxqe+4vJLqhem/iydXb/mMInt8REzPo3zfpC+FknuY7eBhBqLBTn7O
zvRFZ2UGAxNrheRRCCNJxsHC81mNpbhoIszomuLIXqa4Rzby+LlTHEhNLV5JqFyjbduYlx7hMCFz
ssttK+dTRPu93hE7yIJfvg6phc6+BfeIp2O8l6X5pXl4t0vXO/2WpQagbfIoh7S0EQFtdoMIyL08
fM0S+jgVvB6AisYWdLaH1+SfYF0k3ovI1QrzLQy/UEdQVYk7bJETsg4Z/WEFChOPDgp2ImK8N5XY
sJOs9Sba1pxF/vUOU51Fjm+0Zzsc7tJ/ZOQUp0PChKlQaRiE2LD0ipIN0fe4XpSOP8NZgvI6TT6N
tDRrQ4JB9o4uGqooSyYs3ektU9rDt4OiVUR11OmgmeSnFUEyFX7b9mOzCtXo52tJ1NL6wNdQ9rGW
gln8aP8zRIbq51ucQ+5BtDbfgO7SYfajWFNHb5GEpUTZzPHSBWO9whLhX+b2Q9H6KkVP81IvRe6q
7y19nfAN5tZKvZgrNBgNkaowrynw6S51Sjt65925/3Kv5/BvNsiaqHxWjMpExyloB+LekHT62NI5
XQ5DaWRWS8pDnhcQWmaTV5TLUJwWqwrGgQJ7KwleSjm6jsU+CFb+Xl99cTAoSdWoFBEDtWKcKHJa
d7B3BFawr0gt1S4TpoOlMit3mIp8IDRFUXNL2Dt281I2zEXHyGDV0WID+yd1eHeHT2R5Co+Yv1yi
HXml3kWvq/NeTGAP0O5ETbPTOgMFmqK1ChHJf/sl1u7omnFXPoUB0psg9EI6bq6v0YZkyjoNzbtT
R7uEaGepiq0S/TdGGCT0Og1wj7yppBN8OKFdbv8y4c48qqhrfVA6TvAKaCSvwOyZqZpuie8i/PW6
yR9ECxvGnAKnXcohhSb8RzOFf+SA4Rgsjxp1y+yjFYIgqx5ndtuzGeebDEU4TuaQ78QQuZiYVygy
X5vKqxAGmBoQV5kypifWAza2p77PTTn0+aXGZrHr8Gpv0dNfk3P1EZ60YKRsMHsoi3ZvyKA0kY6i
DV1q9dG8dli/iAfwVHtxdrLJofQnLFPZEiCMExQVA17JYRVKaDmrXEDNCJik7KYIgMZWa7ERFGvI
h6k4svBH2I1hXwyNHROJF9MBD2fJ0qlXt4/NUgYX7JmbfTvQkjjudpyze3cKFewU1VN5+nD57D/B
K9hEIk/s5k4/VINTvlYyElfP38YiULW9mostmXgw3jJEdCRema+fAnBRsM/NmlFuI5eIMsdJzf9I
b9kEeHSA4gsx4DF71/a+I3AdI+Gsq78sih2JbkJSVJ0Y31/r79ah3QYZHMGtsZyvB3DU6RqYRkVL
Nm83tR0sRsnQf1LeMzwkM+evIUIJb//DoAdWs+kk8xgYfSOrLVWjZkTd6Fwdlp2JXKU7aMTlh6uI
E+B7QRe28t+Tj917pF1rQSBR/esl830c3U2Y0qjLnAghCLyZFRe/ld+qihCYZAKm/vKpQvpcd088
sMnsOQZ/4bgZY8ejfSMx27cF+jiB8GpK4ZhYXXOxDa9dvebsGMzWgwh5O2VfmW7GOaeolshZ5CpP
F9uDNnOAHXd6W3ouBNFYID1k4PK4a7GZzIFtHSHJVkSg+kj56qEscPMtX4rqpDIGM3Z6HSmmq7ch
ZPXOnAh+WRgjhjLP2dNpgvNKjOuiTxzENMbX97ll1PAPVR9KER5B3T0R8yTi2GzSgqnQkXRyTyTL
j07FEM8NvCqYLGMDcemF+ZbMEAB8szPBvkX85LEzyLyb4CrUtALdYEC6wKIpuzE7pe/wzXEZZ0ID
3OpmUSM6ke7YC5H7WKc07PV0eXgTimfDWDpz/U0tR9KSbMq6hArF/4R3xBJ3msjeqbHmlNFB1lW6
rdUHVzNnrGJTBm4lqZI2vJ2xl9bNwQENOtPeOyQFTOMAaMr88D3So1DzCt8J7xRXnqOZ2iQ83Oce
nsZ7KLNs7gd+uAjCC0T42+X+Ddpx8+TqEU6Jz04cjmUtHmlaBlD5+vDGROPZj4b7x1nNvxdGZsXO
Qfde8H/lg5U8wQJqqo4qXhqj+9rXzlAnZqUDASZ4vP0ByHoILP5n0PDtTBS/N2p/aC9uimPdcwu4
s7zVGAZN66RVfk343gC8LIA3tnCDopOR19yUM3pUYgMQ1N+QKmtxT2sevlLI9NRGqUeen0UtRRbH
jUxo3Rgf5TZKUI1C0FaxZplMR0YowLlkzQahy8n4TvficVJR07ubfbL+G0kE6fjt8g05LlJo5kv+
LYVAfsWE3UNWxvJjqdyjUUJvBRrkuw8vbnobiDOWbL2N3gFoxuf2aaPVEi/bIruiZjCN+6tydSdF
5pK/hFxMVJj/NPex87UfWxfRQBOSxplG22Tuj8kfS5Hq2vxMhn4UK6vQ8Xcnd5hxz4/l4NcBiLjb
xyBmEfGYbBLLv3Nt/fnRXAwSBr2HSLj6+CHfNtUvqHIAjGlOQz9OQ/3U2E4S2wijB6n3pOTh+Zx4
0W2Nzm3D92MrA58/2T3uHWsKZgcTa1gwAjZJKFF0INOCr8cAVChEx5bwWUO6yYTrtSoN0Dm2peb+
A7Ek21qu+QgLOm8u1CdkRxr1D81Tx5zSWi93rjGcsKlv98biiG+Bzr9SLHLrVLGZkztdoCplVt3j
9XaVO8S/yRYAyQS0VkXOva19ALyM4+AidwVHvhtEKQby4E2TyzcF7AF/JQIiZ4frh7JotLSowHmw
sWku6mi69NUp4mwoy+Fx3I/HARbV4GBTNCxJpixcW1oT6LNKcTRbEmtvPb2Ahva0fhwyMne9M/wY
SWPHnGAsi1DKYvfoeI0HVkmiPLvNUtPG+n0/cVh0kPHxLh9KEkDM9t7eUnQ6QwWno2EgR7sSyyz9
7OgcgJW2dCn3tYFQ9TocrKPzJVDpoLXkLz+vHJYILGWGM84NA31X/FfaTFYjXxERhM3uF7R4n3bu
wCewPdDLNlJJCXkrYnSK4/+VPQ52wMqRmflted6WkYcklQ9PyZvr1yu4BlU0jzW8m2Ll6xjnMljW
VIUvRj5VTKN0iKj28K6Sff9f0uSzkZ5uI7rzrimGuKcNX/TM2EYKFxuV58rNEc7xBqF5ORGU0ZoK
Noye9QrGSByc1v2b/xnFVVriFGHwAhov7i1taaT65hC8NZ/lnglrnh10w9DgDeX9D5aLTgPfHcog
V6HikFvqH1TzajGhpIsecAlAlS6QvsdMCMARNftPrNx7sIx94w8ok2DZz91HdOlVvPgaILThq1FJ
9MKRQGptlBFDlyCiVDDcKUCYV4s/GrbkZ3vTqaaIX1hjA4/N31pPeT/Zc2NjKaelfh5h1ivmPej4
V8h0c6D35rAmA/C9MNR1eG/amlv7GVw+Pz4AeSdBORySgXjb0uOuuvsq1MiwV0ahPkCYkBNOg1Qp
GLZMcePET8E7xwGHFRw+8xTIJk089CcaexZwyecOz/6jIX4pKcBRyo8dqDghGTM8haG4M6N7ciYu
w4xHr1GrcagrMnZWErdvsYNZEDbNdBKBgHUIkKAwZNOhfdvqagHcCHkMD0paWcOf1KRJi0FAdPkn
QonsHXwn+lwC9j/JcKHLXSJlwNAE3WNez1yBa2VA2sE9HxDdp4sZCplXkPEVzvLdBR5P/lvDRAi+
C2FSMXe7sVECEOzcm/aMP2Lf/VGsTLqizl7I/atSwipUgmRno/hhxD4Md05YOEptxl8mxY0VvcKH
GmYKCxU9PO4yvWMijoV6TOEnUq++936pL6KckjjD791+p0O0PQY089qWh33Bt5j2Dhr2S7EkDwr+
T2zP9w+W0I/ou7RaLF7dt3UYrjwL/m1I2r0m7pr4sfCj5B3fTeAc+1uc+AwakrfbNWblnVFhFb+x
pTrlXb1bJDFfZiZB5GMhBi+cGq91qLTi5FsIomDKItXZp3Mm+yF5CgIjbufYOcfbEIbUE7A8btWA
+h/qJKUj+oqVLudGG2RkaxoUNIeggqIeqjM3lJEJCj54BwPtZwHZNQW60afxeBybmSUAdDorLSXA
dEYCws3KepPNizhYKi6Pvcuh7WhG566UHV2TLM1VAWNzltIdXDTmFSWTdcdhl0iwiHudO4+G5weC
s7vwZWFsXsufFL9JqpVf+eaFSxzMLnZRafZl7daWtWrJgaRTGtv8J6EufTKWH7Qz5zf7///wAFsX
M9z8nlKMaDpuB8RipMFhI3X4NlzCPxsc9yDOkBEOttqhuXryzf3AKuUcuHD/2zgD9j4qZtvG2235
LQ7F+0Io+A5sLuEoYQkI+igx1eUjosj4E0IwoKwEuKA/zlbwWkim82x6yuqNq/Mb7MPeVBQjQ4b8
S/VI0+ziV2c0dqVKs9ac3Hv47OBKCUr/ZL//CtWCxVlaMmOg7ZcUDwPXvNPBrsOJHvOl6qciMsg9
ni1Zm3tSLyQLbia4eyjbWTJbSzDz6A2G21Q/yrDXmw44+shyyk/N6qBrI4UGxtOiYt/PGRGhx7fV
J+yao0qD5HdDMpvwXCiG0zNHnOiPNxZmY26gHY45ES55k0EcKSLt318dDrW7xA7xr7CZSYxYCEU4
9JJ+cJsmlO4IZH34q60KefeNYnEYKrPmtPXkpLe+5SQEgODN/KNUqyP66v5hR5XHcmOctUt+iLKT
c4yodV7GrCQAda6MvQEU2e3lIGTXfyOm8GE2P1BUyYvv2z8Vht3RNJeB1RjMKvngfDDulcrauHnJ
g/swo7CdzfAnOv6YMPTXiiFjjCY0eOFefB96VzSzgW96PmfDiAWlnsEose3VuyW12/HKhJY7WMAF
b2qwwJiZBzQD0TJtlaRb4YzSdK3KPlImAcx7vl7O9D/u+lVyPTNWsjo/qPA2cb0VUNINnQ1LeSZ+
c3uqiX744T9abDSI4vgRxFpEQfenWyeDRRKPq5wJw6wyFhzIe5oiPvDSnVFj7iN8tYOcQqQR/EGq
NoeAudoHXVcmwvua0gdQRFWspzZDQT/Oz6O47lNjc7oX4z+kHGo9f2DyvWlXHXR2ada/2xcF3bpb
wnR6IGxsSDNJuMYGHfh6raroof1Po0w7iafxmyV6Lz1Y3s/P/V5tdg+vrtQVcHusG6P7s75JQqiC
uVBfiQn5HpCYhFcoYRk4hVhng2CP4DrX+wOoQIf2m3OXOKUnboreNxmz4evSfD/eSMxFJQGynq2A
2DdBWirQmwa6gkNMpBJ6ZHpkb0v3EJGgh4FN4qLMEqc2742yTTRzl6ufT7n0QUtt3V+YxC5Wz9yC
EYeYrVKrg6ToHcd+hd1ku694VfjyWRxPhqLQaPdbNJwc0ahFpiJn0OyvmjvazPOYcSNPqkKlqwS9
eqtOe72ViLaBdDe+XS1MqKoAeEGAInD35pcHa+q3wnErJpJgylesPai/BrFSmarVwXSj3bhPzM1A
15Uw6tvtE42JC9j+F1bxMKXWvB10+FWyyFCCr54YDWhZOKTJJDLZoOGnr/i+fyYSI9Pq2zkGsHwj
XZ1MKNuj9Ralq56OBK9sVO+uL6KSxQinGLberh/yymKUkHiq+tzYhwtUHE13oe4SxQsQG2wmk9MV
n8YYJjf9TZ1OpzY58MCfi6/XKAk2INiRaiW7mgaHvlXDpJ6Tfq1x2dgBiKJW22uS5vvn/Vi46mzL
+VBZD9VdiDo2yUL1NzO5FkSdVztyoV8ogD4r5Bie2n7SwWZj23MjOcVc3MqUp9pDRB66tidUmMw0
MWA3TiTPWGqukmmjQdPNwiVXbfieRGwlmSuOa6Dy0igxDMiDJtvDb/w0Cuxov9xFd5+pQg/UoXd0
Ro0ImPTDyJX6s/5+jDpCP+mpPAz8yhfy+98XIpImGEWDQO1giRtXT7pEdi4M/6SMvA5j8NQc7uKP
suSDwP3WseTEEPXVXdMxPcP9BkY/L/3wdvTOBQKnhuRhR/prJKSR46DZnRA39KwDTjNdOSEBSopb
a5bXxlVDuHDtCxgAPZn+wXhVHmrK7QRjU4mIfAvmwozn8wo/KX9Y1pm9JxHbnc6OMZ4UnOYMJKJA
UnEFOqOa/loqTJ5yycBvCreOeVF9Q23SYtw38njH1f+2LKxYPdJm9tunTQJCOgT/SwiNEg0h8Pe1
66hUW8pA8/Rp7D+eQEPhPSc1+obLnrxLcbBee2xBEIYxxcvwTmZj+z5oeNmncOExxg9wwjKtlGxV
8cz8bVCgs/zasLk1VciDimWgcjUq4DiHmS5dgPqfu7zjYunXpCFbwIAUJEW60Vw4Fj6IHCcKWfej
KLanVemDrZVrspQkjl2ywTSTXyiJnwh8dk+qD7FU6doH/ZxW+LIGpRngikGaTe5+BddEBPSeaGt9
i2Ok6B7nXRLqtUcPB3YaNg4RU0UFIxsBwLic3YJE8n4pxkToH9c3gsNyLaWkWuPXs4hfOyntH4B1
PJwtxtoPz0mzfNF3wVSLC5ZBFPoy5a9zY9erUFhPKuNzD/+f5o4A0RrEnl+OlhA5hsohjCWnx+sW
mb481C8z8hmBueCnzVFLIiECWITVS2Pmf/Qwlzed4NguU9tAqACLELZ+4tbQgR4oemfGaBivWfH5
Bob4lDu2n+I/s+Uxo634KOkG+VcLEjOxK8BJanqJAJZmwfZWJ2XE/5/pv0PiuPzUs8aPolxRqmk0
vdttR4UeWEFAOpIK+kQcHGBVfybYVASEIpv1vaS8z92TmzAprm//8pun3uiT/qGvvjgP8UtoSAXh
2EAuxm0mpTjWR+JU+81Npj+vp2TmqYRVB0cKeXsp+8x/3QeL5bwvXnBM/pLpNmfLaKp2oOvA7SNN
Zperw3KfXG9jhd9XapzLPrN2Epy8yj6d20swlOzMMI2N1QN4pybRrDk/AaMpbpGzZ0s5THZ6UtB3
rkB5FxA7nGukdcG1VsPhMIu7eo/xlumclmKfa6U/96sZkw7vMNYZvcmxzyaGmgpx2I/i3D68rb9n
QRn3Zd6jS4lWkZtlSuw6hleHUVWiCkLQ8NCuZNd27TObAJMWzVCyfJTzsFgr0BX48zS69m4hdSq6
KU9Png75cI06oT6yWuTZpEjDhNyEHBxP0AuebEdFKYl2GqGf+7a8nC8FmvjVNPLymFQclu2T/eLR
PafrdhLaSDzr9jt3QNQpL9gVE6ivCmZ5gIfkXfrCMPUffmc9p4x86vC8EzfOLAh3ypQYuQvrYL8Y
4GZuwcbHz1OIgy17B+CAvnNHjwfNU5aZELKqJoqisJA1+UaiwKLDtWD15mZyKGVVej30Y/lO6uYE
krYUto3zz1rFT99oiLz0JkpxdGjlUr/jyeft40Us6uydIl5JjUCWKE1UEqGV8vwg4tAq2vvGsoQo
LQ/9VX7lgR6/Mkmt2yoVTRGynGsfOCMow5DVRj4WMA1+Y69ICRyKzAZt+t86hsrmp1meS1PIGMa1
GYwsyriDc70K01YkXdSUlcE/cF13emiGS0UzNkHRHIwmTrn+Nk7oVoyDXoR18GDwzX6BaGi5xopF
TYrOoHWHcT0C+3X/ht7I+PmMc6nGmLo6QRau4fLjMulcedeOmlkfQVed6arRbP/f4Fc8G+45xlC3
3ACOg++SymZiKufBVsP15Qgdh7fid0MskBtGiBVNv4kDMDkAHEfYrEyHYMZbDlq9LfF36JvZU9QI
jwT59k1Fo1jhT4FHSBCnqFberrToSzBGXPjnrODg4ffzIGFv9rxowByiNuVra1/3+uAhp3y7SAcY
Lh/9LMN/sltF+cwWp+8TUVapk0hMA22AAzgjpPD8IIerYqYKsdNIXhnKVUigRhNrSlDw4sq7Pdkk
hDYbUvqTywoRWLmWxXnbR+JOIkGyqjj9GcDhPEeE0kSMfhWwHbJKhUVGOkCC6ABDR8OFtxll4fb9
FAK1mKoyg3fGZK6Koz8qonhiMPbPuqXzWHJzZL1u8khmVM6SasB0YjGL8biHO+B31tcL5Tb43o2n
Cz7NHBaQ1H0PFdtXTN1Nls2VdZ5efeEuYSu8Uzb0Xc/YjyCVxBViajmW7/TI7C7xqPyWHEAS0slF
aTBuTY9pdprt1Pg22J9I3FyNgkInqs7D6GHVah/XWoWrR8gtALQfklIeJYOkXlMyuCTV2AL9s9vq
ap/iwSz01e1CrZ0vyMevdDJD8rjwUjWVMm+XMRs5wcKrpa+8X+vGqxWVTa7/snzYJAcl3cI+29tb
+WSeQOrYTW5IyOsdzi905nLaqOMGViU8dG3Y243oe3N6oS3dNh4iz94q8Pvz9lD1YdDw+NZeVSTH
h34/dwsOhKR7qSBl5lCufo2oMrYMl3YX9c2wipVGhtiJZQNzAKxuFJ2gGNkGT0yrwcEXCJYi7mXO
7UkF4ZdM+EBzHjZDgmIXnGycH7vcY6Dz81Kti32S7uBHI56uw74w6OG4RJAS6iyE2tcwIYX/YPBc
SbuAujG3GgaZ/DXdd+Rt7FpB9cxIsqmc7hmWqifaO/+MiLH+cDZhUO8toe9YvpYdkCTgoC67ChJl
7BVwydZEr7TH2vxzFKY/ArhjEZyYGStUp7aZML3KyoSJB6lsbWbt7aMQVgtsPCcshO1t0SZuPyfr
9GwwoUki7/7oAnlcFHFlDrYhNvhItIxK0T+2WR2kv0P8/EU0JBff4rU8W4dCH2FE4c/GtZE/UbfC
gEyx1xkpf4JZK06wbOY7v8HiCeNz48st6+5xqpejwCE+/tl4ptLnQDE5OGAGo3OrvyKz8NhLpKxO
BcKzjgUuwMKyTiyYY669ueNlfHLSlr8CnChf+2p6HKsvfDhGTHGjUHHKwyx+D1ACABBGUTpKo/wp
GcWhG3rDi0NUJVuWD2Afl5i6EZJOpLHrj1LOdwpbEAVqdUTYLI8a/TOaq82pctNA3RDPDOJ8uaAf
pkvrXpiiC9ruq4ETgM7SesCZoFpYoqPrpeu+h1Tq4Z9MIeJSsRTEkbp2SJj/iH0WfKGFT6cwPDqm
t2wlbZvSfoUsibOnB380JPMCN0zYiCzw+tdgWqjnlLu132kKASumXldJIjR9r9uRElUwrDYxa0Jm
W+1IRmVdYX1ARGCm5mN1qXx5KAcTy2Xt1VC/5nc0h30ZoTZv4E6skjYNUvGvNAQTfKLWyICnT/qe
N+Zv9Z1qZrUYTqyQ7zAyF/0mO3DaEy97/zJ3ie/UkAnBcRiKQya8PkzgaayqpXTnTuZgdWT12Wtc
oywpeTk/UBiZKNkDui/P2zcGDspe17maAuuGBAz4R62YiT92fcy2mw9pTeSFe40PS+Y6DB5ibVvZ
eFv2LlB/p7z6d2dqVqKqMcehnayYTLwDkQ706LIoDu6dAbhvpeXrOpwwgs54/7ddRs3qGAcwM/NX
MKkm+qZvLsQWY5uLWhzWAm9pRuVnjY/rp79NCS+6F+Dx5k0yav+0n+iKbC7XvnMGzW0SmYiXZdUO
AcTYTeO3EoY+sEkBWzFo0G9Ik4Xcg7sb4I8wwWSd9n2eopwBeGicEliQXUQxPO9v+eKhlVfA7cmw
Hpffor/+XxLzjA7jjBiWYwL7X5AZWz4+4KhDnb6HwnX7lZ31DXNbjWOf2KLvP4kKcX8/veh03DuJ
rW6ZUcf4cudwriIboqcPi3Q53XRS9VOb1sbzeJwuI7YGnDU2KJvKN8C7X31CpKpOk+i6ZGWv4NSi
shLIGbEtSIkl00fuhZq0f+e6mcxmiw3oLPqwIq6N4HjWkqIyFx3o2PefwHfZqxbPIpc9gMtnwAoN
HvpL8EupYlk6QN4ERfGEvSBTd6NmrOUAw/P06KRvAfy9ycJQ60GT+fmm127Jlm70W+YYyV4+VhQk
k/3bZat4G841kWHE2MzgNCifXGIelYgFs78HxYsQeUYSGKhPUENHIAp+cGYIJIjVAFTG91AolaJm
NelKr8j3Djvp0TSU2mNEk3CwJ4Mm3vjlLIcJdxUutA5UE5hrnK+vi/zMNPijrEIrJXWB/ZIrDN4U
BLP3b/pkwh0VWRjhg4lXM8S7ulUtfkBis/fVPrNz2Jd3ezZkcISWq7XbuOyytll778iKj1/YmjIV
MHB2nGnDh31BZzequyG2pdVWBxDy+WB5gNbjMHw1O/2mVdFBvLATZfXjtV193HSrKKvwsHUAGaYn
rhW8oigjNxQBEH8mDeV5DFiELeZ7WDbLjcZM/62+FOgwlFHNIx2hkvFewIq8EB4Aqh8TiALdbIBH
JePhzcBcI2gYsjXgB7sHBdfBCJF+HkpRzqEjhM0w4Q8D8oRX4mDkHcSPwMuu6bDhbNrKq4HJQRBr
a7Mn50pbJFap5J0HkPonsDT6y+8WXD4rT8+IHPtouhm1hPmqoTj4RlGAZhWSclNSE/9oMFa3PqkO
k6/LTw0/VUwiyEggQ4Tmn7XSFMjMsY1TELAk+kaHbHkyU/P1PSgyS8SKtBPRXxwBQYjMzG18grjP
qJWL0In4WI0Ddxqu8VEJ47cWtMke9l4Sbodi2YHQx67nvZ3c04wa1wvtyNo/4Aa9WJrvaUaKepC7
UVRThvH/HbINVweaIrJZud4B1SuxiV+TLTZy/D/FFrPTphSXHL6jb4XHEPxxdyPS2s/wjit2bcDC
lvO/60Ilstn47CH5dTCsfilyT0WAkETRx0CLW3lTJLGWguOih+N3EISPgNccatgCoUFDU188M9+W
UMP6jGeVGmN8zPF0r67mpX46E6/Gl8drGDuWAHRDq1wrIL3LXBcPV8x8tviyn/G8EaMTWUuuEkhl
LqK4aAw0vHDZfYOsQSbQzSx+pa5/5vr2KDmh0WZaMHk0zAzRrMsjfr0srTZ3CTlHET3iDiSe//Dh
MyebsvDdc87qfMa3vAUcFmL+QhK+4cSa/i08OBGDsPgbcjQLUd3vrJYJrTXmV/Zp+bcDCsT7jUm4
j2M6ZVGkSp8jNWqSh6ZQvIlEhAzbAs8Qd7WyqZE/a7tuItCObK0Pf8ALWka9Dwm6hGzoQL2sUUcY
g0MuVN+od8GOFb6DORlo7WgWA2PIgMW/6tRu//utu0e2TiCS6MivBkUg/tI5FLz5AiTsAuAjaYrs
bNgJiJvNrKt9yEAFWitLT1tvDycvN3pXOabDAzQWTfeXaoRmGYB5nLWFR/HvTK+IMMjwGo74Rb0c
2emQE1VktzDviepMpKL1jxCGtk/ADPv1c5pip/JauGGg2Q7rgRRQmW53mdsaytY6Y3SuBmiriULj
r4P7n/M4CYgF+vjl2j+JOtJIL7xkliZQ6XHlhF3386VXPJKOVRPi4iAk4332T16M+BHj51s0qXuZ
4AXE6qDhCVFi3gjwDTWZIUruehJIYhSsrkciIE4GbVsu5QJwAmNe2t/YdmOHLAwBWpYg1bhu/5GM
funVBHxxdQlKl3ZD5Vgru81lPxrQ3dm8USslC5F8x9SxkVuJ4ZeKmjKaIVp0/dz/uw2rQP0CtHmp
oPOH5mJqBkGXetHxyMmpw5w45n7ZHblRWWK4qb79SffQuLZihMX40MLS+WaZfotmSD9/xy2sumdJ
6PGvsJu3ErP2kO8tHZ5TupdlYX0QdDyK5daEBti8iITc9HA6fpLvn3um19KRfuIPHxTmW/htIWlB
r0BSt5dZp+E02/13cgVFPhX6Rcxig9ndHkAHNKsu3Rr5gB6LqYB0+yrCrmA+3p+zES8BAd+gQjC9
vQetHgjHwn9fWKy5mKoizfy3kekFgFWRChp6eL1L4ZN9uNJ9FAZ5RhDm1KwrANWV4j3mUI9X7+ya
l86mp8fKMe+83cmCALXEW/XjKdKwQnTSxrEfypy3H/IF2ES5kxPQy2mNsjXfnFdsOuUsEOTgwRmC
voQMbOTZodcvPh059PCf6G7JoqRCiAF4EBUFY0RqkKqcIW8TvSL45LLXsl7dYXWbk0afnAU9zgjt
hUkmbLaC4BkE9KykHDEUeDWr7Rs1r6jkTUUBLQb68KoTmNjCsM9iXDBZQq3pP32Gc/cMKuRoJIbn
CWQVgfMYXbQRGMFs2U42rlSlZFIycBhmaSN/RT/0gZZ5V2fuqeC8uf0RhjSSK1spu92wiwxG1phE
Y8tX+v7w3cO1pUTPF6Ir1laeZQWZu1MuoIUu1CeU3H7EJEVnQ7VxcTICm2K/jtAfaH0YpErJ0mgp
5Vbe0P3YqiP5hp/aq64BPu1NdADrguLNY7+eYmyXd5ASBIqqKGzQR2HmKn5mOfXRWBKHxsWacYKL
hD+xU8ItlrbHAoOCAGJmFg8yWETr9Xr7LQsC/HIpLC41KbPTWbgxw5w3M6GhT9OUxTY2aXwpVOA+
MDygy/kPqnvR4j7lM2hwMVXp+Klaytx50V2Mjk0bR27QqemPX/AdrGD4XvaJaedC/P07LL/nhf/1
SUdGTcCHOkGudAoYPJ4KBFZJTcWmGa9iGtYysm34ek6Ay/tmWQiN8LrC53QMdzT1ZjxM/BOZJ7xc
4G71c29Ub4/uf8n09fA0QZA54qPi5Y7H3KD+gXyjOixAfj8Y5uRMUYTTAmz+5M6zjaLN6E56l+QP
K3AsEMa2ghnMbUYJcNlvAeOlN8dS0XnZ1iKlmGuQf/+i/6c7RoiXBeNW77/K4p697iW+axEZmYge
tOgSPSwe4NU2vDJNtfhbynyUJkL/Zk19+EPzVG4WlDMf/z8hcMe71UOb/0HBINt/cEY98wbc/IvO
WxsI0Slh1GZ3NxViWll5aBqZxQfyiW4R3ek2zWCnMwCUjqDKjWXaZ7+UUVyMRqAfz68/QSD6NCIP
A7oQeSLTBc8hbQVshPrnCx3h0WRl/roh2sUM7I7TnH8ET/tClWswVrnO9DBDrqI8niLOZv9ixw2F
K02+rpVZS5rg6ujfCGhN9ATIjFwWY9qWuGusdLmWRgYP3dfDnjPONCdu1hBG12uytfwRocgGzhG8
xuiOJvu0HAa2gopsik2KVQXyU8gz6YoaukzCVrktNi3uFdc6UKvenEwQcpE+rzvn7LSptVaRACQB
jjKblihuMJGd9ZBcA6a/fW6fGuASFZwwOlHU8YEGd0UwYJdJVYvMExj2I7w/wmAALX43M9k/8Cuc
SbwHgE+w3PVqg1/aeAiu5SnxiUP6c92ADDjJQ6KdIL/0R5E3yiHk+HiY062pm/TxMlUGVtKf6Jpk
K6tGKW7Uwwk1iaIZO3bo8ATsWX5qaeVfbu64DJtlM+FqfSxRKI3XRLJdZgwUQOCWf64qAqkXmbVF
1ArQI/JkNI9isu4DSMPntYys8pqR0Tv+6z9pGRJGfxi6c5RDeyeCHxUhDOlhRuYnAUc4C/UTfCZm
5r/Tvr+7QxcVNhL76jmWsACfdV4lN1OK/pC2GXP7yZQZqus/XnkaczlQPOm2CgW537gBoYHcWLBf
qCPbGldL4xmU8he2q/FE56ou5SNhVwAdFvZ2U1zfHyVDX7Hd0mIR9MHd5EIjIsxX/fS930gIimXv
2CwJu6O8WYBL2QAAcRe2AWSRRA67/gSVPVrjjQFsgxs/9oVGDE6j2QOCUbpWgQVK/5ntIMA8xJCY
uh6yKHVCOZjeQGWk5+l9T2yhhHRrKUzNEiMMDdtJC2rkrwHMaqz9wYVa9Rj5BLpMogMQcX5Z29+o
Efm++4dMLlib93Xq5gQJcbtrN6J+f+EJcJPkv4NORMglLav3D5f/c8vCICJXC5ixRItQK0UP+b74
uCHOWInZOiFXVGXe8DoMVi2Iz8EccpqVNklVBDK9+tNLtkE+oSDz9+TtU/kvPsJhp/UjPyUZEJea
hdoo1iNxVNRqXJHYVBmHiQiuYQR69XA/nQnT2im2MIvGSvE6uHgORyGmzrwH6R9dRAfkmIrV0Fea
TkgEEnN3kKudwzUycquH2wyJf2f7hPqZRSdmh9NCBq9C3t8eGnvxrmiM6xCz8WUPleh0k2FXuXOE
L7HDa+hscJJ3ESSuNCiKNasJaKpl5Gaa6HJYSWW+GCHE8xxK98ddxfnK6BcHi6OJtMgszdLq8BVF
H5uW2ox+BPmgGq3ne6ELQo4U1E7NKEOlycBS5qT4CBipxn2JxC8HMh941oqZJ/XEgq5oYVAdoh+P
PH+voOPp9rW302YeWbskn3qfH34vzBULK+We1HZfRm/65WHB07HM5Yx+Vztmymsj0tPsbDXWe7rP
nHAhC4l6eu9CCVej4PGxUCeQYecQHmr8ii74/QduyGqr/qcnwg8aEFtULdDUPfm5XPpEp8mfnUMq
mlUvKh32VcoQeJz4B9I1CUVcKrgwy8RLByUlL02SH6PkKbrh+qN9+BGwX8BQSgul+UhoSDdFqxxE
YnwkAjEyNPN0v4fntJ+Do9taTNrAvOQTMQlu+L4Vnl2iLw1NVBUp40SH9DzY/SpbPld6cwkCq6ZY
vEG9qNoigZrvUe/8ylZo/NS+DimS+waIrFnA0RpYfD8OupOrTMVQysqurfdXWqYQRXFgZqAHRFxe
cr5EIq6ILsppi8I6gaaDkx0TPrSNqcV7UP5T1tScFlgg597aPVOnrmkfbWdgf3nR635hBn+3koAB
RpygxgxHHM+pynZn/+6ajY00vDJkZVCC/MWx/fPi+KaFTB+aUwrZMWXSysoZLXPVT6SVvBkAmpf+
wk3NIZjsM6bJZLmxzJXUwTNiTlwRxSYYgQYQdPY1M21gQOLjXSvsnOePwzltYcTUu2ZqIBFNb16p
A4TXG6P9ZfdgRw3pLfo8LiR1Ji1PUvbxquhwZwAcQQuLDGSUI3RqekZgtsmjwxlN3temTJ4ALJ+X
frv1kQZJnF51N+29zSbVwpE84J7osyu/g6Kw+R5MroNLLQcSdFZ1LKouCw+qYw0Any3Kzcly0htr
rzJnF7OhQEm3rRpZLLdEkr5Dexd7Io9DEs8TEt8RrYgceW6o8OWcuCqdKw/8+kDyO/lrYbUmFApg
sd8k+QRw4tolvxBR5uuDTm4pisxfTBeIEAwR4/dZJmTmCd/IV32WBVWq+3dsMnOTObQ8bj/l0l0g
5WXvAOCBS9k70sHY4SdOJEVuqJVsz52Y78K05owOXsLUvMbaJtY7mJ2ZKg2RE/VcVSa1WDz3ikiI
U6giUBOYJNnNnNhDtx1TOd1Nr3hfUyZqsETtlCZtqF3rP4Vx4shApEtBIx9feDSzgVFoViRT6Cvr
skWj1ax+cJA63VpryWNaGTsmmFBCWo06ZLseQCIluf9EkEJmHtN06bUcRXKqp0agwc6JBoJib2lz
D3rBf/pOjeoxarH7WKNNECf++FMM4dOqo1/HsfA8w0Y/bAoFEZXCAr85dcb8qqY5hHZMa12fzQGE
wLS1PJ/MTOdSOG+MwhmbBLQDjftL5zSPFOLMgFN5hYoszr4O3G4z+rRFL+GufeHoyi9Xt8fvdr/i
gMvxgzCDyFkUeE2LKWtf0xVWpa1cX2heZXxjdPg06a17Rh0VJqccBz75B+m2VmmUoxaCoFW3Rcad
0v63Uk85SThA9zlkjal0ygAaL5IKJE46EwtbPUYN0GLPn4n3VYgXI34NlTOhlIiELuN9mbFMQo9d
Pn8SrpdYqinr7GA7KOx0i3lb9Ef9fXakrLGSvaKFyGM0NQkcub4X4/yHQVPyAGs3SQvGslCUWN6J
Ko8M4cs8NWbryZkuEfAqAdEddRlYwp7VPndW3v/Sq1mdNBTtgdo7RzXO8asYp/TaVJyu3Xk+a44Y
/FrPw8hozthRhc3bMPRhpV+QgeU1Iuspi7YvW5Q6TtJkMu+gYCDjvJ5XM+chhIrWADtRlBZlAY2S
vDthyi9HU5502GpHWxW0RJXIiO8kN5cspGAjAAN+9AXMI0HN2lssBq1vA71pT7aFef34kQ17UDuh
k1dILh5mzAAZiHpNQTxaGlPR6TEobwTO1jTI7uSl3FhtNmcOJv7wvKtsywPhE1zFa4/cTX8y9C+j
oV+OchMcjFdV7Yre+ujXf9EhAZCFvFkkVl8NetHH3Q0yW7kFKfuqpmqf3gllKXLq0NxJD1tpv5eW
5H2uIIMaJ62hiyQ3h1oCcRErRbgjx5+Svk39H1MfkQp8iHSYgjh9ma5UxoL+W0mlx0CxU01nRFYA
QjQQcNQ7WXzA5SmadyFBXgEyv6SZhKh3yhvqTTQIOOOOVVI99kC+kz0A75ro0ORYJA3tbiJ56+Un
I38NOROqi9TlU6EfiBOFvlWUQPQDeOjUSmoqKiAHNoxuefxT31webUBINTlpYxtTxQaBkX3ue2yV
R/g8wPpxHwddsPUvXWL6qPs8qU9CmyQr8Y5/PoSLew1dWZkUf0lygBiyXiYZtnVz9Nz80axzWe7m
zRaDlxxDo2rrH9qr0ewKEg+6pyg/H+QFJltrUtTeSdx+AFnRGLV6tbkCVUC7ujj1nsf3Li2LMp7g
pJomq8wZRaxYavhsDGWbAtpGk+kssZ6mfnXs0emxDaRA6z9hvpHsLyKMmJ3QHn7Sy3mqNcllAAnP
kpfrWIW8Gm72Y2KH8lPxYpTfF2JndEBh1J43/v83ztNHSpjZvFmoRP7E0pmlOaMA1xU1LBHqv15G
YxVz8gY9qOklvxWnROG6WGk+4hsVs1bju8GD10t211mxNnjptUhL4lfnp+blALsIZlQG9K60Zt9b
SAgTQ6qMDSl3dg4HJsRt+AqOXvB2j2P1XQYiLOAl53D/wL62rx0IDblItT8x7dZW30pqKJynIMli
F49OqiJTkqKDIJxydJgt9Jg2/KGZAaQBn8UKarVWPymtuA4xyDDr+WF2W9EAN4g/Bq8sVGl/cv+l
dIiW4B+AICHofEDjPI52EfPNMGhJJ2cNjQi36VhurVhg25GIE37qKOlS+KsADMqJ8reuYfIS2TXZ
oGXwgLsxtS7Tyg2hpajVoJuOVXlvBVIz+gl0BYjOl+AmVP0tGI+Pp86EK+H7G/wq4FGAWbrwcpxr
ambPDvcnbhLcITUQErLE6gCZwrNdz+EabgW8N1EFxZroBi/5maqHuxL+lSKk9DFldkLRJTPhR055
0FNNoN+NSKkcW3JYh88UpMrC8qOkBl4DnRojz9jbWFGHcZV6G9akwqZYAdoX9bF/kwxotteJfUwJ
/npilw/UiqAjq41TW+ydj0OMZL1Tu39HymzJIhuCq2/tURpfp6vAVGL2q0ZBP9begdM19aygk1lc
qLM7Rux/L87Qua8NZ/XHZk9eLJGCJ09zFCcby96EAUf1r5vROb24eyTkceIPXlpChL4CL3CWcGN5
vU5r652/NXgb1cM1XacclZpPp9kRuRJSy1ygIziJww102DxavH/DKxrwOLA3gOQBUcEKBaZ0rr6w
EDZsBy4OLJ7aKfZKW8leTGoZpwsSi55nyW+qXPFIYw2KmbFVmAUGcXKHilt+q29yvYorXNh3Adom
mfyI3naxEEQXw1WvHtEdGGndQxquzWwFewcwIVeL34JTZsJk/OsqKeMcuYPeFDBSLCDJW5GFNpU7
m9dVh775IequYXInbfXkYkRlIoztPJ7gzYlsLAMT58pU3Rf1dVLRPd8Rh41/8ChvLt2FALcvZGCU
Qu3DNVxub9qOWbmf7dEY6U+AJTg/yjfhIJTu0uKPuwKqEAU9VKLWXl8YCf4HZL9UqeEu/9/dYdH2
8S/Qn55pv4R2BcE//3Z3CVwjrG+4pbWmJ4YLWmB8mwCwLTy9CHUC7I0bBPrIxFj40/+tuXna+x/H
iNg3u7tvcGKvSsHa9gQV99ym8NP3yz5nJoDeevZ1+JntUnkVLu7Pl/AMQ+qdNGjSfO9zI6bjjLaB
xKsI+K5lLbY38ruKgZZjTVVa/aaovPw/+a5Juj/n+NZLctwj12NcDPD9Un2pMXzw5Trq8RKSKXZc
vAmz3Rylgz7ud+V8lbbwW+QCc7p5hnWLQySdtGsLyU/iaZYc5RCOjs0Vk6ccQxUELXwrg+VmwJyK
gFjtSRIb1TXRQxBgfkhV/5Y6QoF+7WTbi+0ywhMTT2B/Bdz2TEILkowNwpVYl7aFTj4ORbvKSEGO
0E0rl+7QbgpYt4RiJT3e2JaqThQnZP5z29WM9K7TSZjpCTWvvT2sDVE0SQv3g/jywRq1t3juGbC4
RCmFmCf30FUeL/EffD9vzbu/r4fo1oMjU+HDssAcnTCC4CXYs09oRnfIkqYMiHz++EfiXqdyEWCJ
7QWVQP1ZaFhcNe4E3JJH81xSRhN0yI+GQf1N8psCbjO4m57Fe16WgSwhNpoAi/6eJKZDQrbFwWp+
uMA6kht/ffh4mtdB+W34NpzOmitbnW/TJsFsnVHreOjwb5FK06cMLuqJZ7WX4CIRMEJy7KpPCtOe
2YxYynuPztVf6q6U+trNoM2XEBMbrge8H27e/WMqsoX6MDcyZJJYcBhCDS6otfJ/VsuJp8dXLmMg
Uq4w27aWa3nLauRE4bzD57/eA9zsLDpe/UNvji/jWEELosloK0thSDYm+y+PD0TEDa5bIJgEe94t
uFtU5bTJAP8PorucR3teFAN5fnSYlPT6AeaYEfJeM6makGdgRkN7URyOuU+Ieu7tJCRpuo0hhORF
QQPP5GRklb48bnGr4Oq3pLwMfQFXaZuKqXFfX2aVl2A66MfUqXGedNFuwbrm0GYrdJX0m5LIdgDA
63/8qGJSH+/HMRX30lMZhvxj+Nza42Zh2li0VYKayi1tmFcHNi+A9WDsYOyQt4XgJp0jBTuWrJFW
alOKIw6F6s4FxciE5cOYiCaUGv3qiSg/mHQ1dt41xybZiKaSHHhJFy7Jm4V75lBgDBevqxo9H4e8
H88GtjXqCb0z3qxgshMJV+YYva8tBd75/olKa/b/XTeFuQ5kkTsHhYY3LulsFJC9zwMFgXCARTSb
xfdWR1XqvTLA3imfYMKOkklF7jTAAkyyKGj9VCzaobpt6sTXnuGGunsiFEhr3r7a4HTmnF6paVHD
ZC8vem8OBjyPWizwCuGjcjwJ7X03s2w4mnJ/+xbJQtqtc9niRxrfNH2OLBthf1yjYUPU82nA6Dnq
PBO7tIsciZw9/2geTgk01UTT0FX71BrA8oYAL48+/NQGJjBqbhctW7XSGQ4NziwaHHF5B+KqmfW4
iFEoS03JLIj+OGuWcmKlP/zerf61kFdiJsZVZ3YfEMLPTmltHVgq9gyTqWVXRL1/UqFSQkKsSZGz
L51akpMytXJBZ2TaslIMGhQJVqHlX6SrrlL4/uP++1tPFteSQlX/tMlSMNWz75vNTxdkrCOVHC2j
iWjpoojosnTVy1Aoh58ioipOahxsVJG8aFHd2HOUYX4H2SgR2W64sRoIIoU8QfK0eY2fbo6LGkB2
IzKYSEBLUT3q7MQoxpOrinTBCb3n0uZ6IyjL8M2p+gqUM7IfWyqD636gnli6VOex9MEzkPaG3WNt
tJgjmAmgSRUC++a5YX2BCPCIHEIRPrV7hJ91hra+KyciBgnLEs1ATgZwYG8SvuGMHLE9Q4jsKGeZ
StksvnVoEFfVZPVYADnBOyotqty0dt0SCn7bFHOQBgeh0nKRCV2KTYVWWnQLwB92oIN0LLel5pv+
W2K30L8N32IwfCEwHcf1YfRVNyzDVaxPWuO7t296opCbGoMH02GZOMue4cgOqer76j3b28tJxB6I
qEZ1XGzuj3PcGC6JmSnm46Q3XmVx7oHFafYEzRkwkXXCTl9uP8zjyeog9IxJWuQWPzeplXL6Yuu3
ypaNjlZ1FXfOJdEzTtMmjLs+KwMpzg0WHJFrXn/2MO6XgRZszIO0K5Oq2agydVzrosFamp/67m+a
lTkC+M4QPwFF067n2UOx4VWLlamkwOmVmYtWhvbI5iGUgrXk/24rMkG/DzzicJFIk7Mfoe5jN4ka
lpc6UrhqFWtEXXNL4owKsXCPUxXHdTSKAB3/SP95dBhPjplu2HAuaCVV0B0h5JDdLLDloUmaAVNQ
iiEAMqjeo7uKlFVAoRopcCw/iY3H/3ueGwZ8mlgw7u8a79E/zCw6JKeFTmL3TitTOtNb1i7fRCZb
cbbVTW50mSSTsFaLj2VceM3w82wCMRxULs39iESQD0NN/kIqo3HbPFrs1CyJ0dgG4koqkHEEGbaM
6kuIt/8SeDzTdz0vPPcg0q1QauRCvk5Aq7SCjblgXbCn2z6x/mHEW/HEYffmTJ4T0MY7YMl2WMG2
BVIvE/D0qzPW5W4+uSFyEF3hPRzNU7OXcHbiaj95a9lmb1xZdfv4RJkm/GW6+5idB9J1vp9gl8UW
5t4kYJXH9Vj+diRs2XgEhRIpyGEdGnCisNSE1I8VBYyyQt38ASKgcjMSsdhUqAizysBd5Mn1ra/o
upe1i0yV1NM5NuBehdYqAJX8rq629XqDnQmhFjZCiOjbZEMJzsV4bYpvg92BUfrVfFgV7PdNHail
9hUYC4QTGXfGvFJl0sV+QCq3f5oZ+MCk+grRWLcG0PXGE7EM5zFocSVQuxenn30zsoambH7adxWY
7eweAJ1aJmeSk2PAeA7HlvAZFdnzDLUaLhfC29yciqhsR4nSF/ymee0/Hs1omw5+Cp0Ca0O0/neW
CdEROE/wQtElLEOBgFDXAhTy5aaloGcW1QMsIT0FWh+rVczkYTg/mhkCkDoJdmfRJLL2kS4OiHEq
r1c+SW6X42cn2FJ6x8kSGhOm4VA0Ls+arx7plsEokU0kS6wIlAakxenYLMuBwmHWTuHNyhuT2fA2
jd7HM9VUotvQsGX1SheRWYfgjWGtcmWQ5WthlpXG77td2Sz7nPjZTQUq3f7umji7ypUki5d3QZ2k
bKOneZbt8KJoWgFuJC1ZuTlzvLuzUdqJmM/0HjdWC5vH+XCnAKKCqtkZ6ImlTSyXtunqYtN0Zwf8
UFxvycQTn/E86E/CVDj436i1C7u5GgEuOiViGngXgq+KcrpuKOLwZ50H+cAOAxlLCOci69gSEAFn
tbsGYvNGO+WT9sZflid1up9ZiUBWZmL5CtiDCf8/V9QCAh7Ah0bEBsjaw/QkSSb37JjjDAYTlH+N
LqfGUS3y7FOWfNJtFYwz0tWVo6BdwyxoG8blp3VcdXJbuF22XcOe0QnNcfh6suHsGv7UGGTN+yWT
vq9iQUGtmqLwXIbrXUJjk8v52XXB5g3C9Kb5UJTALob/jxqh/3/Q1AQmBwj1waLi681hnAHYRUwJ
05a32QLcGm0+bqKmA3GQf5tZWIq9Cbqmq2F9u8pqfqi2ZoNjmYlUzYabLjW4oX4idw0Bwo2/JATe
93oGsPnR83bLTx+khjB3pt+5OVIOnfzYC8zMiUHRDjWpiFfhN59kXbyotx8WpNWYvSLxT1ftrVol
n3iDSTgTQBtW9GkDfVgbCx7Kdw+8Jx6V/3MzczaXqyVVd4ffoM+ZmvI4Ztolh+cWuQEU4RN+ZIPF
mDL/JW3DFGedRM2O69lMXTYsX2q8EuEdmuV4jbVxzLahFfEnl/OiLKsQ/v8dDKljtT9RMo/QUQQF
r58jeUNP+07l28hWjA1ti946aTJHMtzDjOxYDR4f9vg3onCYI6BoRxmRXdVIAtWY81rBYuEaYwtQ
VpZ4/q1pfO/SG7rhtHSYLWS2du3naPRJ/QBIITZNLED+KudjxnMsaJS4keI82Ce8dqAVpHAKDDED
yvfLHYIuOb/luz5kl6xVAmh5AnK1VclO8ZMHXUIbqb9WCEABt3HsFH42q7eoW0fozsdkNSkANTch
p92oxsTcnrHBV3CKTjN1fXl87vLLEZYtioo8uYO7Vwl9lFnpKtg26NWlvfiu3uqyBnjQHSkA+0yn
Kdc1l2NyHBP/TGHvyhYepGGv4zbWnlixVl84YvC8cXOr1nbD9seoIuhHorE7yEjmhCrvt//En8jl
ZjqxTwDewOEYMZAful9CcWYpKyH9QnwWWZv8hx2mFihA6vRzyUg5YbdydyKTgYrPB1mYjGMBALhx
9EKYKebM3mzkqf1pz9YQKWfw+87fQeDogqVWMANPxoz9adBuCP3wRsq20XBJg/TgdXPyj525YZBd
pvjesI+gqjmSuYNVnNje/RIfDPQxH2emZSKTPiCzYYsDkFkMV/YKRYG8/VfTjTd03KdNZf9XyTno
JsNImcbk8w3EvezyYu7zLgzMFQi3QhocrcuYsZJUbhLdqlBTasA4ldGAY8vOzhkUkfGR2IVTaAll
cvb70lzzrS2VhOFqZ79dxZQXJGHUG2MTlkKMM7dkEBX5mIGwjjT2fMSGmbucwurYbiPy3cTrXY+Y
0urdjLJDhS9bEJ3mcvFJH47tNX5iUiRUAmhuVvt4dv7sdmm0VBDJY92U1vjek0T0tb1mZt+hovCt
U0IIJJgUq8cplAm7n18TczNuJ37M24bTUFqgEGv4uXp4CvsOfY+MOf/k82oFvuq/KWbvbMQUYOr7
p84PW5SCK/1BNvz3mCsp3OVW/0D36OIchVLZba497VE4bOEKnRT5yCaAarsOE+F3sJwHSctZJ8KK
WlRsHftuCNFzu2cutgn3wGDfubpWpnmY6GMKlA2A2sVX7G7QulVz76scIJ4OUyVFzU5woCLWi229
NYAb5LJkKyhM1aWy0wClyX1PV2pspL7J+NNLUqRdqxSuhNEaXvE2k1qsSMsgtdwJ1hkTrolmi9s+
TQCF0C4XCCUpHyxdp+QOr8aODZcN3ioNtYRfigowRd1ZK0LJcTLBoxvTweqriO8p+6Na5UOIRgrn
/vssZRPu2o4ZDMCe9SPWscEELzjhDG3di1AG+mggZXhiYgYTQPeBdvrRfcIsIiCQliYJ+nZ9h5Wc
EUuy5WyaYwOxUjoIeFdU9gQFCSoDpvBej1hW+dWvuPEvKTtRlP/ZvlmqgTgSJS3kJpFTw7+clYNE
AyaWnAgEUgXQQs1ctpx0cnhPDiKXlC+mSpphQ3zQae6OG86AtJbVPJyxYw4jKArp+zUyMRWmkOwB
VJhN1PA0TggD1/IUdlEjdJreMOwA8mGPKBqD1CGoM2TspcCTHWW2N1PtKiv/lFi+5irgtcMSBfL/
x02Jgagbt2Wrfkyli6e3qGJo45Le41r1P3oU9USKO3opnQ7VicV+q/L+WGsx3/jYGG0T5w8hmQO1
BI+d48MaocNsbgYGW2F9f/KUkx/YcTpCW0ktfT8RUwuSdrN315brJCWfZ3C8VO7zuUtev63yY0mR
RSG+ea4TMZZ6tn1XNlmS9kLB5hftiH8tevo6+VlC8DHEmdhCr1vMZTwpCGkkwcDi43F9nzCg3ohr
ifLxa+a0fPYf15W0M5UsGcolRvH4KMRn+ZzJtoLPCb0oIcgVSte4+22XAvsSq2imI7It+rKcFOav
ArDGJGCCi609pIlSIzmOER7kYb8N0EuBrfMoqk9Pm76ccrNGzNCjkpCMPruvzJO56qCpVbnV4fvy
QTFOcbmRfTBzeMATrTaByHSQE3i9v3M9oZ/We0ZFElT1z61c32lyjgDN+ePC5pispCrV/XKe1puv
pvERuhMLQa2ENDN3CqoYawj5ci2VkCAEoFFmRZmTdVv9FfSp+3ednDP7R1Xpgu76xmy32Wc1FgKx
3XK80lf9aOFXcSnACqunY95A4LaPVnUhT/NmqJFtslTumDYmPQcjVCZi9Tah/TCjhNRwm7thWd3y
6GKA59TyG6aIqD7K2F3ZKHV/MqlGN01QqTRgDyPrLD6LyAX+aacRI+lexV11WseKTARynbxQBoDu
91/w81BxqduOiYnIG3SJ7G0nY45oJzXDvaACQaF4u7c30jUHhoL+rco2JUbai/x25UQR+H6NWoiO
9uXNP/PoxFs+A3PN6WAjHA8t26kdERHBnTRcwREiQcmP88UH3mfQPeemEEcWVV+oONla43I2ss1x
Ha5bMRu1MCXC2Uwe1Y5iSn887V/IC63Lehe4Ec25jW0ywRMqnc6juRJrACkvEHU4jHCr0V8qtDyU
40EFYFwxRkyDnW9uCAUeoJJ2/oDXz2Q5rXSSxMn7QMUI9i58qKPHZvyDSSXKZyG4E/q0Mu5jMQb9
szFb7cjZmOIOat3AQ2rNpENJPXag+y2h3jx1HCRRyT8miANxZj87C5+Fq226j0cSsTTt5Pi0VpPM
hwW0TJUFIdl95N3B7ZjHOW/Zb6hWjTReYlIqqL608x2Ja7bDEgtgJ3sWmQrRLIM8CSd+2j84K6tU
RAiae+5lC+uvl0xuJ2Kr2UHpcRopONWstFkdC77+v6Zqk2l7D4/rmBu7UPRbLsTfl53fiYIHadjk
5VncLQ9qbhsYV5r3MaFMyd1/ha3qHVtzjYqG304vFQTgSfkyRVNqeB5Von+qx1C0oX68Z7m6ZB8H
hAQboinNtPNCL91HEddlLAihMbGdZuAN0ffzrb4T0c6jgstqLU58xPTJ2xZbk6axVAgZMjUS0FwT
/mR55GPCMWmCypYihRE7TSbOYzBXfi5kQ/4JaGB2dtqx/gwWzPZecAA9kHOLqLtTCS7HifbA/NJY
/ioMHdJ6q4svXnsYOeaPV4hnozS6b04r7clgip+OONE+u205UdEObXCjtgPVxSIBlmCCUuu1dCIy
zsOtVI7892i497QwimW8DTAoVKHwFWUAGjyXihbwklz1COzNtMcvxkKOiglYF2YgX0P5qoO68lSG
kb+6KenxmPbnTyD4IKBvHVpfeZ0m2VEV8mswo/r//eHcq6BFvMgFEiSI/WSNMLtWuqC7MCJF6Co3
GRcafSOMyL3o3xkVx5qs7s1j00vAE8pMQlzZraHj6Sv6dQrLJYqWLOWuJHOMQVr67gO74vfA1uhV
EovrqWyPRDu4uE0LkSBePQv2cspYUJdsq3NL2hLMva1w7nTcoAwuo4ipDRaqov7O00NSXNpJDWFV
Haga4lWmhl5mS8WXpGsD7go52/6o6fRwg2Vwe+cgx3xDd+ZbwFsXBN1zDmdgVeVyi9ovQzEsMow3
mG6T69UZOWMXdgFh32nHyCPvXTXjziqEbbtMGUKlssgy8ZUXDW6ORIJNZyp0gjPKsArT42Q3wbIz
jMYh6SqikyS940WiFzcOMtFbLn3vVhggc+/g/iATco2UU84DkdDl4BLPAotXHJa31GcqybWm3X4p
2FbCruGESpGitpGEcvzOAf8DBLuu6XGIld6kr/N0rdTiVUyrB8Oex1w0zUsWtBY8YxRksji+3jiG
4NLzyhPeD1PBruqMXjjevmkxVVDT7UEKyMXnRwV+thnhme0cJiyw81lk7S7OV/dPlFHXLomZztsf
Ba9yHFDLYwvaDMKcwwhpPT23tzCuArfg0p7pqttbL/pgc1xu38L48q4+ZEEiQDN404Y2ure23iKS
ZalHBFZvvF+EhINzmCvlAXsa+AHquzJmZoWZxYn4Z5p9hP+eXytyIWMBTdKOi9S1lXxYGjNcohMj
j+G4xU6obRWf5uosdl4Q335NOhtgPToaXgvtQi00MweUckBv3DjApFRlOHgX4QQwxCJlEankFJwo
QcJOKjLjdKkc44ASjzxcDimlFe+muXIPUaJ+PZts/7NqC0QO64O/FNA0gUD+62i/YE5iRE+XMX0x
xNKqWV3hpIUKWNjSZaqVVo9+GssSKvHGaLmm8B07+Fp65g4PQFisjvXe0jAJ0GuSZUePOWBtnP+U
sZdXcdoN6nrTRpVlFWya2fK8DBOzIzzVoxK+qyJnyH8WOid8LhwM3AWvlhz/O2ZbQ8ICLAqFP3Db
+iHOk9tLL+dbkLaOCp+3gBZIIDqqR9yZ844nxMAixb1JzgfmrfzQhHRVMSreYEwVkjeP64IL/nhk
M4yXrqA5ezden3/w19ilgNDsZOxaFmlFsv0klwXFURoDu2oerKsp52yNwpB/XSGIfJTj7BeWv0R9
Rrz2DVDcVQp/C9WF5uCwUhdAeRVX6PY6GdybSTysualDkFigh6T2plJBHsKSopjLBOiJuUl6UFm/
32oBK/kLkTkG+SwD9CnEkx02cniIEfZNbkEorKweyFzB0lgOCWkupoZkbZOhcEM3Cu+OUTLLLj/3
I5xvtN5wcB1+MPIzXfV/BoD32wLpYxiSgFtzbrP17N29O5MxZbmVWsCkWUxw4EkJlMWwtdhaZ33N
BfppI2vzzqvoh2f2y4QwyRAASsybHDxXFZMT9y1AVOfyMGg+6xyzyKDr1m8CDK8a7q8oMnhWDoAh
I4oogVElCTvW2+fVN/AY3PMQuw2sWdnXC1wP1ZanSIw6jBgoazJzcc7BqWV2q2VMy7YjK2wVIelj
cNamrHllwcCfbIY4SQ7CkkuhA7Z7Et+HSOiTycJOEnghu0sokVJxRnNAH6KhXZlQymExBxaHZWAq
IGcXxdaF10WDrKOlpmcLd2oh/pPssvGEMx8FwnQj10UL5eKfZyXipdggm3AoNuPXpOM34KJdoVn8
ci//f3J5OUjy25HwnwLB+rKVP87//EHR0t8QtYnxVhK3L0uq0D1A4ZIKpRxTsjOSOKpbVjJhl9eZ
bM3bNz1ONMA0buGmSHIH0xA6VXMoQT9/fh2sCzxP+PVwnwKPRDnQUgwELdqTl2RIcWTfK2AXl400
qUVQapAVatWNvltU74DB7USiyoaIa55UvmCOoee13tWarcUU2VmiSQxOaiQixNnEOMTpsR5RfQXK
rpT4ikpCatOUz+285Dde0qqxu/99GpdNybv9El8IfMPlZDhHuU85zY/23BvLRZ97o6QygYnebxlA
es3zI+39mcgvtJjPAHU6PLRhPPh9Jn5Qx+H2bkazS22IXRPFa4lTEw1j0xrwWC+HQtAav8umn9LZ
BDFXuhgf+Ptl+ydC3VkfoV3D14JpWs3l4QiNA0RMtgHKvmTNISke4U1+Frqhj5ymxFaUUp+OfczZ
wuFvll6U6DCKw/DytgrLEyxIIALVG9tCnB10hX77nkC68EUNK6vL2+FSLdbs2fcxVN8Sp58qM+eM
fMvta8LBsvBaNcOcYrNiFV0bMfEoFMRCZb6M63s3/rf8dYS5hYaOpzIY2Is/R98Z4akRSdXYOzvi
a9cE2h3nQdFNXnPFlKk6u1NPfqus7hAUOzWqXI1JXL2sIH/GCEU3HmqRRNf0iAovxRiJAxDxAELH
M9vGH1Kq7WiiQX2Rp5O9q883A79mWcEYf/+EqbY/8gRHrJ7Ry7gJIoUJjIDHyQFI2KwPjZCz/TH0
1Dheo33xQT7XlkQbnMBVy7C/sXjCGMJzg8sDlrBtRUStMjefC9hENnyUFbfO85uIdZOKfAYpvng6
JKi/R6aEFV0vZUBb9Zh8uvJZZ5UU4f32PWoomwNqYTXKS1D7NISPavYLs4MJTo6xX0Jfqmp+5Q/n
bmEsfR504Sfh7ozg0jYvGG3y5emOjYm+QtfpsiEs2L9fQJqFaUNTn0QTmh2Pv1y3oeGtL3LsdCDQ
0J240OMP7I1TiIU14zq8isnUb5Nr1YGRttCHddPxel+iuIObL4fw+abYw3b3sWXAykzRXzYtdIqZ
2J4MQPC5aoO1OyqO5TuaeV3KMPuPlnA+OVGaGE51EySDs8CttnCk2QUwBgiG/Wkxy4E9VjsKnD6D
jDxtZY1vOAfGWowB1RqVcOjcG7Iq3rNzD1cExtflkEDpXRisbHvXu6Sn8s1bc607AJRPIO0zaSJA
2aJpvutB0rTRcaN2StCqXm+tVfOcRhKIyUvKija23Vb0esJ+ijSqyPO988m+Xj/7X2CiT/ERqfnn
AzZthL8kv0MQSUvzIwldSPv9vvznNP0LIHcI22DrZ9LahzeWbadyfvdr8LCyx/Sw7f3tsHdD88Qj
fEm5yu/YllIx7ppOm/j8V9waKTnXOXxXx8DHlwRgXe1W1wkG00Om0FewpE4evE6CA8u4As02b3mh
OHYUzxH/RtfVXj62wexAePwVoFdxdVajp5VUXUm8gdmNnhWcifk/iJgem4qnFCNrS/QRIcWhgMKT
A8zm9PjJTvWbBEAHM+ojKTF9kkv7+/cPEiQ7oUExQQnfH8xC+0QVxSrlMuCPh2qE69TwfzmaCUYd
Bhh5eEE53Ipe8wqYnaJzPTWr3wTssAa65MX3B4xX8if1LDcNe7NDpOqFFAg2iRdFF9q8dB1pepV2
UK9MJJvMDNRCMe7nJ86RQ0hsleSVbhtLBGnDHDKLHRpUf1T6h7PRIkFKuAHkQDmfjWOw16a1d5iK
j4UWyb1GLBPYuKG98vqLb4qzXUl5Qpy/Q47ofYuPYzl/Run15CsHN0bqXVAdFHHzvUZxEk42rLCB
+Rk6P8k2d7zs8siq+QJk0w0KAoivwMe5NsX81GzEH+MMHS0cCO9aSx4+rbaa9ceTn9egjKyxWVpM
BSrYq+H7htKCmwct9UjOEx5AZJMZ5h4Ejp/XK5Bi593gP4XSB/hV+UPrpiqkSy3JnkCeX3Ws4pOG
eczNjhyUKOIZSyrbTsMh20NsEI4pfi1YZdkAtMzr+tG8BGNqA679dgUqBrEhGHd5LfUyc2Xz9Q+D
sRBrcMC7x3ntfz/henhlYM6fGwiD8FUCNdqdB6ODwVWWbwaNv4CHE64gvrf4r8s5crmkVCr1heRU
jNuMct+jCwf7fR4VubLvRwxs99GYzkWP/Y95fBwfAb0xGYm2qhrUdr+wWCxHUEVuLS6VOb7TkFo7
Rdva5XAxcymmofBHSIezYMIE2i5qHQqv1PeqVTbvyrzwPhSHuaF1CZBcRRhQVU8aQnMnclTm3nvE
U6yQEcz1gwFFfQpp4EQq8d9ESQMSipiRID1OQScqSaHQo2CyCQOmcAW0/1RmbkAj0VkEb1X4S883
sCziBROQyH9ME6Ynbs+dZu7oRwjriPJgoAp753dfMXyV6wSc2B7CvYKhkjf7vmm4t6EH0sjcdruu
IIdNGZ9eF/nN9hvmYjF7gpkIegEbXYeBPqRYCMpxxX0ugDm5vhSF/lVNjxRtcG+kTjPED0kDuxBW
lS4Qlt5v4zFMPSpMy0Bk4zfaeTvbbwyoKQeVWxVh12GNp+K1yMw9Drb8e9LuywV65sgSF+2y6gto
91NdZXxwjen7cHqMQ3YNjdomjK+3i211JBCdtENBopf2naCA5Vhtye/y54xW17N0TNZlhydnLXrV
IMiOR2MM0jWwPvfu8FMJUvq1ZnY7IAg9G8pGhtbWQPkkEmx/nd/LBHkug1bUYib7moxKQ/NQuL7U
I2yR0s50Hzp9MworAZYki2DNvlaMYlCK7UFia3rw0gcQ0Sldg3LGxnxF6PXeib1octCC3r+GgZis
AVWZvvJxmGch+B0oVp/KvTVA35DxzvPyNrKh3WGicBIm64AoQlhNAnL7pyq0lqLBnySw+5boEBs+
BoKuT2AYe2g6bsJOw39BAoNQ0WtkrQsSuiWa6cvkvgpX86aU4yR1jpat5EWB5GJ5NlpF2zA3qiFL
TTTeWt6pK9vomI/fcHVg7tdyS9oYqpeJYfMremTPebf0o9Gg9DN3M30zHAaX0aKm5WSoch2Y7TwC
EHgXeId1w3QeRZk6Wg3mJGC5j7WTB9R6bUNJM8EsFfylEPLK3bChYrzjoKRWPyoxtSG8lbQeuz42
ryqgz5IgyTj4rMuFWAb5iO4FP5iap7LbwHeV0qb2HnMS0iAxHfNqiUIjMkh+mBuj31MuyOAk8xRN
/wv4InNCitX0ExPkLYbC6yNb88tlElh1bN/X3FH3q4L24CyIBdlA/Ph/rxPiAnqunnxiFvAz58Ph
S4xucS9uBRBJyJCApbnlongIYpcgE9YgtJzAr+jAjPVx+lPwOOAWC45+tYJ/0GU7uCAsBsYwXJV3
+VroXevXKHnx2jBKIGrgqXzlo0Dw6L6fQFsD6Z9pfQgivp51aby5bxQLWMJxO2r1ef2XpMRflTCX
hB1AUWBCg1oSPJ7Jo0bZxJwMEeuKEda46egPEDIkZfYsnx6s/I+H/W4QqcXqsgo2XeqGFgIzzvG0
J0JhE2rxZaodNA/TRTJRBb0xJgPsizkqTLxHq1PTvJirtZW0qs3JPwD6A1Q50uN679QXkdh5qrFA
IAIhBRAjjdDZ2bsJRx8wHS29GfpvJEOb4BR0C6XuWM9C+GHSZQ8/kCKl1Lm7aACBh/SMpaOaABPp
w6noTmo4lT3mwo7dZp99siUCPewjVIiumuZ028DrGAPhl66Qnev9g6t2RYSCQJDSTb5KWtC2b3A3
UciXHcF2GDOP/CtHy1BTGeg/0mxlfqe8hHK6jmXfVGX8NWevNLynS06YLWUsJHg6uArgV44j1IRo
fem0ILoyLfjFPkmbARZyF2tEAy89gl5H1o3snrY0iNLHtV+LbWT7K+f46KVqEe13Qsg7VZp6KwSz
lQKr8LvFo5hTu6sNSxNVZnqq8a7P9dwubRdmKRLjAH4f5hhQ6KXFBgGXPfGNg7/K06v6sCLmKLHh
RbXJTqyaSRDe18lbXqa77zmO2WeFO8iVbdXxDcB/RWNfAI5tlaP7TicDSC7n9QZaiKdCJP6xmQid
ma5x9hOAczGdWm1FKoUhxT+Rf8pVZneKCFi044ffCfUGHm/1gUl6jtpJqHrs1QgeshZUtkGG+XDQ
uQslIi+zWqxi553LTRdZSie8/af+r97TTNzknUUG7HIR/R1W70duphaI7wosoaTVg0G52JysULzp
QxI+vnqUfJvE+4w+6vMVPNkp5kjYRg2zM4TxmnfKDve7/UWFz7XMU0GN1Y8wwVRtHWQWXYfBBQpP
0mfuRsTH2Z3sj1aowpXpVVda5PFxiUavelVa5lB/+7duE3P3Qk9QCh/xKLITsJ0rkYFEFcy5AFHs
uuLyYjqKS5icbS0Q7TFM+cZ2KXJaZ/ByB7hn/2qjdE0oDanrSRLdj6KYB9m+yvF8uGN7HkJkcQ4k
iXFRFk8ck/ayix85TeouqTSuKsrtL6P/3lwhbEom65RXfGq1TKGpccw2eC3ceNcS2g07jAtRrdxi
w8Nl9KbjEeKa6vGCVdcdo+xLWnbzQf7DI8RRHP/6d9tWFgJ9BxVacz2VR4gf8AVvdCAffKL/tTYt
1v0ofMccow/8r3/oJtDh8olW1UfnW3rMHijbYBH4HdwtU47hzLdyTSKsD61wm8jZvx7LvBD/G0Hp
1uwJZl5WeWpu/T363vmrgCIeVA81hZneJmh2dMnwyu9akgElsB8MxNnFrmT8uFEBDegLegLr1AkX
VxB80IyGXwiK5XRiiDfPwyOcpOcftMfDMn13wshEc+jrUS4AlE7TUmfYL7bpzj5k30cf5M4nJh03
wHOzhMNB7QQl4YxM35mh1ysFcbt+Zg6YihTqBlw0jZIqD2y08BgGLQ0vt52NXxw5ZiQ8EEkzIdCs
PCR1rqa6FHqWqtO30f8aJT0o0rwaQOH2uj2gHVPkK++GP8QF4NRpiJ4EFIWfaUEGPbbsxffhD2px
RdVP1yLwnm2H91um4p4iihc1K0S2dzwG23DCmkDY+hJixHk2OYJPeXlGr5/PxdC/SAera7FE/lET
JGuYKmWsndXv9iPtnDV6i8xE6M/tzWW5d3PyFwLbwxvCjVmKL1aI+OB/6iehg0uEcSb5sclSz8FY
P9xTXm75LcO0HMu+fAowKd/sr/tx302P7VQR3uSY5hF9q1Km6ygxQvi+gwcN5DeKq32Hpa/T54X8
Jhxeuuj5HXviUfg30qcWThgjZy/Hz3UGpFA4ZYEvAj1gOm53l3kbE+Q8mMlaZ0V5Quut7jAKS0GU
3pYVcyAoFHDAyjhdqTsQHf/+nA8bFFFPE46iN+Avsg2kSwg1xheTDkFvQiT6c+haJN7ICVuVz7oi
x2unSXkdYpblNqOaFFCZIwp3ojrhN4ddm3bCMeqkZ4Kmv6RYF5ggAptWLU82k35nM7iiq0W/Fro4
b664fJEY7h5A1R+USgV3bDhBGnwsUEvOzxYTIFgtcAFUp8+MnHyRYTA6jJBIzL+IKiMfrIJXClsc
K/T6dMPLn/CZE21s6T06uPREBTw5BO0yydGygc2MUbKt15JiUuYejAXRiKQk75ojVfC5zwKaCK2V
c0mxOoGgrArzSMDL2TTJCjVvoSyeYvybP6JirlCE6ZjA1AEYfWA8s5vvjH14EL7+yM2HMZh/dE2F
iET0PyG9myrD7lRFMrca05ksSSHdbYBz3RgCMYuM0h2qDP5xMiDqb3S8B8LZGJ2Bk/ON/96vyrnX
KoNs7WcZo5EJfKuYVaT4otb9Uq7zd9xqQgj5LPIAyt3gFUJqmSUbNBDYppZLf8p8nOHvgn/czeYI
Xfo0aZH6mbmWB1x4zBP+lInQaRRiFpidnK5zjzJxta9ee5+P83WM0jT/Ogcuoh1WavQptrHpNyEZ
4kcXLL+6JaXBPGxqEeugqJ1YlVOrQJgzCJoAN82Xvs2GkmYBFzVPA6z8jwOUxZvAzVWwpQTBKLGw
wji6+lu+ECe7OpOrRTt2ENUuZ1hjFSGWT6aV3hFCdvBkpn+oPCkS9gXYkKMMr+nA//15TB7s73di
z0TfcFP1P5LDYjaGOLWM3MjeDexpSId/PbaRvuV4R9eccS4ODuJy5gnjilmbO4a6p6UZZGlcuJWr
RvLBqNrc07lPQsFhpSEkLaQ1k8oe8rjY1fOvy0ExJqIsa9IrX5YomH4KKAFZMzy0NRclOFhtUA1g
B/eCjnOn2PimyCcU2EeYUsvnzyq15s3SNRXfll2B5uFAS3XFqVdxOPPhKB5zxyiCmkay03BNCqlz
Rh+3oFsjq/DClfoVinFpeCPqjJUw1bHzYilJK+hb7Nosg7v4+IZM6xkQ5WiiTy79+KGq1mOIkPJa
BIaiMco+TU6ZQjX3mLY9ZuDT9ckXd4L5sqNrXh//7tG9ShZKfE+rhq+ZBujhphL3nKIa3avfGRB9
8WE95RYgJmrggTFMxidVkC1kWeuWxn5XUZZvxZ+sS4fNks7KIC7ugDUSbIESqq//xm3r9rGyyJDR
EEuPxkeh955vEZeIGFAiNgO/ojuzV3HEl3qDSOQ6nJXYconuls3erY1+/41YKJla1RYTHFTHbbnl
q6UeUJU8OluIZ/pzVFpVS2e3WQjBKLI6CYxo4EMvB7f+XxZbrXBqrkXJzb3Jg7n9brwts5h9JD3N
GSDffzGKOUZDpVRvJIBeZM0oCkuhUPyUuTKIyyD2BLT3N22adVJwP0BEPA6cprZX5SW00c6KxXTO
T8cOSOs8KvQyI26BARhzzgTM5Rr7YiF+n9YKOxB164twy2mOrH6YW0GV/E87fA94He5ORAwI86na
jecJNf7setnF23D1RwjwkkUODOsQ7BJ5LudJJepQxcUymmi070SVAxF2/6PTb80lVkWOCS+mC0h1
iisCBQaqBCMMYR+tUarDX2BgDl2CksmvCHxpTufmutjrqcwKaLUI9PAnoIXLDe6enMd5yRUTRUoP
v8abtuU5bXu3SctbmcfIn3OshGXBnwZFmIdh5yzIykYRlDoqxHFTQdvvhbO5PCykk+0zAfDspHHX
Y4IvEU4P553LNQJQCP9n4vJmmxIWoS+/NqH9cH/tlCXbg2c7EOcVu9nqXDSQZV8+SKz4eLyoDL6y
v0jn3AK9OIFchipso9L/IKX7L9bCFm4f6iv3i3Bg4PCeufVHFk3rPE87vJf+MO4zRg+0KdJfaBug
6hqugnhuX/XBwzkCE/SlMwOIH1osAVtOjHN7WbO/Og4lnviDmo1ygaIHE1h9hmN9Ea5eJ/6RpDDi
GdZkC4yDr/MXvWOcbbAU06XH6U4hfTyRWvxeueS7RVxfWtkaaaz1WBiIw9HsbjLg4UqX3Wo8NmmO
DtJsSpUZwBEQg3vA9NrVFoEb9sxlFtwt5TMailVPMSJZxFcKAZ7jQx4e42u7I5QgcQbb9NXCHy8K
xg5IJSSK1wUPHpdxge5yaOg/0/S9Rfd2RJr/Cd9vepE3fS1k5JLkpI8//qsVQ9+uZJ9eToSLcHQ9
5jbsGwTe0T5VPdLhtCio/bePf8a0mNaDp2862/mKE6YP0PAOg8kb721P7oVwQcbbfjm0QCfUAriC
G6SD8X1Cnqc+8dRsZ9vsJqbaHL2l/T7bOyby004A2Vp/fnSM2CYeg80R9G5sChzWANGQd6uipq/x
wx100Cuc6cb5/9LmEcgwjn+DRCFsNfYsUTlR5J6N8jY94aDTki6Z6V9mfh5hEhJ9asHHUDPuXCH2
CSexTdSqOyb0rtI5sJ3X9sebXkoOP6e632G03O/wyB13rI5LvOKUzvkQyu9WBpsdXuS6P4NBqBZo
epceqYL6HVQCOtIDXWbOVQxV7cdk18KAuOA/Xnc+2Whn7M9sLe6zeIPaqjrwL3MFLeBvVdnvVeuB
pjfK7ApUsDSux1TgPgPpJTICGFJvFYuO83DXR+4K73EzEA2EQfxZ1tdRcFEr2kEXMRlLEWCMyCY7
D7RlPNQEFSw7p7/1doUS3O8/BA1seFYIxBFiSv4u3NWtHVDUQZgkmgke0hEXNmh419BwbaNg4XmK
0yllXeOCwD1EQ9GhQEmBu1Q7dInGukZuL04qUmQJyvu6rDBfjDsBI/arqDjmIucXoXUQQZcwyc5M
HnH4BgqDnFJHK4UjMdigR2zrRkZCkYLsnk4QaVYyJbdi2JoF7d8FYD+ZXnESxiz6u3xpUM2qFKR0
WyA3QIzZTx510/BmIJaeKUkFoaqHJWfdSmRYED0+as/eFXRGI0BE0U2V+m2mvfk6kfLXM3LDZgQ5
kAEtrnFOca6wijOicX3qZRsx7Ktuxt5lOQjZuhQCL2iy4af87VE3TWJiJdPsZ1DqkQ9Wu7e4rAqf
h9bIPfL08FCTQfceN5wvoOWY8C9cYP4xZwPiTetQLT1IXfkl1KPFHYeanBtDkkjRgSermCqRt2sJ
lhctwqP2leObOL+q+4f+uw4CXY0mTxDsMTQWpjUJOAlt6yYPV1CFh0t37cWCWev1hbJxFMjfyEWf
DGwGPQ36HwOO9jhC954uTeM1buWNsBeqxH995wO2lsrizl61mwCwlq8rjTZid2ek164+QN+Ppzea
nC4hKPCiZElXMekyfxoKxDBdds+Xh3ijgpQiKmwU3BMLeLedRbfRU0uYJlgwoVmL8uNL/RyLmHvX
msKlLHi8pxe/R099C06atrmFJVpKi4bpdyY7777tFKhA8n0GQkSTTE4WvF1ktvY/u/kMUezUTUPF
yLQfYj5jvgqUA5aTlJfCLagA9+tePD29dqZgILvo6KzVi7mg71nk30xaZ0+cIIfPWv+DTTZgX8rQ
sqb6/exkUABpGWVo1z6dtBdb4De6MyEXn0M/8kWg5OSl4kw3iaro/4OTwIBgV8kmCjZ/kLDtdBYz
NO4HnHu0iyqxbqEWbQuT00LRw5UnoOi6EBlWAEBFo6UZW2om6EqsiPiK3rUQg6osnE1chztiqqwY
ky5K6bFaqkUA7cmAh6oGaB6llBjdye331g8u8ohNRbRXqqc5SscSOU7silv53gZZJfR+wgLw5y4R
oHNa7sLCNT1oyoTt3G7iUR7fY0b1ccrIgD1Wh9h/7E0xAClDaDfrwS8ECgZsQiENfpD+m+0pId9T
18dCuX2xmxFK7RhvQkJ0yvohvqV8XB243ZVahfVhcNYaAqOtVEO9s/ExJnSZVnvRUbFnk383Q7sI
ACIHcv/kd96WOqnuYz8kVYxqnkaGpSF0KNyNrW61Zevc0+GOGSzgvsk3PMVawz9VOXOe7qmlzWIo
DeqvBm0aAS7/BypwvUr4jsRxYIJ2ZUoudISE/3kzqDpQYJ1O7oEKkmoKRM9Kfq8AzPgE7gSY6Mgy
EflUKyDURgBj5tx4w61C/t8c6lqnoY/hDu2Kheaxzhx6bvRwPRgreoKF3cdgtgXlqn846Ftd4X/L
SGf/0mkYELyhO/3hJiWv9jBFEsYVOkc1kGasC73LpxxAEqHHIoovT4m1U7tkfPBnVpM6vP7k9eSQ
pE3uO156fSSCbOa2B4d8bo9Qa7kR1iFS/vtxiFthPJDt3OwadE7Z1wHjjEgBx7rAVSDeWJS3ra+U
6c2wQwvzZIXVSU+P6s2j86lFHs63/1kbIAH8qE01wrFroirPI04o1TGbi3JSRwvHW0bXeAq7/n4D
d3R/3GnEILzXcYetUisz9MSoivJIQ4pafR5zsmhbCDDMnX8eTh+qqWoFm0cVl1mKYFcYNs7OQ2xe
xpSAUJpBUuLkkC3SDR5GV3PFXg6b1P1/lrfomABAMMjJiejTYcVEUZH6Bf2kaJvxLhqOJ/pXiWQG
5WGGGADDXyzsID3QzlW9eKeWy2/nyPVjO5P69TaABSgxTjSjxhcAGP5kA0ubJasTY0iQ6YxhjNWE
pg2BVGHOtFk71Dy6kSL3Ckngb/RmWz+3DJIiU08gHaOA6YFEnvzxee8nQhq/IpWp7H+d1GLVdQx8
46Q2XTdqUCkJhQZWEFJ5TR7EUN0XwzqDB6SbeJaAf+MZaQQ//S2r/Sb4Vdy8lbp3xkYhfTnAmurY
maybNsZG8gl57pjuxw0Vb3C2pSU+KQO13cN16Sj14+MIU6RhiUpfOoWoHKgSnB9bs0wzrbLk83G1
Gm9Hwq2+ku13w/cFBeL7nnbWiJDs/3x8YkR3e/Dt33WNs5krjGlxs1CD9OFrNEToYtKKPBt4Us0E
gziF2Qly3rsAbg1tPvKLWs2ULA6eMBz5wJZAjvhqw5BYuvWeSO5+ZlbZuN/ZBRP9i/s95EGwFNmV
flFSqGee/HRoww/x9/2F5b8p4054f1UFyXkBoYjtF6g9Pt2LNVkAsrkjOinkxfBjT+YTh/ZPyblf
WLIqNccNhl/T7KV20afk65QUnh5B38GZiw6tfrSEz3fpkWabssgqLqA6yngrc6DLuYHpUIObBgql
hLAAquqAqVWMBRpO3tGh+2Ven6Bunj+qyhULUbDnfNUdxsAbUaA9xr+EPuGq/kPHRcdJzmmY22tZ
Se9J8jduPk4Q6nCpGaxg7xcdIFsh8ZHbJFVU4k1G890BZ8A+xvjC5tsaG3NnrK9psgphSaUiteZk
jYxBYqA4LjgWLCatDmvo9KvFVe+dp7qWuH4ewHmXaZeMSIs5EBIkxm1yAjnM+sNqQVlXGF5LJqQU
uEC7zWt6hg1B8odcjVAhPC8gf99HMZ/W8/uBzQGnlTKoRnkJzvQurLFJ9DTNedl1bbLFzkVsY8Wt
f26KxLM4TrJVe+J/zF7176A0IwPfpZQrd+bKz2eM6b4R7/nUPPIL7PHnkmdFKE1u8OOwyU303S6g
Ga3WIi6LzPiyMBuBtAUJqb7FrmKiiAiRMyyrFPHIRxz0SstOSoYUbpbR/Bct/AlfTpe6kD1EO5YT
3vl/07TZmCmQLolL63ACEHr8qFb50neb3pWxijEWqgyHrr/RzpA80YPqJ3NbMe4y13nnhC4RssLm
5hr/pL6V9k/QV1lURix24Z8Y05N+ocMSRzHiKEZfFt6efX2IbE++PdtYoJN8oEJOzknqBUmcGoah
vB1wawEHF7R9aRQlKXT0ac0o4WhLRQkxTOy0revaHJx2Ch1CaGd+wWxDNWIJRD9K2S4ZdxmPC/t3
D7rciaxHt2zb/zWCqLcrelBt3ekJFthjkLLo7RpYG+wRc0E7a+EBFD1mcJXWPb3WDKBDZ0cKGFFu
9I5omgUOCsQALjD93DPFTZwVFAW8vAiG9TDKrCtf7SbUKUmccA2+JXB2bgkMmc66tKxdOBqQCvHe
g9j2dDDQOlr3PVnkqFAgw9PCuHtB+NZrtKkQ8I1l1rgmsymvC8MFfTFBh3GLRvPjSekmqLbNPsI9
g54z54KT177RSfUq6zuNYS0gsDHdvtbM7l4+GGkZ2S5SOLF93NX1OSaBOSjLCGP4I3SZHM4nOR1r
LFE4/QuSJPPUSl4OZKAuVX79o3aZKjJ6YYCRTBk1xLZyYoBrGYs5K/oy82NQn7XoanLweIwPlTew
E4J5hrk5JM+OmGmPSCb5pSLtaKAm2WKBw1SvsGnEv2xHQcgcgytVhLJtSjZ41/2WFm2jdzwuZ4Oi
1ZHMLcX/WH/E5pEyY4K1ORI3Uq8wgQqIWz0YGeaT+Ls/0jZlOHzsaiqc/0kAwRXH3hqZL+MCutQ9
2GBCNOkwKOH1YSD/yKnRBjGBOT/vRMdg/RSMy0k1rGa5rgg9VOx1hYn4pMndl63eYsYkYeHo4E0p
jUdzqjGeS8+PRMKjspn3yt+w1RWAZm3Tn67RHzp9gW83KUMwW8AISJexZOHxrSuXFKRlSwoUI18d
hqjtfgXgaOEQeNe5vWGj7NGEytoHUyAXB0tRtFfVkMe4gdTPdmmBj3l6AjeJjsnYydSESS5YXbAj
lhq12BI2TXk6S8pklkDZtKB1dMGR+GJoTYc6HBBPdalYNyxH5xrHun7hYg52vZFkdtflkwjRRgsu
BREWef0HdV+se8E5BLeHpR41TlxKLAS/DQv/q7awfs5YtKSjfy4tJAwmbxYBLeaeX7VUPjbKZ92h
THpd+PUUbHsmcQiDtDgv/MxjLxpsvqe0PRyqOmYxFQpMdQdaV5b77WE8+KsIAFH+OQWaCQOAiWGg
v9zazLPrYFxeKg4mFwlQHg0a/Gtk0l5LRQqPFiP+lEJS8ZeKhP25aJfZk4htP3DoCAqBWIpLWi4k
VeHhn616a2mMa/0gEdfAKc6e+1dpqbnFyHAgGdb001u1stxwz0QCoWHx9htCQMb4Hlo4P0scpd7w
Iqscd6ubREpDqKoWp5kPZkLedBd5LwmQlwuOkZDTkYYvNFuxPhBCDmW61KXNOUBfTRjVhfOMtOVU
E4YFE8H/NOGPBC74LyQAXvBS7olttFJx2XdK4mxVadGgM3dsGZHEf5P+gHDPU4nUrYkYoCYP8AO8
XyIdrCcE/PzjHDsWw1ePp0/1jqb76zzap/yX6xDq9G90hhQpafAHFXJvONSTwUkCXYaL03/cCthr
yGmyyulhpwyeUx7QhURoN19FDR4dZuOP9HzwrTf3kgzAiUrLF+6wuxjf8pZuhcWqGodtMKpx063g
HzyR0GE0WkxEenyEsp+82BsBYAbffAuVVHppdX9yrOceeezIDyBCSdAFgG7VJkB3RkEgosT6tcuW
klwAeJMWBTFTEk0KT49xZ/xgAPRKLb2jmAj1NNLS8YbNzFCLg8IvZtEj6aVu6jHV2Fbjhhzl03I1
j48xYf+RTncgPznsrp8P1KzArQ3CmSM82wpgLBnBaRCnhLnKMktMurfZaNMcEJazC7M+3DJsDxiP
LAHJ6dtBOugil9mzyVgy1htanF1+eD7iNNpuh67QL6QomppjYX+l67c9a72PuTuxw9iLJ8JO3nAu
rBOH1hWAFRt/Q/yhqtiLNjeQ+pewvIOBOM8eMQhgtImbMy3psezQbgKc5FgryNFw94wGrNQUdN8e
vsYDLM6j2pk7JcaAPfpJ55/07X44TaWFYl4KAqeuQ4Zpr2FCtEdYDclty/xyQsFyV4xydmO62NhL
LZ7Kn9dicw+z3RoVh5ZVGlNIbZ2Cj/dS5ie/RIye/dnxdGHff2nfs1pQnrvrb32HzOpiRy7dmE+P
bcI2F2UdEEGhW/bTKV4XPwKvnFG6vfqZo1E0EoevWFMExzIBWty4LLMBq7LCEKwXd3k4iCO5sss/
fLtT8dLjeucXDYrA7/DubNOfBtxyPPGCOdfWBq7YdQGbar17rE4Q3/ddcXe9qFDIb0mdKzGNRxE8
peOsa/uVuwx0eYGtCfQVY6VUjSvlNwmEwdlq9vHeQN/UXOPLl/sDhq/KD02cf8l2ZLf34XchI1p+
1QLPAAhCS/kuGgl6LRC/KOjTfSS0NpxDiHI1ASM4+b/5qexPfxL3TqsDBojUUBcc8QNmBiLjwN2r
T30IWo05ImuV0Prhwo+LbwoPG6GcTi4h6c8mkxsNc3EZMxPVU4Ps3wPFlml7G4hHk2N3KevT+b9V
bSYpAsQdDLtWZX9DmvmrTwITbHAu5Pq726obcD6nb/1cBRIoc7GMBd69q43hzhNhErWbVRJpfBWY
neK07Xhgcmoy6lSmHGbPQKMqdBuW1X/Y9nTD2w/Mgzx9Y/+YfG6FteWYZYDeZLhO8Jqa8k9bPkc3
jymXeKnc0VI8/SlfsxpEenEmVdJeaIJoppdIzM/ZTv19bPrFCnqiVfhhvfH/8WkyeRnkPejAlZzh
fxS1etYuLThN1Rnn14kze9ODIH+T6JZpLe6SHYdZgdQbnbiaiOs+Vnn/94KBfyZlaC5r4jiqkVB2
Lsk48Ml6kzMWqT3JhggWs3WGamkmOSdH9+tusbbI/foB1M1h8cy8dzgjDvtObyeXfw+SmGxnxYIt
+y/dLsYGDEJpF9RFiH15xjQlTQ4Dj9i1qEhUga9uGfA5B5ib8B3CiX40ieGEDN9dPuBZabxslFtX
7ngY4p2o++Enp4F/yK8T9seFKupxDhPNMPf1mdztBrBWF9GRzKddJzjLeQhi6C0evSlTwOEp4aO5
mE8dNFABZmyrCqZLc2XXJeq+YxtMDS/N22/Qib1zFOXyXueivJ1Q9RqD6dBNmlrVdGoHf8Qdrs3M
5HZzDfzxL3cAX90ftfiOgyWLEOMuW2Kjrot6Z7PSHAgcj1u55PQqNnE/7kaHzcn+iTkJQj9lK8tV
KtfukuwQypi5JD72sH0ollciSjrsJ30g8bqIjgKNsDuHO/oInJV8GZRKW8H3pUksxXE/XPurBaCN
gZt0p3QMKuX+zb2L3lQOvTONYc6Yi0iCbxFNhogdWm6EQqFPfJM4XgjPp1kZl6OyeGFZEAjzjvw6
plC2X4g9AUu9KH/iVCeWu0AAq5CuqRL7gTc6Zwg5PHvax02D5vCz9uxyU0UNk6W5exwnO4IlxT4K
EAUNNC1t7jycOrBGsDQHKWJySHCooSKlFDPRoElNlXfb0Cn60kXUhG+N4oATnmqFLZ18KhBjSdNT
J1OzX3pxy0KAjtStxaxjUVtMsBkmfiTTuRFfSBIifR14vyfZvDeOfeAleW4ijDrxgkYr1nJAHLdO
aWRLqbzbVIxgCK3zKCiEV1/JcQzopkdyjt4NprKdOzXk3N3JnZifQoRpuZnRbFN+u/OlIv7tTrLG
lA6ofcR7mS105y7mXmU2d20Cb+q4kjW/vX9aIFP7m75Nfu0Mh4BQnXZSNCefyooQIDikqiVXKKd6
K85WGJOnbtTgtF/XjfGOvGxqWvAVqHm+YaoCv5b87wEo6GthQvwhnu9InKhZCRVflG35LVffhJEt
uQ//tfd80pckDHzUnBnmViATHc874G3P1euoKCmekLuNND6H7w6D8jyt4O0MpKwS8Q4fgOHbvWym
XOunZnSiVdH55Wx9juDsYFtrGQJnnYmJpq2kdCDEzmA2an4vEQhJDyy4gI04Ajp4LYW6594XtFBX
TytubFXzCOcO5LjZVSVvHHD8GKE+6ZU/bBThn8qKbbruc01nBN57nvO3NVP2dUBWFj8ihwF0VSVz
M+r7pG3Vb88vwTXAZ4KYGwLXlguHa/P+jhIRRJwWnTaEg68M3vrNt0h7RvlOK+X0szofFXn0WT2+
uka/L1Mg7HCkiztyGYO6VCDv1wXGludJgJNVDJ+93Wg2QtxljW++e8vpbdpYtN1t/DlD5h1rtbH/
vrGDC47rlH3PPV9wnckVd+1xqy5n8FwbfZyin+mDge/wpPMcncm+6ya2pIT0BE7QnwwZ4tdwMQj2
hgnqjDl3heS8GYpNDYcugC4tmpm74YMbZGfJ0g6UOgu3KjokoyOxsoZaTNLr2hXqiKijoMG8/tNC
wwkUpc5fJoY56GLaZMONxVPk5L4U007I4Q+5LMJ6iuPit898MELBKpsbuXb7Uh1RwOK96J4gkgID
LR20j1QSAcvSeALR+AtyE2A7/jb3zqBKNWk4sJ7lnR6Hn7Q5WN3kLJtvhUcndpj9m16aPFZimJLL
ZtBQQQF250b1RH13HLjV2PZCLeJB4SH2YYILe6Qw1WW0u/2iZIbCj902UftjDQOY7RTUoSIzck8+
0/g5FCo+W9A3eSAMfuf8BAOLjtyi6MnDERyN6TnnNSrPnImcioIhFrNu8qQZ0osvpJWJQnq90ISn
rdN+TRghs2Ssd/bM8muQJdRG3xTO182lChuC+aa0Hf2FAXPG6ZGT6/FSByg+qXMtkph0QMC9cusK
wGRcTIx6XWTBYn5wTqr18Cq0GPv9sQba7RCHFG1bL8+RHqatoS3VaJ/5nzI+YFwe35KLKJWCl5Tx
jlRrBRWVT0WXpqnITmrfz2HOhmqzG19Rv4E1KtK+61lNG/NcNub3K4psFaqjnQ4ydVTaLBZdW8s3
r06NSp5uyytYz6P7Pw8OrVR9ZmtXvzr0MF2MkCX7nolUqSOFMPk3Vw/TQu7dtueILb+iX/easJq2
woUbWjSo7gsIv+WdQ3Zy9YDpNwdWxgPMbP4AaXzw5PJVg4yiK8uOljvWlcqmB2YHiAB42pZV5orV
EmWVuocXQvOBbgpyci4+wkDKMrdgGrzlTeweMqmtrP+bRWcnV5YnRG1/aHqgwTNwD1tRiEttH2Zv
cMhsDikZOodgBR+IgSXzHN9h1MoQjrMem0yNK1mvN9EtaB3zGylMR5E3w9Ta8/NSntulb1Rt4LVi
0R3X1BnTmbi35URPrImWVWjPIc9evH6vanhZdw20m9Xywi0tJ0tci8pOFA2x8vWDPOvdgmoAIp9J
tA4zLO7Z7vSaINu/2wqJY/VA4AP4PryIsC755dVTeAWXQ5EA2ltNgFnwjePJGrYrJIOEil0HaezB
7ogSBLcwmCxQZ0a6m2Xm3aaf15lo6TVAst/8x8APWxjokjyW4XCpl6GG8ZJNETq+1zRjRfxXrLQG
1n9rRjwmldDTUJRlgHIp87S044smBMDqTYUDk2n43twxTgechgr2/nyZthDyxD619uZPrrArnDBq
Ww8t3u4aNl+k60KkUj0qJQ2IAhfCKmj4gLkxMAVdrMRrC19e9C/nehhcja2ExPXpcMpYBZ2tG3NS
w29CL+Wu7Gd4PHPlmy8uAlQr8dHoFQZqndB3FNgrsvoj6RmfE2GOd08UCntCH/E0mYNHrlDv7sNr
zFvX+5uURlu9QWGDedr7Chqy+BH7YGJLNZkDUqnv0m6ZEph9uho5tXQprdyj1J5CqwDy5zJz+sGI
zApxGGvPKfdlFkgacdZxC5R0m8nT/mbMUg87p1r3TOBHszOI5T5lj9TRaWLdbyHRWjR2bRQLrxJR
yYHFQ3fRgBpIP18GizL7cI7OvAFniFqpn0YMpoZn5QjBRXvO4bOSjr2BlFjftK1aYbYK+3LgO3uy
9CN/QfTj52gsaqKvE8f7gOGpA9WJuzIi3ysf19/Tb4P3j8APMzUYPJnIeln3M2URDD5haXJD08ow
TkYQj0Q5n5rxjwh5bHZ/4IWYMuxl9v2XJahxujXXrdBCGNjDltkTtiZOIgn0jUm1+kVROg67nrjS
5n0KI/YN9lhWvlc59y5s54w/gjArL3ttWHmw04HsXjbxWcnn3l4IPyHh+mbMNDr/RYgWWNXC/SWj
sccksj3GJW2LxDhpFZV9IGRiGAKYyyXn9dW8KQnM47iErP+++Y40m+1rXmA894OzPUjUTPB7ku0d
0De03ujbQhST4zB6mIycIqV1hsjyuvqAoIOL5uac23HJVNQaMJ21YvoPDSTMHC8jdjoMteqihD5f
jE4ZGXUsu+/zN4SweUvi9CcFG6STmQFhwXdvD/33rJzj8O0ZOrft3T/gV80S4hItI+6hLJEMPyu2
x2ekX7OepLqPnw+GiZSsa2NwTS41OTnKG83M/0trCoI/vMWAS06g4BiapFuDunL55ndt9413pGB4
2L2o+6YtrjqpKwTxn77AvlJ11YmL8QtSLIYX6s58t5WLAPW24jt4BJXpWPOM7p2vqwL0age5UCpF
UiQ2T5bWqLUF2STfXwuj4V8/AT2uSQY8vHdnGBqq3or0VUrQDKmZxTqZ3CIX3MyMdTjtxr7iJkTz
/WXqHpr35clBmuMGj8TU3QFaq56+j6dHy3A7gYkm9TqPB1puIQzA9Ize93hKIUKQj+pSP2NU3IRI
KgjDUK//tzL8pzXQjMeFoM5C0O4UONn7eZhdXH4TsZ0tL/v4JuRvF0SxUMLiGjgq0ikYxcGC8EPw
Onv3SYjHY44ccGmY+C+QXF07iOGk2vyV9ErfP0mw8XfifNB+pLYk0aPo7tbclFC2FCgDjrpXoM5z
baF3t4wji/pKe6h/WpH8zYX/oVnLzJ+sE3t1rDV0pSjQuOTjYeiqXQJ/yjvqNCXyT1w+gdpJep0O
6DzG5qKjyHVMGnd4kxbAM6yJxJn5LzMwZubKtySVs+Yjmy7kwbA4EhaDlSkE9AUmpUmzvd24iyNA
QisFfnQE4vprWIAejN8XtHC6WtWPv6dbvw5GOGohY6Mxrjn7SeDlGmHf/pPpeVuSR1alU3sOuecW
dQoa7viRHA1wpdBSuZzlUz+JBvdBA/4GuO8SwWbk1w7lKY7LMPTIEG9ZkaxDCfu6wszRg6MhKc3q
PQyxaM28+D5r8xH5zu0okkaQKT7+3yCJT0HvAP0WRhn3WNRVGksVy/qt8vVn+jeWzRSB8C3iJn9S
8jT/tcvQwGrAQ9VH04YiZzAoznMbkrYHNyMywNHckseGcC7wqrGscjSo38a+qgRxtVapyGfx191R
wnqSQ+/uHQSbCtxf7feoeFG3R3DuFUUO79YsabOLy4JUecT5rnewXXBBSU1mO7cUUTdt0f0I8t53
UQSHnbZo+z+Vw39CZFo8LbUmK0D4GvHBEyQLzj780aydVdjAPXL8xf76wGxhfCGVOVddJ6BwiLVu
z46jRTcvmptPILWQhz4gq3v8olzx7JVsMYwu71ypA9WrU+J3KKPyLaROU5LBN7i9yqydP6ZLJMnj
hiOzXiJljapHynbgRWWIPk5LArcJbcnKVmHM68TkDTyfWB584VQk/dscDj1I7BneaHM3XXm8WaiI
67ZJwj/7Y/x+q0/2Q27PKAjTxidiIGBD2XvokCaP7QGI7vSlgQGzfDReOcrBzYuIgCzYKXmtekWB
VbGGqEbuwNZ7Rrri+HFP1jEua91Px+4tU8caV7EVIijO125FRxQmzkRJm4Y8yG3c4s75xAweh8ai
h5IZlisBA4NUsiUx2cyAF3IMtfXnwXu+jFCIUBFWMFetbx9CRJMJcnt6uKY56GGMwWyQkO8/Zm6b
YmKbhjU9LDRP63A21s89j710dPFu+br+3W1aSxdLs5ihn86WbRn085P5EHO4QrG8L0OpnkNeiVLT
pcTsVZuiEbGaveFyzp6SlBKUhOtPEJ1KZ9WsEznMOtYTedaRr9PRnBcZTyNaZOt6EFpdF/PEbz+1
c8d+eLWNeOEJ4h6YaF7PL/bt3QHg94l0YqlJFiqUOfx5B2JZweDX5HRu2HRj/DhfVM7xQ9cmpBQ3
3HhQUHvVLoHhJcF7oTCzcS6CHSpW8hJtYm5RIW29CCBxhQyYUFUqqBmmOHJjtujWAIwVf4dQWXVk
d55NqHCSCnMK2bHiWnDBYB0QAV3MiXIZHLoF0G2B/pW0FV15dFy9eWpFYPe0sY58/3gdc10SzWSe
4OgFvFAEKyURTam23hXhA60T3rSnIaFifPn3v0dEFVNVAS5KbnkqFALvYBvOLM/TKqX6vkk1HXCx
YleXH+UWAi8FOfhqa7PZJZqwc1CEpYcC1ACK5PWK5mmylAsIN9aXquiJdmxqVAW3lFj+2OaDpgxX
ZCF5UEhdjyHk3R734SxZPYJrzG0cHKwgRTLeuVnKiXj0JBgGeNIwgfFfsH8G9Udp7vtxxzhyZuAV
6Mtn8Yoqrcjl+8z67jZRY2SxY2b1v2cPqTt3uvqVSiSQEScIwgwq0Uv4hoVKa8gC5yumeTEzJ9Mu
E6+x9JSZ6HJ+rjkASdHoF0qWct5WHWm0DXhxzmE9mlRdq92cPoRaFT0KxmFWTdAta6NAoUo7D+Er
Y/KJtk2wCald8jeGsqGbY71IwwCWTMzx63xCV2sJUzscodyk+O6XSmPpiGjg66uBpiPvEaU3sQl8
2idysL9Qf57weELmMszDbdHW00M6D0R8TCzg//UYPr/zSO/JxuaEPsM96pO3r81fiYf1TMPghh4d
nVyI0XFQqp3ntOgevTQzwiRrlGvK+zoqbn5G+lyo1TeDvYaIWJ+nRQrbLTDVWLErjmuvW9sjHLUI
ruqJQ3h2mWyi+7j/OcCjZbJ+5D1ygJoUpwur113P6N+q3NUlgN6g+Sh38zjM0ohtFsz4uB9uP98t
0jrqBWeMzp14DnElUqJMIkRl44dhtWgrfvW1WFyiEavy0MXthQWszzpKB7p/WiMDwyBH/QmRdK2u
gCzffM21Pnn+hmfrKt374/FGcnES2Sk6IH9UZ7Yt3Cl33bGekzHGUQwb3hwJxwCmywpdkRJrxmx4
jm41xdZsR7JyBG5JVy1/McGHawJQgA61/cuUiOauyopesr5Np13H5SZXLpLgQyCWt5j2L74MGNX5
qc+Nzei4OGQjvBXeZh2Kwcatu7yi2u0EuFlUa7jOcK9JpNxZSLC1ZbRyFuiAdiIzzj1WbhZYS3Se
syLr4QOSja66okI2qyUTrHV6Ce0xVjqdj08GFvQcZ+KfcQUjzpNQw9IKrfqs9Kogl7GXXpaYfjqm
6XcmfVKYS74Fh4G4GCr4yPAGfevzDHBL0bWtJUxqPofH04MZyYszbOpnOvS4TxrHJ1r0f3GXgQqp
Pe1fZboRUCY5h38VUyVktEdQkQObzLTUYlCGg7vI2rOMeKXuYlDIUax/SqAgc0SJTRFg7Nia4F2/
GzncPNoH+zBFoeRxLsccO/I8VXhMPK9syu4Ytu/2/6At07N12JYyRW/zZHfOzRBQBNsQQ5cNG6mD
42Epnn9c+lKEgccabVIO276gjZ25wf0ZjEUVmAFspkTdiL+dq5xAA0x8W+ZWyjEp4H+JJ6+t9A0o
k6085vWrD7ZGxDDzM7uNp/2c0Vli4OOFOoyorJk9x//MMc6WSvJVUueQWMXRuWFJI/7mgyYZW+2d
ka78gwq/SpwfLSvK3el4nLKsn2OFDNb4OdWx6x02LfiXy41lgXQa9BpOPQ0X41g/F3sgckMMEuyG
1Q9tgl9VNOCOUBVVW3jD13br059mfOzwnMAAymcbC6hN1FZj8v+mCqNJ9gpRiMqJ60Tpk652WYzg
uzbqXPM3zRwfJZjPREQn0sUHUF3q4hJMoyBL6PtEPUJZgjBtinxKam8+rnu2FiZiweLSqx3rCohG
lRzzt8s1lnbV/vZl9P5Vz0SYBAi1Ob0R31+ECuMV9TYUN9XI9fEuthxH6tqP+/yW50RWMj34sL+e
r8+vaEzd0myJSc36ZVJeTh/DK2diy04AiMLX80tfdV1C4y3bBJsxH3nyv7G/MB+3t+LoaDOXTjFv
AvcELY+11a+E8HTj26Yb4P6bjsmJ3M/BWK6zW8qNanSH7mL4DsTyPf/AhirVH9FV8G6Eb+nvoNtC
zbtxJzEFtJ5ZiUuLndv2J4cphRvm8ywve9WR42M7CCdDs415FE8RkjzPyIvWHxcqutTdgdVhLwiU
imGlO8YisuyMpd3MDqfYM/MIRwOWH/ABOpy2eMJ3VYqWDtL07eIOhNz9Wa9bxCJW0kIk/d+/IahB
EMoY4ILPgLtodg5CHx1yfxQ2YQoVGOJbsnN3hIRjJ9HgkKmCmYZu9mAv7LgtyHdpTJV7ulFHSUHI
RFHXx4kPYZn6PhUxtIp/nENQwd7oOtmAlhYcQ/ttCrKxwaHFeoyk9arPLc4mFXski924SDmhLpeH
9P54t3vdzewaBlhk7VGtLndG0Bm1CuFCn/jA+t126T9r+H6NrwlZ21RuX/aTINJ8aFDsgJV/cKil
efSaKIP8ONSLxFZtvRPrVJZlzZ6bh/Nkbh4DXIdjwy3zxvjX8y5XwnluSRGTb6RXkUbBE0BcjOt4
ZNSxTvdDKwZrYNpzAv3D/NtS65nIkR/xc57Qnp2JjmPOld9NtCbHh+/Xvwh+1/Kg/UIs7DredQrD
qY5jN4aGKpAvJnSgLh7IxktH3pp1YQFwLsGLcIuTWdyJqf6cY6nQMDd6/5+mc15UJouhakrrDAcX
dX53nsVI26v+UEu3kh9eodbtOd5PG0czLYgZ4A6y0bim2fg8NnB2rdpoOVMfNeiCxsCF4aQwhrE7
I8c6NJw5FLXlupNey35N7E89Wgt32Del5P/xhjhdKhNYRQycU/Vb9VxUTJ1K1HE1Fd15srLwYH5d
ESOQ3MvOYglPrLIVA/8pNQzYxpnFLwfTdOO60fnTLykIiSMcH3mVR5k7HQuWJWw0mHEiNSW+3LcV
aVPN0vIwZa1rhKPpPUuV42/0PI2Cea3lDeCJ069USpQy+G+GlS15XNylD1AscykFZjmOjqWKQvOq
P/Bp4dZ3g60X/Ew8GIrS4nZA/vdcfAzQccTMBmQPDloJ1xodLK+MGNpQPRgwOnUF4BwSxK/OIUFx
+WL01blet+/H3+lwWEQUjZJPmmZ3n9BWXTgr9/NwCs3oXVVA+ymaoOpObgaUCe9OvjuNji0QaS5O
23mDrVV25RaD3Ssjju5bjgyDgAPl/2UU5hixon50X3aXnh1HN+r42YaSRudag/SvSHEzfKNb+lVv
MYgt7ubTKflfe3ttyDWSmghcxBGXNP3Kiz+omXPBBL7XqOonxWb7F64PnM951GsZSfBCc//GY8TC
N9hjx4BkwcYFjTkKca18V6aWnw6e1ml6fk8MTK58g88v9hgPOiBixpsy0jsoh3PcY5W4D4rNjxzY
Pa6cQYCTdZNlsg/40+AioIHy2UmZ81TljT5qg9anylkXc63950DNoXZ7xAZqmQb7ZygPvAAdLbs+
nIFy8xLh2gTjtj8+4cIXTaPLD8pTiAb3dbtxfl5yEcVZ+25Ke5cQ2Qq6CY9ksP4nt77QiPoYLwij
ngoWyGNQ1mpAgGKA/mXs2lFTPWSIkY1uwaSzgBhNEikP8iDwuNuIFR+ZreiXutH+hQA0T0kNUwGu
I9jxZzNX6H07DrbWZT6IYpkspsnTGMzNNM8eRyCOUErycEybIC+elQisEvgwrT2J6XWbYt0vmHrW
zsdKMY0TixljVmESOCem1Wz10vKlfWpu0FGeJyE7qz1UcU4AdyAoqN0/oPnSyKMrC9CULhzQ6jCt
/CBGLdZ1hnBDpDXqqjntXgGl90WH+4MlDIlYNPrtaDHbbdblReMeGev6BKQoHanfyl8suLow1Kj4
sV0jEgRqst3sfXcnmBU9ZQ85IcAY3ZG4Gk8N5BXF8L8j3bBFbf20cClTpcMR0vx6kIAlcf77dR+Q
zy1qiyYsPsTIB7au1aVHorHWbYhWY9DiyZhDDlSTgABPyQwpMFwY2s5LaLh5SwTnmIxoIAXQiFfw
m6gyPZjBQGAs9V9O0joaWOKTKkNl6rVAllI07HWFcy4u8+pTT5pjmnhoIF7TjDjcP9Hcx7qPbgDE
qsZci0U3tbf72RtR4MXGYPvXSoFv6bDel9G0W8cEYbftFiKpWGWuZWzQWpxte+Hww/owvdGj+bjD
kQQc2tVopb9phnCGHBNwoehTSczuX1vpXTtpaekvnYqxorr15th+eBLgbUwX2AuXpbFo5q+X/ySN
ZGWA947P/6MUGpp7Z/UvXqI399d9qsMh/C4ZsqsaDsBvatjsiA76mr7+QatkoMqIA5ud94WOiIP0
p8SucnbjFt48J9/DBw2chQBZ9R9dX2pIhXP7kbWEgG0VRLBqA0eOgnhFlI/mi9O9EyxeE0GYYzxn
40yvbWSmLB8pgsLvCwrqIrIHpFoAJawTu2iSanRSFE+opiJ9drsk2GquMag3ABaqhxhZRVcnqiJ6
hxKIY3jpdlbn4RXHlwqrYHIgocgnHflU+ffKXBz3uA3BSg3yivBRE+mjKDa0LJEEKL0OS6VoR190
5I2OMpAgUKUXPgb4V7B1ZyEh1cmIlcAopUbKUshZ+9tznh0gnHH80glyzRehWkQ2+FFkuRvRyTdK
DS3xgA8R3FMNUZPjxP3GfBjJnY6BvNwwsUSBZszC0LBoSJ02LSsJyLGJwNC8QlP+xMvM6gD+vmrx
whCEtHMSZ0rqWmmTw/1BTGj3C3kYm9SMBd5BOE/Rf321bBs06TQ8JOipaHqFjiwnUAeRTPJFZzyr
hr0r9MRxu/2RIVma62sgm4Ulnx0fMSA/kb4KT/pdn49NIb9HYnN1GJRkYZeHfTdT8Rn/yQiksClt
L4t7RwMcQ74856ROgX+VWHXbmdK7a3/r4JZiE/XM0oi5oTnJxd5OYiYXupGOXagVYemyhn5kgGZ6
M0DDsHVpIRTXPzJKyt8ht23Tf3pm/8M+5k7Yyysk022QsRPYEiI0LTvLOfYtLcEdQo3noKJNtcRI
97QpWbmA7X2GqyDN6rXj+h1c89TZ91mSb6G4/aBoS/ANEwBTFDy554xad1s4/tNOPej2QMaOO+Iz
kOjSTE9jtjFDVbdq4lWp+Kug3DQSaLEKnsQu0/j1WvUEP2JsOAJV2Fhxqc/+PTizeZh+mkwGbZ66
e+UvG/yXkx0G+ZtNbc4+UOKdcMMs0BxlrwElXEk+D0+xUsmAtAzOkzsDUt5z0SUMnTvpU5LRyOTJ
n/cEo7gw2kyddyTrL7oD1o0ZR/KoMYXKxK4l4PG/r5orSYwdNwgPYjtB4ycQebjYYeHVfcsyTCZg
EgnaL/gd+EyCfNqQVTAjYsAXqC0wkfvvyuww3B4Zs660JimijiP2xuZ100B28md7gV1umbYCoWQW
rOJyCzNLVHHUkNVllNStCOBPsIW0bhbw18rFZrIXj07saAQomfLCFUZLyRSm8wKKbWnu82USRfVf
g5PqBlnPxjxfgwCqANxUp4UijbJ0pIKtsuJtU82pGKILb62RzDuPPpqfIwia++eZA1VzyVHnhnqu
TZRhplZSSGrJDO6YUyAQELVSvbJwXmxtegrPBQbPTy8BQCdxhTX0DpFEVEuZ3b/ety9KpypU1Xjk
rtV2Nn3a3xS/A7Ihfn1sKLxb9fTHx/Ij0r799QT/9U9FMloQHHfzbbuWotfZj0SVJuwvnJyEBDtv
mwwAF4IcbyZMrhUSdgX1azOP2ZcTmldSUrJkgVzpDKV5wIQrcAB0MSnm36zzslKrJKGaFICQGNeI
sj3L5h9ZPMFyjqL3Y0MoZTGMaEFm34VrGATt1wr68u0SPCbRmpL9rM9TwhIAmVN98QtHHvypu0Sd
PnA/BsJkdQa4hZld6T/HlO5uTm4c2GUjx3whF/IrMOPMujKSSJueLOapPZ6CHYtbSlgrKFxCq/Ms
xD+rR7r4pbMAZnLzrURt5A/G4UAQtdEnOy58x/Mraem/zM6BSEOVHyvkFI3GIbB3dNzeG1cLnZJA
vT3xh+3tm3u+4ty5douGo/rdlvPrQwSzKMNXHdwFYjzyUkKhB06ZomQ3L4plaxkhWBTSiIwDroT/
q4YXEusexiLtWu/7R0Aubowt0pGK4THLJj/dJAkGidBJ3FY2lKqxGsRYJnW5HF+e3nCRZeW6+46n
grkJyHbqY7WVVLOINHq3Xhmp4Spg+Tz9FbUtJG4RY423MGCaYlsNZUvKn7InhBdAnWipT1aiM1pc
0FWWVOWJoS5We2JGxT4TZ8petCoh/qqz+zTWptZt3RlujjsYy7DLg6gA/ZtQ5qzPG3vRjo8oEI6M
OPSOC/y983/npVqLV22Gh+OL7D+keAOEH7PNUKgLcRHSZUnSRzaWnBP7YpfB55wsqIOqgeRsqJJx
G6VqOmxwthRYUf5oFIzfzGxDBpfEKY4nj3SWOs7Jh2fHEkQMypO+pKOU5FVXf/J0B1t6XYq+9Q/t
xaEMM2iAeyiuZS9pdnhoDLi9XkSBTzHygWUOpuRwTZxXnCS3TB1BNLjVvv8Q2MGf6Ok/saBIyM4P
n0Bp3WQN90KQDS2lP5crz8PuQm9cqrHeC0WjtgLtJt4SZTVAgdMB+xDyfp+3KsyL8Mal+p0r9Iy2
mmMDRt3WznhurLhH5RhbLszqzxjhwQAWmE6PJVX37UDWpweYx5e5vUkJSGZ+rhcJKKili0hQ8uER
X8Dywjd+Gy1QI3N7QJhBEyNX1u1mcQQmntpcqazFf2Xv3FC/6ysR5DjN3ZKqNVQBnkOZ/1zMQw2O
9IiSmwyWy7dxI2hOZ0csEInAGU22uFhpoBJngjwsDRhGjxYkEtwgLijn8s+aju5n+xObZOW0oJew
yNkCBlbvQ493HlHm3ykC+zRHjsuqiseJxaWDConzTJ6GlZ3spY+uDHE2MKZ4VhOnk/Us10jMaRrh
gKUiKXexOxd/5VhlHP4rnOMJfZKy607kJ9Scgg0SZ6UsnhX1y1+ERSSF7J8UmAJmvcKRptrH3uYb
vzLhkSzmRB6ghLz5pE0NnzkGLM1JHK1CLCxY8DMotshvgQ9lgnqV4+2qPriIVbmRwfkEeZYZHEVN
UcFU3dOKRZQIPvLGkr4M3iy0WjdninF5dSp/3U9NF5o1iwqeQL46eFHeXCKhz+cVrmVpvtePDbex
3xckodRfrdSq9Ll0ZBvci3gp5UAKo9pWt38U1FHPVAPW9l/u+TYQRt/G0UdbR59wvOqdnlrV/DvA
XO8O5JjslILPqZbhGeuu7r2jTUfc4aFRb4ogAAleiWK8JCJLwP8GM9MhI5AHg3qELULIGvYsVVvh
akZhBc2vUcPTEcrg625K4Hpv+IT4OY5m5nvV8K+1BT/amG4JSehZ5x6QKcgw0iK6rH1SFeAIthRK
Zbss6xbVLN1Vneb1+lgfzrOdp8iKyzB6mgrqcIgKFBe7C/XZU9p92h64NTbd2v5c3o6TjMIAUVmI
dikrsc7B0y88LLdwXqNHhmTcE4AcTXPYkfTO/vJ096keTzhl/pgcjlq0wXPUL9mrIZ0mVdxKhe3a
7500lyd0w+ib5akD1qWROE1xltkje73z3WPom7I0DpGerYslzoH0tNiLNjOfuGOmDFST9Smmn6m/
cjvIFkp/443C28KGgwCQLUfkcawwXj9UOpWWGVNqyUm+Jjln1+AbhBPWu9UX0eWXgAQsmLmLwGAX
WRKu2vAvtuMI5LVXSUcsCJldzRJ9Kk7V+FrQJAXlE6uw71RakOq5N37LlAWYeBKIZMk8sdOCv+Je
J/9N2m6nv1jiOXbk8KNhzJvEkeUxnEjhfyr8ra4963l0FNQI4ejxO7IyS1Z1dEyZjQrT1koCdI2w
K5XDiTX/wU7m3tZ78aY2nIFdwtpejll1n+ZYNHedGWgkC6iZZGiE8HxEinAay1aeFRo1QU84NpYW
KJ8tkX+k5HGbwbHy0phzprwCwW3q8ERNCNaG+PLlKw9vtxhTzhY9LmeL/Nv6DuDqgeJnkhK0jlc2
Xjx+8XAmHLWJ6TAp/fs84WJDqzw+dvFUz/3tNOahCssBlYjealth4xAIwF15MR9YnWyRBIgPNGwK
Q0EdskTOy3LFKFBCD7d63cArIHXlQtH0l8kbjxp9c70vUk9cGalDmYNOC3tmchdaKdBRSZjzpWvf
DCcbDjSfyTNdT0V9zMiKhZ8vWPlA8cUFE/JsYbje2KsnzobzWyJdqe2DJuaavXn2SGUN0rkv4pOY
E7ZkHEjpsl0Vn0G/WMdkLW08nBO+9tlM8wfBavUfDocIYTZVTwg43nn63+1D8whVTeybpdN4ItNv
zX/s5XKlO1mIIUyF6VBBSpbjEYtfQjIX/9ooJsj0kWXFvmlCBwyASJm6F1+mQmBAmMetlPu5L6se
knFGW99eYGv7vc7V/pEWcP8YEuoQnuNDY7XRlwqDQqFqmD7SYgOG+Ii0u/+eVK8SXYGq1QpaiUEG
UgOT0gP3KC7Q5EK6z7N0M3Bpb4B9wFqYtsxdoy7j2T0V5iXrSfhLyRHikAyU+edt6wQA7UzR20FR
pxI4S2Aat30oVaqb3PLlnmjv+yrrzSohXPvHuw75+NdY4C0gHth1FFuddUkKnCtfSbXXc6qbLsn2
RVc9TFkTh8QZ9a+ADjesAiKZSZVhCERSz6nLtf24gSuj/azKMD3EYTQ2mLdMHWk98O7HvxJh+ewo
csmEnee/KTei5u3byW1DuYbyEKzRaOjbyt+F5a6nJ58zyQxz7DsHRGENYyWgoPfgNsC40gge8Lv1
m1uiGwCNDfFkGjQSiJDvbXgo8nWGZlbfabp4pTObrxdxtn28i8rdM1sK9rOSUz7xWSPT1ZGjRvli
DjsxcVPi4jcFQfYX8GK9uJKDbFrYbko9lb1BgvLa9laayoOcyvE8K317rAbyNAddBrwPHXzU806a
8YyjALLSYOlTZoHecIvDMgkgZkr0AH5f7aBJHyqdDsCHXQNjCti8U6B66VmCdZKQ6eRiFGB6KWP+
z8eckyNRPIjftBDCmJCAbpwiMY6UKTmaYwbQfRwsZdGKZ7Dy1bhNkHEQ0p+tjA7EO6eQFW4BNEt1
qb5PyBQYEypeuYDQ6yD9nzNbPmR49mXlqqFfn4tCgS9zsJvzEXQ93Fp2KlK4cLKAtXz2evGq7BgZ
F3ydMLoyUT21n085HdvDpwIRq/z4sJt2kl01fXfYPQS5wsnUgwjSrQoGgQTOjUsiiyGbhOcetsi0
COIi1IDIiW2BjhmS2saytrNb3nXZukCwTaO+LjEx9SBB+9f2UwRX4HqduhMVe3Tv2DUaDIwBKObZ
HX0x8vQDgy4qzg9/B8+oYaVmLvOjb0vHnBR7GGH4fl0BiBqFLB/me25rtoLZEbDxjez6a9whl/ng
4ecVJ0uwVtgmEeEFtG3+40NtOKjhQUIm9CkR//a1eoMnlC785KqGN9fPwykzuPcwm3LVex0vaLeE
jM7O/xlnANSrM4YCqBtYSfizshp1/hveFemaDhK2be4zeejv3ui9GcwzzQMei/2tqTjrtHuluY58
SKbwR5r33/g9ZWGqdmw/NwZG3bFyHx+AYa5xjBmfPYr3AyHZMkJzcstUcgcmv+X+xOxLOVUlrw2n
WG/e8wPNEYPZdObhWsvYtUmWMtukz4JfWnmQnoFl5SOSVWPdnTCFz/oL2J6kKMZ2PK0jKhnMRx1c
Oy/LB/fvdSC7bI9E+9g9aEeALC+brZToMiyoFI/Nj6OJpXjd3hquCcJJSTUA7yM2jngIwIWKg1n1
P9D5aUWlrXcObN0vAOEDa6E0dwBCsFTq9Y3iHhQeMftRvsFBsbV330fpLMrtcqWeVhL6cy7ckoTm
8w5t0LkpGf8f0AvNJzbgBYe5SpuVNkqlyQ5xrBQYYwBdzMG6dNA5jIs/lTPLHIYLG737khElF7Nr
f0Rhud7HXjG9Ri9HXF39zwNeqyxE8VG/apF7DqiALionVvOYvdffTBipr/CZb3NKMg8dYgYuxxxl
I+zGvtPJRSn8KJSm1kqMQNHlHzPLj1VxGUpF9IZO5chxI5UCk1sUmhDD9p2gBFTVEnTAWLudEpmq
ZtkNnwav5BPIpmgXxiI1qjwjdO9RfNwA6oeiY0M6MUfql1X+yhGCgiMuhUvqVFDFBDGPj/qEE0fB
YWP1D24QwtGCup4sxP9ZeE1Ds+aV7vHzALSbT/h0VIblW7ktIWdQaXp1+zNf9Gz5b0EM3p6eTUuS
hY1wutTT1oecj+erWNUiQzHd6n6JfFM9hMOWOSd2hc9JjWu+UWFK+ebEPGSb+Yg38equT0Mz0GAb
691AYS9C94TrSvCDtqtlpLVBioPvsj6QLJrsPLboLG73xu1r3i19y3Zo3Mi0xzHNdw+WO8Kr9ZRb
fFWOL6QndJ7TtjTEi7tWtDLdBrI1U+ulx6AQJ/zMpFXJmroLRX7IFm/Xe0CosT+iX9pp3Wy4YFUW
Wu41Tz8aUFXcpglKiu8Db9sRxA0JvEK4R9KiZ3N14oD2cSdWTKnqjGkUpTf3XGomPf4ZwNcwlg4Z
8taJkYnrXO0JuN3FvAp7mo3UBc1hRuxYUR8ddPQWKlFAMJStFBcbowKPrnTmfZFPswf9PGvZiNVD
wqPlXrWdW6ywjCACOMAuGkg7UGqGD/5XVQHdRfqnz8qoPXhLNcDp4um5Bvh6h9uRWXAvrJ92+Luf
Z7iDHt3Ha9oLar/GHbwqllbXHssH5GLD7ue1FcE8SNURxxQhVW7lSu3GtnHnvW/RwCym7q8TtKmb
wwTC5hg9uQvcdQ8lJXrzPADTMrjzcfFmKTwdOTRekkbPF5kAlcIHji09kEUv7ohh0Nn0FxZ1lmSy
taQUZU1edFD4lkN4i7K9v9sgjDvT6hLXk2Xsr2W/B5iylJRO8CvlZJEMKVWFYhNE1B31+PQ3PE8t
0O1QYSSHm31m2P3tJninS/ohQWk0+3OwvLI3ony9W07jKyQuA8KjeNA5dn3Z+e8V2nNqBrovDQwc
4KImp9ierWxUsaiE+1mpfZwYi1SxYDVonzfGpHa1hBMRGfBqHqKYWc65Y50ZFdYCDnFvHGzKuZXc
OwTwgzo16bwu1WQWUf/vro5gRSyriYaAgrnNRrZr3gZ59ITz1JCh8Kjt74nbOIZUlIpnZMKE9B4Y
xuGscnwcV5VzGKgTT4PSGjzkDt904XJnagNz8vlF5piXfio78CDp6lWYenuhfL1NpigLbUg3Ry0q
f4Paeqx/DAOTsYiByEznUHKXdkXHVW/WczNkHFQ9e0h1QT25rDa1aw3OSxwMqloL9lt8nKKbqS4F
Fm1q8A2Mw/GIgU6RASmhp1ws/LuYbC6bHYc13QWQKIEHa5dgYWCzE1K9K8fLeAZi6HhwacXP9cf0
vY9LhV1xvYYUuhylyK1DWjX9mLixoe8UdeFFrOTFrbd21xzLEYwg/Zg75Uc3B75ALzzmJvp4KQkJ
hD5bMvO2z+BZ+nKT9MtVfFdC7OQKP4FAJpYLD6Y5XiHdf4Vm9uX4JvQtV/TrS7l5849+9ExqAChO
UkW44YaZ5vb6/chrloG7tfTwnvJEFrIiYa6khqI6VcxqBA0GG9vjIjJEu0MTo/KWJadm6bCRB4XE
EXaQaT1N90nqwsYneW431rGnF2Hxzhstb/RGImpysIdIYLp98sGjWFXPJ3N1eVR7aMQSVmWmXeHB
emjx+4XA+IUKrd5XAILsjUZMSmHZBKIX22fKJML7kacBFC4QdacKQPePbhF9eS/AAV1EWjsS87mC
VjE/M0fw7D6hRwVA22X3eQY6TpHZLeRaFNQqjCwt7TQEGLDm39FuiB9XUCMV/TGiSA9GSXaEGxok
ILwEtjeO+tP/PB0ZRMRuxG7eK3DhO3DvpUn2sgNdAIKlm8XK0OyK0lS9eumNSur8B6cMn24wDOKB
o664rt4qWwLGARaJR7TreWRURAPJgmjnGDjWOtjUEdjf2P2zASKphcEgeTPMEma9/Bz+P3t4rk5e
nERvPiLNB/SMoOB4nuu6EiBWse7dDCT/svNaASJtu1s2bLKG1DQPuHvwRqdNTXNBzyqgXcdctwiJ
B7LJ1ZDnEu/BAgxeARF2TGPuVmZ35+Bsy26tlUJTr+FGJ3rFfoIz6S+ZGokIqZnXb8rGJLFwSURb
DyLSZqy7pay8UhFbh7zd/hwkWSUDTibQHUVJTTtWeaTX238D4LeDOgvXnyhiQ+xNKS/btk8jjeya
03n5Z3Ba5MTedOWbnMi06eGqAFZepoezkNlKz0EwuWZg4V/zBe92o9QsfeY9YWNmH/e0NLAPE7PZ
UzG5mpoJ9OZ+U1hWSK5cFCisCqNhjgKBQY6UlDcfcRznlvp32KJH0hMVxgXR3CXy939eipJYqexb
yQlGNGgi7JW3jcWQXVH54QT/dkCLVigmJdIr6bqsaN47Zb2chnKYB4/bTjSBIC2ye1gR8mUk2Pq/
dT4VNjrF0UKxu92FZpeogo5yFEu4Sr4w8EzlBGu0q928epmv4/AlzeHZKf4WgBJKJ4DRou+mYHO4
WZl8JDKScyGeNjuf6Q9tS4Y00OFUUyT/xAjD4W+A+h7oYKnmU0N9myiyEN6RcsPgnWRAUMJKk6S5
hz24/fvwnPuyEnbkuq1ySv79jf3M+XzLH+9l+ajwEYOKkZwndCK74/yt/kwj0bHmsUK/hhNscf8N
u0EI2RMjEsWIIZ1T2jZDtG81vEyd+xY5CIBEBjLC3zHb1DztGKxGbA3xHi7ykODYTB1lJ2CSz9lv
l+5DZXaa1fFR9WFDT0wPGGpNE7LWcLEyxxudcN74Kym2Al+Sz89xT4y2gM3Abf5G9c0V8oP2rFYW
QBFXkRxiRkzRKNLeIa0hEttfTlixhmMfuMm4F9Uu7GgjEOod0n/nFC5gD/sKdZZDKi4ovux+U1AD
snaVe235OX4SiGXnAtgl3AduTOj6zdu4Li/98BDUdNcMGV2wJuyC8hT2Ug5dnUL1RCCW+pMf7geh
9ScB/juAK+IaTToPYUexj5DYhB30SeEhPSfom9wJl4YqtHQDlaaEoDCNlfDxe8uSz0T1c5XO2uMz
jVnn9UA+OcEIw9gVR6NvBc/IMbO+V8sk9OLO9zSvPWn50FwQhQOjs5sK9ecXl2TjcUPwpSrgnzgQ
s027pRPNAGLY5zEmoTMz4/AOunjTBah2EpMkoxBhueR0uC6Xg746HsE1TisJFCL7B8rAPNPfVcdL
+aQw8w2rLprKijbofNzHiM11aJtY3O4j7TkcYZqHPBUNnniIXI33kJ+gtOxMYUCs1vAYwhPT99+h
268PZwdoKaVdqkDLkgLAPfmlpX22YoeD99zJkZ5Xj8j9Cadp+CRs2If2W3Rnn8lwKsd4t1HRCA4U
vyaQj6TdBQPbDEVC8BSAMyu7ypxHcnjYjggjEIIOfBMN+Zuk3sF6tb0cdHKGbkC7hW6Mv3sz1ZE4
9s/lvhgo5LGoTYpyZVJO9PEQ/iDotHpNaKS/y60WNqxN+ZukviZQkusyIf1mFYSSA3RhKbgq3c0F
LlfFPrwO3o/RW/0V+Wf8uxrrwRrMj81EorE6wdo+vCA+raTXKx/fiR7kqgJFJ/agWXEbnU0DOyg4
BnidPzL9x7w/9tKocQwBtpUIICW8qbH9gW5rqXZQKSGqy/WKMSBenApYprNlz3YcYO9Umfq1yKn7
8Uuxn6r8gXGT44PjUAPRyPsdQfcrCQfSt5s8mJf9oby7tb0/4wjsKvy0K2U6eMNd9vZApzjwPw6n
tHemaqGmqPkMJ1eA/JItt8PraS+QkyRYimfNdB2/1vlF49YtTptRm2IPeNpUR7fEWgZwriq1woTA
CLiHE2TIapyZanC2Kg==
`protect end_protected

