

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EErsftIDJVF0m0AzARUB1bTNfa1D65PKFzXVCO3IcVnfdNzarCrieLdbzQivIMAadZGQICQFGhS1
QckM881Qig==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oVVLyVCgNzQviLS1eG+3q0tFr/JK9RCUE5+xAA69a5PzCR+NN1kdZCFY3Hih5lupWCZCqlSR2yxj
T/gFuX/P5PwLJG5+6QmvoI5i4SAxY/rHrl8XM8Kicu6z19CTYp1SPiJ9834l0f0lOlXlTmn836kA
Wgmrcs24F99177fCyOw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kW4owDNqb8AMzEcxlafWfz8koQuLn9mxd/TVVOMuiv8YQ3rvx8K/DGu+WboW7BU9KyEVtBG1MjQH
gJKixZB+7AY25kT/0NwJhM5YyjG4KdEl5DSZuDhsBJip1w/5m+kP4N5/vcsnGSfB2gcc5U+hEZN2
tOLv961hH8596MgBAeOrfvnWa5SH9SROtve5GcJIcP2+J4rtDHR6wFKwG2xp/9kU818nQ53uY3x/
7USyyE73h57I6tiR1+FD47Z14CKQGy+J0+yoYnuxOAdrlqmEtQAPiwIuHmV0R7zwgIucScma6/i1
zxERzOQ0UeBZqrcJuNAcQN3PnQ03sEWGfc4Qwg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iAL6wKTA9iQaAsMi/04OqmErqGG219F3T4DtEhjCOkAVV5xns/q62D9v80Yu9LkL7GOPStNaimH0
0fLZZNbLN9aXY+LXsOjLmXKIRD1NJHFD/6y4EmfJhRxv4wTaSxMi35TYjtTPOpBQ9f3kiGqvET6q
oTK12b3zP6bRyeM2ZbhHWjG88vLFxPuV0/g08KIWxnwsizoJce9xWIbPH46yn/atycdYeI6hNlt4
AsWLZjzzPTaNgwoNSmXe6Z/iHwOsFgDluZ4wunNLVxH5Ru3KpxGf9jGPoEfbj76tqe2kxC3Whmb2
TOD3EfgrtAPEX3iiwhkJ68FGwrBXobVCgJLrLQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AYk0GVXSV/oBWSOxjuGlD2oLlqIfBX5t16vozwXg1+siZJZSMUHEbzptzgNoTGyAuDaMihDY3BLO
EtrWbX/36HzF6OYvwf5POdt/VXMiD/WmbkoqBGEm8hBrg/s//Xc8uwTP0aCjxNObZuBko/Q25mgQ
30NgIumW8FqCkhPd5zaKXjVEqWRkZbVy3s9drUMCg7SmsRWiURkSk2U7gJHgxqNeqEvn/U3HMsD5
przVbreKAnJv/RzsnAueSJ7se+zz3ea7TcdOm8FG4lJPtFHb6jvhIcFQ6qftny2xQ/73EGrSBx8k
emkzKeZp3UgSKQV+dZEMJkjg6+hPhExCSG3ddw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z2aYnMPHx9JY2YhtHwU80KMSOWZwPC6TzLQf1GQQ4Vnr361DuLoPMu0MbOnkBR90QGDH/qF7P5Cr
Ly2yiYO0/eJzmgzCpSyJ27rzee68zFBRRDPmlOAN8FHZvnbWm8t3N4kjdk2vzG0NcvKGeDmWVBg8
WX1YKAu49GjIv50pk7s=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZhLzhPI8pgMrQMSYddC1+njODiKwQHec1wBB4U5W8/l4gRoB3jhisEMfFb5EoL+ePeazVA8YvpBO
fy15vYUdxOsCKx+vVBouvB0iJLQJ7MJ2yB0Atezf8W/dnulTtecMT4xYThtmLmUoLpjc/XY+sv5+
kYuBtkUrJcr6xJNsQtV8JIkAU/9rh0McphkltAYVfKvFQQ4iPL6Vn52nStdWLo/EzZRGxkA2w3hx
RxGGI0fCa662AzFgfo3+9jW4FVA/MfRfrEnMa/qSzvX29NQHmhsMx87TbESpFUhf8rcOf4pNxnvZ
Kz+Rm+SekS5sOFDAnkaGJ2fOU9v6YhYC3w3/eA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
pWAKVmJWCll9whDRGM5qzSVQzapQvLsSsmM1Cnq4dra+fhdRitw0chHMW7E8oUAr+TSzo3swntOo
8zfLTIRDOv0f0KCF+GN/J0vVglj02cs2vexAs+zp1YKKsHgd6xxD+xpGwVYv33pzMvyNQXmwPQbo
vLminacbx0eFJt4KQ3LKfe9Ce8DEQqL3d/AdV3k4A7nwLQsdI45dwXkwOaPOrKlJjz0iBvFgzxAE
9sOpDEIJKf7/ePVG+rKbhhZrIvX6HFoFaB5MCrmfqAooRAHKUZ2qCqjZmvO4JXG3LUxSVxYBprMn
vMSIM614WN8oIvBB4Fy/p6gK5MYKadUyPvl844R6DNeJ5FxHenzLlgKeOr/8s9672MfKJao2j87p
QbMBLyytKdtzM+N25RHaHPLM+XwvdAmPjXuxdSU4ryDOjJ310sQTAlhakb4gKS9YcGID4aWXaX2Y
RhMxWEoblXVBRUNkXWsH2KSGW/3hfxkR1yYJ93TEsbEYEGlOuY6uvuhBRZGvIGfQvGSxcZwbfOpk
6LodibnaFkm8damfLoRyEony4TVYchMsGArRRRSHFBYTuTFOhU+EKpAqByTwvgcpYe600SAQ1pDI
o53evw6oGJhy4Knhe+Na3ncoRYRl2c7tvb110McW3KvDb+TlCgYsGBEx55JAk6bO92mhWE8ysviN
XUpY8pGd5XPlUBUm+BAQO5Qa4KTxI6x0SsJHK2ok++e1GjCr7ByQ79/8Vv6g2JXs4CaoHADtIl6G
9bYAwd+e0Cc0lcYbIvxAdKNRa63he9ArMXbPXTObUkwqNbe2z4dFYDjhiiEsoalLJgY+Ia7dP3oB
0I1RerqoRLNORICAqtAMSy7FmOEUYGulapMCnmsTAdPSdw9A6GiKN+EwNh/hwk2ufNew8m7uOOGT
y3NhF9bkkqzCsbIXY34rHpBVRDz7s0kNFUgVYw4KqcFb4hBJwzZgToyqQEUkWU3qcPAvgPtzSdMv
FxDtm8wVOHRR8exF4p2D4B7qnPUqsM1ujGAwadjrM6NJKshnQ/r+SHuogf/dpwg+vQixuqwrDCgJ
t6Ui2BdrcQes3hNPXj/2zvHT8sU31egzEoIvHJoay5Kjl+MrYednShMzmj2K6Xgeb2/d0ei4YJv9
Nf2aa2DkEqdKihAVrnSlXMGeSNLbLTRf1Xmfx2SdkKvl0kjorgIN8aP+3tSvnLhbHwsaeNnv/27K
GMFOqX5msB7VtqFqhoDKPmmhYod2GtKJ2QYX+XDu+79kk5LDXxnv7NqaCv43OS78hkBXSUIdaGif
FP9ZHZN5Fr/bJgIEXbl+gtFN2no2Nxdpl/xkRiY8EBGLfTDU3wXtBG4eDRzFht24Hyi9f3pEqN6q
KWjjsM15Kn3P5ow0oT0L7A0Q17GWWaWlClM9i/5vYfBE5vDsWEalpiU9oOft00qM8DEZkmL/FHpR
uhhVuTzGgKuNexXpxmidxBdjfqesW3W3J8hcwleRLh+MA9KAq8vw2O4h1W2jhbLk7waWB+nSjQrC
MqVXdrnAh6grQat6lhGzPQPos7EX+STGB7oLpPaVghhM3OzCHcX2PJfBJARVY183uiUNAjb2lY+p
emHvMuYh5lPDNGx0eJWl2J8mT6/DSDFhwEPWdwNBeIDHfsWtWbSqhRJ5aBVxTw/p+8ml655xOZBu
77v02p/CFimsfIhBojjEZu2aD+xSW3wJSWJnXpvZXfqfhoHjrXYvA9JmyU1nsXGH3yovWIlzKY+7
lFDi4HHhcgLxN9Fxw45vKbOVFeASPweTUdX4IYRdn7+h+A6uFFE7hxXWUZTo/VKYW3ZepzaKy9cz
nUetU6NV+0ZgamhaCMb7OuT6i01zajBtbAh2T3YZ2xFOqUSGUXE4aElYocUbwGBNGqpMU3q108Gd
lujbElK8q4OB+LK7m0l7rabzyQgsBrzlhDU49TgSCLGcVNlv43ULMjbT1ws6zd/4jM/37LhWZrgJ
L1QAOC+KGWuPQD98GD/brCZEqHJVk1pA7pgOBMrDNtpBXRmX+VuKrkyYlq3maJ2sOyhGmuHQE7nn
Nm+6rW+x6S+4HwZgfu7EGdJ+WLdIcNjjCL3BnpNnAVibxmcFc6Fa+MT63vsI+M7dzkoCJcnZe6WX
1bSYiB4z67IqkZfacIJs+rKhcCDv/dy9gwdwj1OuLdV5SAGQGAhpWFMD/CSZayhKIWjUD1TnKhHo
be3nmoofYl/MfBYgZvpWtSWnhT9XeBPFHwV94p0epy19Yj9FW/I4g3r0YTaz7TFx0O0lHRY3wXMp
vkZ0rY41Zf4j9cUAUim036OCSCs9Km5eimNpzLw1yVdeQW8kJQsQU7z59Znz2otfsFjwPTTQlKmS
3mFtMTcIovjwMDjYxUCPPY0dEMTofEGQiN+XO4i2SDNAvpo/psCaN4YDT840UHVGylMvglg5vSeJ
UHPAtjfJd+cb4hPDeI6bp3OFrqfi70O03+xW0AbAoYDE9evsYM4irxnB7o5qbKcHBkqR0jFTE1kH
DR7XBQRUIKqG9zmXKqFhvMqicRzaIskXNJc5Go3yOh8R6PGxXDZkJ+BamoICAn2aR+E1VIUuW1/9
KpQ5lbkZK2j2n5saFsQ3Ese/PhO4rp97qW+Ls8zyhxrg5zcq7sb/AZ/MIxmMEr00uSmJP8DHXAZn
Jznd3e3tCV5xQVvuO0FSwp182CB9mo9LkM5mICDdpPG3aw3UvmSSFm+k0wZ5Vbm1iIa7y8ayNivR
AAtFI808Pa55EwBQixm0ZGpaNkR6xzdRDCDySImN8Nuk99hBA5bCbuYOBQJPT4SEe3jDTdzpzOS6
vJNrH/CcLBYk8668tRMYoWNkGNuQ4ip+Oj87qYiKQVD+LK3GnuEcpptQ1orfJXunbl9kwET2L+V3
zeMB6CZXsaYD167B8Ll2+SEwToWA6xKvblY3VfHq5OMJAXuavuAIDGkzuo6ucxQOnbaNRpTCSowT
gPEB3SaIVzHP0AAmtO+/CgnPY2c+EJLUN1s6GyJuyVH95VbdmTsgM7c82fhf7cw6dgfT+hVcJvgE
XKflxbwfEw8Nru0eWRBnO2nbtT3gl2Ju/2uAXgMcoRs3v4tZOwpz0+FhOqiNUi8K+habxltNJ7bl
uUJJxlklt/YG2cd3kFuf2jIio/mcKCHwhItAYyjdH49IOsSr87XfGUHQyl69LjvELj1ST7uT14q1
Bw+j65JiOc2fUfKArFCmr/qEgOVNBbBIa+K6ukEZHDCpyAN1S5cbU2gaO5fZWTrKdbxoKTP7iFzb
29b89Hl1BhbqiNsz2K54AQjaxoIIm6EOfOqXzd8eCfv7dhM/qQmcipChKU7Dxf3vYznWdrz18aB7
xGDpFXokc4ZnQ86tjlUa4rbinH4ck6H/3eQaMVhptMu4n8d4KJRNyTtYnfCgGeCi1vL1i1DfGa3f
pHRVG252QMcXykwV4NZ01nB7vrZHZ7YPcgWtiqq5RfNafxrdYMEGDjVBePvMOg9Nn092ZrDPjADS
MTlf2dmvXHM+RlwU4bdLxAIDFAJF3809bb+xrzCpJ6TNPSYHP6UpLZPnCBF/sH+V020Q0vne3gzQ
7bA4ic14934v04hGxq6DgsN0Zsfd6yDkTK995PDd9a0YU4cAF+c6gW7ToXmj3TBAwZ0DdzovWF3i
WWAezvj9UxEAYvAT0jTdJGQFXPJqXgN1oe2sQEsAClVhGpPT8A45Lf267LfM5f1ng6TMb7loe1cT
SJqfHXN7lcYv4N6soBp7iXji5O9TGtD1w1sO3sLIEWoydzb1FsFTK/sZSvO6bcgJ3vc3uN+5maUZ
20t4/OQjGGrb6aF+IPFVSOkMhwGbHAG0AeZH14/NDzAxDi9Cl0hfjF/lTzDHZPRwrmFFmVRY4O07
V9nmBpB/SmqnLmzokfU+z4bFd5ij9rbq+shGECjwOninaZzLBJlXiRuwaQsQQPnRlXD2FFGol9/k
6y5qTUnPHMv06dW/guTLN7rXYBtxyUMlUOwnAREHk59UqKkKueU/9lK+rAku+9ajhYXpSx67gPtJ
9zMK0BqEZUjWksw0aHHiSEzln3tXdZKEfB4ENB6Qors9Gjs1ATBokhROpd7veLB7YV0lEMY5BOy2
MKg1tQI75soojdO2nYVgFSk2EDYh5qAHDH5LC32xBtb2Px2yDi0jd4s8UB6eS52ApygDomUen4PF
wPluJomHmtHy6odybaLEyRn2YYkEL+pzAfj4aRwBhbOpzmk9vasFtI0XJUWN8a9L2eKud25ZvQeU
AsYTfkkkvAvSEzH4s9aAePxktN806SZMOSjVs3Udy3kJRCzTw/ZpXf2fwWoFNYqVSdUyx/0cjx8T
vZ9z0ZkLwXUnjXOGcGTHSFAruMA/7BdcF4fn5uPFlX/RgOcg/hkkVlufVSdd8PsTFLn5hApZB/tL
bHW3hjXrmjeBa9/fSrDYwdeLq/zg+TUh91pMj5mBfBZZ8YQDM4tUvXRAqeDb/auP4OlrWcaU/lby
0gV2n6MdhyLpt8zZGjGUIk5eg/SgXcvkFKBIPj2mznZ1RW9AhDAydOZ+v5SQDOrjPTgUpOGdtZOd
Wl/luJ8SX8RYTgc4Cte0dtOfpuuJzREPY9/J7nQH6aOTaPrx+zjqETHbCd+ZYJlSak/FjPupl4nN
RZJ117K8WaXYwIXewFL5MLWAiadM/yagxaGKcnfxXA236HsZDO0H96myoAKquZRs4T1TVxpGg0UD
raLqmM42Z6xZGzTDNpNUSGdfVEtedDx9iJh2vhBiCEG+iIT3PfU+kAFFvMIiXT+kh31vsAHjdHq5
blh8XAEUho7K4UfUHFJXJ+oIjvZOUbZIWJitwqxOvd48ebEjT3nFWTnaDiN6dJnrokJIyIeXOhGc
w9Foo43kO2ixVfdvQo6oKKjy1GMmzhKEwj/+TdKFgH5xYGRizQE9oSlIAptrBJI4yPoIw3m0yaSC
dUwmrYtWq365qVieNEMMiJVQBojV9lBHO1iTBTwphjZuF3max82Cnhdznq8bq0VVwJ2B3dr8dXQN
fNtuB9nmztEPrPNd6X2B6YuNxnsUsy6oIhlm/awxFAv0jnGQhNduQ0aZELHsYGcvS2CdVLCHFsyF
TLRVl9dzjvNqZrtk1o36PAsOAFPfvx1pRoIlw1XOQE/B/fGIO2ENf4Ktp1wenISObzuATFX5Wfzv
XfBBxwXGEszXWnPhUYLwY4NioBuTmn1ktTxSlDWflOp9x34isLuA7o/9fg4yqXhFGumN8vhUueoQ
zKURAmY09ZuZWwXrqJco1O/TynLb3aZREFh15njfgj+PWuNU28ddmX4biV/k0rYv1O4+EPbxNSPt
Eka9N2VxhVUDyza1vNoTihcn5Vx2GS0gAtiji6hRUs/pX+sP/jzlbVbc1iun1GWQmA8tmwGUCPx4
sPMaxoDwDH2DvBVrous60oI8KQWZo2yx12L2pJRAVaHMHdKWPgEDmi4Fz3WdoaWFa8rIJzTryK/j
7njaX3BCMDmW8of0RlKONjiGGpBmz5vLnOmt4Yd7guMO1oVezdDUczAb0pNrKJmBNLK7BRJPW+kk
gXSlcJQg5WMLOBgo7jsNeJZmHgoXW6XEuf445qPKlvKwgbtuHMeHTFJTmbk78E03dhuT0tTcDuM4
4GNbIM0hrOZlz5DJYIY69bejlhWRttHfFD0n8t4CkLON21rlC66Av7MCaHQj5pR5LIAkwAtj+PEY
6RZ/ZLDHWWv3cbCvxJqGoxWLzchzg+AxJrHD9hxbIKppQSy+bVtNXHO98GZaBONQZ/zJ+gZD7wEM
pJBaA75nE8nZP1dvEXbHpIBfH7JHQKJ7UWQJ3YOhcb5wH/T7wMe/djK5K0BEy/3NbM/lzDo/x2QF
c5dnMoXhWB0TDEw9ei4vQMGzRQkggwHFNGffuskyB1KSYAQDQK4DxSx53709/T0FdcmwaexrI5XX
Ejw5jofLqHKMZxA4+Ujf/T/cxefnWrFDwJhAFi4cYxJMSdniiEcIiql5oNN6GKi60jZ6D5uBkO79
3sd/XEkjXSEdcI46G5yYrRV9aoi5GUSvlxw6tr9CS/wTzTh4W5/vQwdFTBQrbnOinOoTXAmw25B0
KxGU6Uuh33jOvbURLkp24vTlMQvwRtv4O9NQHpzz/ZZRPsELA8aL7RaSK4LjcGWfzGJo4QBQI6N3
94lLmHZwHzJinoDhY7IgZtTCjsTBKp+o80n30z/Nzd6G+OCCPIn204+N0yib4iOZoP706HuY4Yq7
AlaHk9DnBW91lvuSLQHOjj1h5hhkVVhPdFbl4fWuhVvI2g2fkpNDneH+3y0dkU9jCYrWcu5oi3kt
2ncZ4VA2Gn4CdDwozhS9u+BWBfOLXRy9cAHektFN8SI4Lni5uiAFfOzwVWTVOENrZhy+udUYwKXf
yb5rbm1MUvkPFlWdKtNa7N5QNyDjvJg76NpBS1xdDtDBmYrO2hNOznBQce5X9AfJsZaEq+mnBVnQ
AsO+6S/JwnbqK+9POi035/B93X1L+f+fHu9GyOKRuEXuaa1J3Gsy2O51osd9AH5koZJRXUFwpJ5k
i1M4K759Om+RG7/+pvej/hZMQ82LASW5EP4ltGKujB04E1sA0byjli0idKHQ6E1D5jAarUuMXvOS
wL059uaQRzkV7UPuY+pnSGMgBIOTQUCATI+Qdf7ThB/p4o5TrLuxcq3FWl22O4eM8UYOOIPMNu7E
fdCRNNQe7r5fSI/xAnAX3wm7OkUDs6crSEWgmANAdGGJMLT9yhJpHc383Da+ZFeLfJlAjBVOg03j
l6HImDaYXlrE1UdYsV6B7/lwerN3z20ZIzyUNoIR7gaUxe+cCIaihtPHUGcooNBrPVAA1sDSVa1X
SkJg2iFcc4e4C5JcnrQ/TucCkEadkvrRrONseauA6zl/laAy2aNrCcAbsieDTEjRFrnysTKaxhtt
93cIUXubGD7CuxS4q/zx76vADKVjUUrTRJabr+OVMmyir2zfhhSnLpbQ2CQrGymdQGt2NfM3mSro
9wjmrSNy4J/Ql5bAFco/NegDsvPF8CSEUCJXlxW8Ka+A9yd7wd6esrcfCZxxs9nCszUgd+1OcKrP
oLTfo065B55GBX3NTdFU8GAKF4N+UmWoOSK+tZUTWSYgBRCnvDZGEo2OW+O6AR7qsCRtHcx9hAbr
ZroaSWMiJZACUOVD4LoCA5R7cX6d50ISjH8W04+CkiQkbEiuMaEXmfYDQLicvS9ZaTkwR7vH+vv5
8JAZdHlBs6gHJejLF/m1ZwCGm/tM4UYjzX2twmRQuypI8rmSer4JFiAx4jphnOHjJBXnXBC/MCjR
1oY8+e2l3fQJy8r28+V6To1N9dOy74BZMI9kBFeTVh1F6tFgaPyoo4H7pqupjlaKh8+HxczfwmAi
SJCRl8aiZ79M5Wy4S1iCrpkUkBR+v2wwpsLwRtTxZWCfhXSTal/3lpLbtgKljYQWw0vSaWpAdUh8
acQFbmijl0+PrrGSY1+hbSZPn7GeZGOeq4jTJ5Yxqe0OGXr3g6yfxoGPq/6L2uOKcHLDpm4gAUvd
hAJmQypiMfVVCeiCCIP8FPmaE089kgn26jI6aklXxe03i9cUi/P1IAAI76hgYTBvMtLdwciORRzs
6oPNnXJZAonu7fCohFq8dvOLmiIqE5/ZvWBJ1QA5uQDsgxYOh7EPZ4zoo5/c6ioxUIBnBL1n2CGf
biNLjFA4Vh8H7TTZChTCRlJvCcxeKZKtoRcav/6PP57mG71Ggcbc1OIjvvcglh2kB95VXt2HwpUE
goYvrwuRTO1CbIEyqpHWtunMni9kA/mqG8G8eIRh/x3MhpZA2fC2a8AKK9BffgYu/+J47+qvA3fn
ZcyytbLsDrE1UMtvfJY1YEgNsH3Kkod4LZlO8BbMJBa4TfBiJfRh2uk54CYRx8MFgER/uc+y5kC5
UqdlGH0F9v/hKaM/lJIPm6xNWaDCtcGDAV0qDoVFCqsB/Gxo/fdpMjajweANtZLIxdH++DyS3rrG
330iDO+zvjwfkkILKVUTYsFg3yFM1lJwplgnDsJ2u755WDs+71YGQ05QtWyIdg17AgVHJSUWEFjv
9GPLTEl2Ywf0G+KI8U6wkevapF+Zwkt7ds3OzCo6TKdwwjSoo/3V9YNaHw1qpeBKsnNvo2z5I2I2
znP3xA8PcdbJB4pCjg5wBepaNY6DjP5W0V2S2mTs9WWw0NDrlDIhqZSfrRxRwiDvvk7ee3jRGMqJ
vwMppn1GuY7UpWbRprvLrFge7glqClKJHErElqRUUCtfsTi1u+8bZtKciajLOo2pC4JfPTMm0GGp
Hcbhmto5xQvVxEoWqF6I9+UYNQhg+lGGehSj8kAt8SrnaMX9Teh1hn1X9HWHTFmcdRv5wigGWuht
H+mpEGHADLDHw/dLunOA6hcEP4AhIP/YNznhihJvCvPfK5JCKLlaP1LoeCKoevyPHAi70RvPdVGm
IsYxesa1GHnUIY8e+Wk9YPCZ/u7fcI1YK+PpIcCDgQsVt/2tcr3uFFt5lCB7VnPNcjPyy5JSKhg8
IR6OMm8oqJxx/RJkltRrTKkvSnpIQk2AnnYQHrhbx8PXzwUPOiTDrPciTHFVNoqqKICsCneboRkr
3ddwnofbZc2OAszi9CqIitcfyy1uELtWpY8QZYBDmuhhJkwAagMcwsCu9HIW1iglC7Ouz8zGa+wo
w6zqHdfB3JREGCl1tRV3JKaU7OftDKopsa6+PhyEODuJYnG++UsrzAefB+d8xslu4nMTx1mTc6Np
3+8s9dAGQxVcBLBa7ZrJo0QQwJWZJvqUobIlUisdpOcBACVb6P2UiNSRpoB5FJhoU09/+IEyL0io
nlipi1aJs0w3G4k1Oo7JvYIvgt+Vlto/UynR30L1M6is3vnrLNwlMVboVYo0VRwQ9q9sCf8aejvd
Z/FACsFzeoGKwx9n2us+sx0CChgoZ2AqJxL/uydBzeb6gQPSetCfGswLk6jjU9twrpwgQ4UZPxfz
4LpUxQENs65WIA0zzAncqpzSpxtzC0bwhftpHYbmY5ux19EuoYVJzQiHHnsacB+y/cd1MTo1ckT2
8OvDa/Ac80kZhLz3yhVCZkG84UwZmVrnfBDU0cHD+gddH0uY4ZnIsJIzu/0VRtNPz7gUe7atev2n
G3/sqwX2OEITIrH081zuH8iXSHAE+yOlD955zKZQY5x663GfSe8HdJ+zBNg2UAh/CLDAscKh1LD5
ILLfCC8n5/7RGGagAfiUKn7vsNtXNF3KKoA41OUtgAIR9LlPKyjRhPpGBbn4LFaTgxFOv6QuZc6D
yCAvqWinm/EF/1wXQdh8g1ICjaKBi8JG1Y+WDUIOXGXf0lwKn/ufiygKttjK1bZ3RRF+34cM0jOl
WwalTD+TrVU/qrF/qNrJUWq8oY8kahUA0mdblHatAZBkwhfltsos/Ugv9KFYWMO6wCDhVLusZb2v
Y5d1W5/8LdL5gw7nsNiqonlz1Lzm3qzGw0PNOq2GD3Cq/N/CXfOLlCnLfgRnjKkC3NB9TChiTFht
gb7gdRg+/A4ldV8br8Y6XSIZ/ex7bIL6Bq0fBltO8XEMa/zazJij1mKVDcyXp9hTggfSxvy5713X
aAf05JBMMN5qDtDagqYdNTiZh4SzR5UhwLWNUaq1WU27vJGjq0DPtakfuFEp5L3gx0xuDJhx4PoI
q/Q9iRkT4NoisEswfo2c2I5e5yfEz2R4wqqM2DpJjqiCFXBYjrSVHT/Vu8T/piSzaimGaa/HdK7L
A1NtLieDEgX1DIM22eT8Svl0q4GkahTTuh286/MggMriZMZ/SUaM/GD4n9QUq31cMKputsuF2gNT
Vk0dnyX3g8LxVMsVny/hNAC2mxNtMsffbMNUyRvkbLNKCsFJfD6Op4v8JA8jDsenPPlVPzkgYzw5
yA+9wFIX9w8zLfi2yzkG6Yq6BODKfrz1VKMzptjKQr2T4HqbRWiApS5UbY+WPHFJ6W13Y6jN6/IQ
ZpbcScardYFE2u2wMlznftn2OwZrnyJa5TrX7Nm/deOyogmDLZpqnYQLSd48KuMAYioy/Qe2MHT2
W5KT4QGTSEn0e0oZh0++OT8FCG4LQCf89PI1WbeVJqmhOvJ5NhkoO+8dOWstU9/7YBvOPoQyCyOz
0ADCHjbXUyXndZzQNAbQmJGSBZJTHYU46qOGC5viNgnKGRYCfz/P11QlS/2tA4zcwJPufHGLnMDJ
Rbgs5Ci5GfXywZbVDvj7MqvFYGfjd1o6mCnHnN8iJe82QwzMGAjEgzNM+3c9sYGFwxbrJhLZ8O3d
RS6+qYe0fPx+QT435ml9GUoBQ+0MJPK+4wso1pzmgcntV/PI24SjRxExT2ny3bSVlNXnpXKwldrA
eM3okMLaz/oldCL/tJkXtXRoPkehtcBdYsgF6uR3dn4ITZ2bp+MhISj/5sKNBKQuKLsJY3sZn19k
GRIiIIRaiVSj1fI8l7uurwNMCHpM2LJzBpNfndxE8bBezcAwxnfF+IW6esuLGWYPjPJlAoXCz1FP
b/mcwKV7G4cC+/7iAWQmsYgt0uoBLV1F6WqMnX7Mk85yiO7Tfq0RAB4aAVLXZP+kNO5QV5+LC/Uz
PqyGszJfgrOcmTIFioZjkls200wQXeT3py/NSh0K5sqpJwsPWfIsBUNV67ZIkmuofhfEF7ZcHdJD
AeWFTNrwWQie0AjcKCLc90G7B75r65GwhkL7P7O5yyzhZciaASoqpGbedYA6HBvuIV6gpijpeh2w
Lfh0xgbI7vJbxeYo4Iyow6kmxM9ut8uwMfcZfNaKTZYZ62z3/fuEgsG4a+acSu6gCV4CGekQR1Ve
OMWK//pLX6Q0kjyd8JUZO2chHMiaZxKoY7ZJeMOODuAB6cT+M+ykPyh366Zo1Rmpw3vUHUFX8mP5
kr1OFyLBrk6ek6KU9mAKRyFNxnWGJg/ciQ3xosUS9nKSR+AVj2vHLYwytjqTeN5d/u3aljM40QEB
OFbN1mZvcU0Wy9yUqz/+uN+lHwjuiJo8fGblz7rWqIhS3RIAIY63Ufp62G+n42fNoZrXbE+wgraN
sbv1Mc5+GDWU38iBXCnvCd0Nb5xIJZNbMqhjZWAP84/p9xkvEKRO5bVMkG7CTINyPlLyCs0rqDPl
60i+tYIzcf6m98el6okDmuUzc+l5SdXQVAHVLgHHUgga7r2uHj7ap/5f2Z1MbSDO0Q8cMOdfMb2T
/VOZzd/RpUuGh5L2xucsILPHLMGWpsujeolpsXpVBILZztoaD/GRWTPydCy0zhJL9fdDA3TxPbEd
dpP8KwtYxrzQLItZ3+bf6fnofU05l4Ojk45cYdhJKUNc526WlmxWqggoh8zQgRVQGsX1Ye+Cpq2c
qu8uURAqpjTIq30mjxDhuXKW6faym0WDIShOa9jUHzAdueFPuDUwNYZCKe/7SN+megGQ8Q/f4FKA
oCqBIbfqcvKSHLTqQkoRTBLrn8Aafpl52WmoaDA6DtSHcqgyDxW0d8xUfKFUVQjXBVw+o3cGRh00
WzPDGlfhr55KVxilSV7frWY6qustsqAxNEL6l8lKFro1Ou1CkRjHDjr1jNxoOEeYNDmePsXo8xvX
+F5uHs3oaKbHZ0V9MJ2pnP+83dw3QU11p417iznQ5yeRst5WW2qo8pNNACq22V/AauN/xX6RYDup
D5Xjbx2xwRqgOy21z6h6Ejfhy0mJNBVaj8SnLZgTUtq8tkzKE2x0bPlTYGvHVBmF7dfiWdqYKSNo
ikeSqpHhefUFZ0VVO1ZMehhkErIdKMPzGkUf6S22t70WQiOEvxJWk7AfCcYfaKlrHlqtC7zlthyz
tFw1SIlhIXQgk8deMDg/LDJ8LwFGuDmjevPgA+OXpo3OyFIT6g+vPrkH/RHxY/T7cmDDZYkW5j4L
DEzYfxylL5lbp7zdCFyNYW9H5zQoGEMaDn9KoL4/c0HGm/k2r5bIISzWtPf1OV1BxweHzzESDPMj
Nj2OnDoSv1W0twpunQa8dgqPFDIDM/3Fyzy8/nHsp4HfG9RXQvXUbAlgLNTItMCHNwOMGPu+Arj+
p+mUKR/YxY6VNwgEi+p75Q38EacN19rISDytpt9hcGMMCHJxZRdZ8YZN3y8FIsAUV/3Qmqaqfur3
NRH28qeUhKpTCDvVkqnmZrDZdzyprXJqPIT3SZMgrR6DSmS38Jf0qgOeftiKeMA2gtp0jWeoiaOA
tjjGekKyIsRqB7nLdFjgOsV7MhSgZqwt6mUCbd55/ABopACjfxFxWasLpdCSIeA6eMWpmjM6Ganh
YoeZ1QVib2GmnrYsgO50zxYuP5zTMNRuTFgb6Ei9Bl02OZQ/YKuDEhUTqXlXizJ/lEgNIkb3KZb4
JgBpsYJT7zo3Edwo5dp6dqAFYbAOx7JKHajDNf0yzN7KD98KNm1TsCkfMHMNRES8ZxKuoRniez7E
X1qOlb1YaGeqMZCiuHddkEkUpoAaEwsBr82jDQV+QpyNdy7hoqR4GGiUmAWbiy1T89wxL4U0qUDC
LKmZpeAIFQ6HzHmlGVKXHDmrJ5+etQN7uTh4a34827kNOpQz2kiZP6QweoS0vt35qkowgNfSy3/T
fOYBETiPsTyPmuuTvPXfxKzSCcPBlPqU3YqqLnwCgiimTwVJlyUl/4bipqL62JjPAKfNxLKxIli4
hAPD480ogt3pTF/5aDaDZ5/Fay31ooCg+Zi9Rkgq2fOLB8TosHtKCobRSM3m8XBhOqWZeSLuXGSv
Y0gjuZyKCDfQ60aaV6B6xkWxjJa2gSYgUYMgOIxbK/rkuKyOBGxTQhDR4iAseaMaOxYJaBT8Xw4J
G3Iwt2tv0tyO68tajKdqvtflfOY0MnQuH380msgeuO5sSVqAcRTZpT/xd6zBrrX1AJ2dEkMSm9hi
KO857/RH8MZM+8VcghQZ5IUuO1eRNXrZmr41h4AxyWolF6Weavmve38bXaaFejx6qKtJNV8sLT7b
gLnUPtmQD5cRAKdNWlk05HNfwxrLPJV9zIevHhgo2pexIHX7rGMT5cH1oBq12z8rjmo4zdOX08CP
JABQgRfa4t0m7fgDzB04GXUtv+1I0+hoDQDLUMcPGR2xXtkVFS+RjZy4kiWf/kTwigfOCMxnEdqg
foyR6pzmwDkt4DY0uYUBsUqdsc/FbCR3Gimb0yfSmB+jMKCKXXBgPC065ZLb8Od58m1fNjatJ3Sq
zRvy5uoJdMbGadPW5qQMvgi0684di2oA7qyEJsvRgANmSC0yyKHqBUqtsc6P5a4U9bF2IOUrPFO5
oL49O+NEHu7Xn0XTuSVFQ9bN4PKFuXuxH4Ghqej6fd4aK1nJQmbfZBTktfKsooMbttPgQqi8gOJL
y4DuiKmRyUbMakcFhhrm0poGpih87gpwmpdUiMJ8D/qpa/4F6YiSFkGHmKJF8bAV75h3MVj2s5p/
OKLT0k/rO6PQp2VC1+4JeEutod+cZ2meWOyBWVp2k+vrnmTRCy0kLTLqzu2rGSicCVbrmLJJOj2U
tgpHsc7s1kIFA/yinsADD+AsrQpBZAqgR7dF9RP8Sh93CTWa6Cdn5p+CNlYeSL0TfXz8Qbr0kAvf
Fmio4Sno+5pBc2bOONZhlYS2pqbJho4pYUNo7J2CyB/YsRNGfD1owy9s4aLO6VklpgZFz0vosB2U
4NVjVnLxwHsIa3Lzx4tn8+T3lEgfIS/n4SiWTG4TxN3u9WLwC1K7zroYMBtpZt6iRbFxO4+aCcFY
JhWXM9+2sxCq+8MKdQenl+SwWCprIUgB6IftH8y8RF5iXbRi5xOIy26iezL0Vx85pz8KYF6L8cCj
Nj+jPqg12mndazpavEJpjvboqZHxl/P1HPJ2+6wOAVAomRT8ZKkDXz3+wyJnxCFUZ93C4qijgIZz
sR4hzGsneGfqWQ0C/sDISp/8cLiRKfSzg2046GX1WfjUtUC/ca5DZot13hjCAqFs2mFTXlsCPo5w
FwXnucC338OYsLLGmCbzhzXDbwdAbpQznlsgIK0UBjmNwu27UKkNkB2q33ScOjWiwGpLVEymRi9r
tsxVxLfIOvkZP3jI7a74GMPjlSvtgprrfeMDF72Lnf8wqFX6HwstNjrPpYVTR2yOYNTaeqClZYk2
53A3VbCO5s/ras98KBkYpVowVOHwPNog73z/t41caRa3uQat6SpfqWOOy9JRT/ZrYqJZsIiSGswy
4Jq7Kccr8X6glhqSoqTirLDhqENl5rUrP8vfdmmOR633KS5nfPUvN7GhiPLap9uQbmBUn/HjIkTd
KxM4CYIIgKg70Usmz3E48wYk0oHQxhFSk5wqN5042MkC2d/GipGlxCpBT3sOeL6hQQyrn5hX4SEu
qU9DQZ3ba6dUixBvQEiNRJrjEqlxrB3Sb3mP2+XYzGLxNEUgbZjxTSSlVQVdoAXlayGpjHqR5XKc
yxKsMnr6FElDc/DSY7YoMdim2iqFfkaMIIMV/h6HC9ygNIMINilf9KFMW9BSIlXP+fWDBEXe8NA+
NE3J4Lk0vG4aCyrS6Dqn6o3Me4GMPWd3WmrtYtS9OG9qeYzFFzYVyam571PjtpGwD1j2rN+sutxf
YokOWEbUuJd8jdJpfz1IS8LUae4r8gH6/QeSW1gsJPWAa1a5uqz9sv4GmzVYOuumspqrHtsZLJdQ
Si8Hv1JIvurwIIIa1C+RxBbMrHav6OFcxkbrvbAE9mQt0Gt2/FV9KomhuGDzSnqZaH/a4pjcWLdx
ZQj5j7anF/0q5SLwQzJkz8VR/4JCTLIZzG3hJlH48bb5Tk4OEVVd90nCsejiTU/vdJNUzLX5Fsbf
vOzYcXdWAwlOd4ocwfsJfZswArYAOjkMkNLHV4Lnl/6/3s6cVjBi3x2aqysoX/worS4/sFilEDzT
F/CJyPkHC5L6BXI9/kLLGAusVtMGG09+THnTUMLsuY1/4WEOTkOwjAVUUTpP6cHQzRF6sZXcKs4e
aYJTNzFPKhnZLBtfMAXfI/E7gNkaqk2Lco9FP78ATYMZf5qVJ0A6VNNvf771fP3vTFuw0cXtvN7l
v6zWpx8ihhWLkOtDG5J3kwD80brPsgjaNe+ZyqGiOotqg7f7ca2D88tzin11QqVodbLt/i8f6LFx
0DmwxNiqSe158qb2j49+zdYOtHwxUxikg2VPXX2WYs5QmUA8OQ3O17tROyaFIJHCS5+L11G3Lfy9
iDebtdBW4JQ+YKk5rs6hqA5tp1K6NUQFZhDfhCgLc2YCs/H57RNqTqO3OOkmK/xZu6kpa3Xaya7h
9ZJgXo79eFy+5U/Hz/3wyzSmGgMPEF3vlUpWfqoeSkQnQtQgTznoVOqn+Zo1vvcHzRdBPvVsAk8l
XABojGz+cRG6dXpVvws/MLdXCrSrBvqOm3Bfy8+c/1bIqi/osR8wlPvSzzGrKQuLsiPU6Z67AvlV
Zu90y9ZYyvVjGCzZBmegc5KvEY/zl58CSgnRzFpz+qUgGDaHEyUjRFSh4z57xUUUVQV1kcPaiPZv
eD61yQyrkBuIY9JU0kCnUxk+eQJbyJZsttq9TVumv/XjUOD0dx+3n2sAPecPSCHh3aQpRAYOULHH
jb8hCUCqNhb6w6OWV35tHv0tQjScmim7Tif2RcQ7+ta/AtxFRE+8/Q9LYF/wjAwEHWKdoYB2w7Ws
gN7GDKJQPSE5PrTxyvwI2PmA6ZbclcPR62VazSQVcyorNUz6nd9II7iRsSSBXKgda1R8ynuBnnFh
sy9WQJddSfqWtejvQP0Dvg05NSOF6+qNbDn2mZUlZTQor9fSARGbgCrwbBj1IEQK3yUMzVrCIK1K
cDyfb54RhbpqN+SoXW4+92TNaAG7yagldijQnxm7+40MgxGoVJPlGF8EMlw1+70iyDdGll/6PiwY
m7Bf5BnCZ/XpUQ6TDpjIxbKny0Di1gGJsWP39yiPoAoCdN2fC2pVHiscRQqvqTlQJpcs4KPcVX6Z
FiCHF0oVfYpuZc7CjN+HIdCA54DSTrgIGtudMFp6z7yzg6gr3uLWBA0ef+jpfkVt49YmfPCVt91M
nYwIPgtJOUwpybPC+v9khJN4KiYeKmiVOI5l3NuwZzmRsrx+LQsy9k1xyx80Cd6KXlRpDgG2t/Fi
1XjoIEfjMYUWiUPVFDPtTVVk+CLKOWLT4J2HPfcWIeR8uMlxT73bpHjlMwsMSpJ77qfrkWdfWGSu
f6uyvGnRFwPfOlyba/Xb0fdYLwxmjHAf8MiB1Ze/gkKlq1vXxWQQnLB1w8BTRoKLHE49RXkgL5ri
+1KzvaEi4uPunyJQFQ8ZRfSPdYmV43IFNLeMDc+pbf3d4vglgSS/stejwJgBFGEWt7i6a14AL7RJ
Ud9wS6doypxZ1A/cvek5Q7Ws1HgHMJFVsx0ksQKzOtOFYYoV7P6LICz9rUjj7ZzM8ENQ7s0TYK7E
dS6tgJZ2P0vJfmHp1f3mxSUWdL/j2MiX9QAs1paCeBcHpQIQ/o01fFdudGykR9NfVLnOXhAt9NJW
5tAc5hhSWCpns+FF79GGukH7y43k6og16DE/PfZAKoxFYGk/RVE+wVn79wLkra93Xymo2IjPEm/a
crSNRsZf8KKGG0flzikyVCT8G+ywrWl0z4Nr9l/l6rHCzVXH9e2li8gS67QIh+PqXxCTXtftOIG7
jGfbDlduUDI8k6ynaDfNYltxLl7RM8HCmLsJ5aNjCJl9062IC6zHgzgW17fexgze+yl1IgnAJJqV
9qU7KX+BZDcZHxCe4xAMr8CRn4W71O2KlC6TcbCHzigT4BZevQcMTJE81uKj1H3dcWY1LCujbj7K
Pt28GDPyWEfT9YoFjpdGsSIG3df5TFuGhu8hr9LmCk1eTL2mdiM6B5W5u3dpRtCUEvi5l8xHV6hd
PJT2YtpkQktS2EPR1ymp3PI6IN2BsNC5W32Opq3qxosCL1doROkMHGHp9nZ9iPmDQdQKJEfW3Z+T
qMbDr+5g76TK7N8d19xR26O1GxupaDpAn3134nrQ+gZmWIgb/RN3LPneXpBgT29WSDgKTJWVP6b0
EwuYb9UNIXtYPsxMDEI98JkpdDkyhdW0E80LykPGIk88g8IfGySNOpAr2fLHewYOMDN6hWRTCM5I
v8oy8QvpABoZzposW/O73ZFXAcvBhozK38HR/eUhxWTlTdTUpmZifE1a/TB+0odP5fEZgjbP+UDf
HI7fbLCZ9jj6wW7ivG50P/YjjOG6zYrYFJBjD+VNRNUeKEulZV+spBp4Gf5nHuiYbK5l6KdDnGPE
bkUV33BMv9rigjJkPo7xJWoWpXH9bMsaXlr0v5hhk4bc5yUrgXSM6vryi1ER42yJb6u8QZYPhtmq
vqRHgP7poQJ9UNwGrcRc7ld0PkcooGRZsllSPakk6DulMfMj/v3mCMb4+H40blzPo3T7lDWlKqMe
NvHMaow95fzCy1tXnUG5oMl7aXl+wZlVb0YOgcKX1NyjT75Uo+tbcbQi4goGtnEd9VaC2qrxg0ZQ
iuvsEoDDLs4PMAvaag4A+SXl7UuSTY7/zqRoDlZb9mt46ryIBjzwDbVyhRL7mp7i4Q6hhv68Q9C0
Y1zb4mKVPZLwOUsJj0Qb9uD6L4zs1vRbhcCG8sbTnBn3qWUGUQmWSk4x6ZdyH/E2iE2re3nppGd/
DGDSYPO2zLSsBBdiRBZO4Cq9ZYBU6JXtdz2kCMijZU2rIDpoGlejxBXqAisnfAYUCqWybSWwiot8
0K4d5vEyIVEtQSfrSyPv1UoqaaTv0S3SrQBmB8jH4+aSrgniooUrTVw/m42xQTyKjokvGmCMvXTB
oFCBaWedWT322C3Gklhgtx9JRbW8ZX0BOdYxn5R+NWJ+s+Pz+cVqhOtNXcaWDkaOdTNsedH87PIg
5hnjmiPczPqUXwq7iKK4ognhc5x90tlc7zpH4nPZljfkzlHAMd2aClWKHJoZH2FwB8l8QnOMSwQ8
8BWSydjX29OUZFUnh0A+aqnaxdNDWY8lUecHutdz82LNfHfmeVAYamVbpjw/DlgBn6kpSN1hnkaT
gNa0JWod21dGCWbohB7QqfMCcwhXKUxeq2l+OlaYAyBKr1+OQAKy9OTvK5QCpTNv7tnjWIVzlESP
ki97qITgjmsYnYwzzHrjZ+JqNnRa0itMRTQJuqG+g/bPvJSuc4mjVs+umGLuxWjKcVXohSDArDnN
4S12RTCQjEjXjauDupEeKXPQWJC3I+5tdPdhH8BXFgTfWcJ3ROFCnz9HDo7w1aVypWPMMA99yRz3
eESW1WEnco1irIcC2T5Y/IzFKX2GEJqkAJL5rQmxrXP6TO9RRO3hovKoo5yN8ZqBdviOfZPqxHCq
QImLdI7d4OeB0eXztPymQlSLcZTP7V/quPT4rEYbWOTYTuZES+I4T3WhL6Lyfnb4pk9Jb4w3OhJc
X9ybQLWNfPth703nvCO5h3Po0YYIxRFTXIdfdKG2h/izsf3CtMxYEbhmgf91VlJZGvNA3SRrC8Ji
3lYToRNwXI+ITsrtio0ETgGvQDtz8W7DLLBRCNFHW7gXj3/h1TS7FsaZNtPRd+Iv3NGa1JnIzS4+
LKFg57fFPhUDWiWL2XL/kNCy8JZShVxhiI/xnzYeARrfIjWjsffMtAfrJ0WRQJZA/pEL00aA66Fx
aVyLudsz3gxTVZeI7YlTdI6TnlvkGFlBi5be8hGHE+aFtVBoAhKmBLjUMuuzeLLiO8DqsE/Li7kM
+b93QkUOUDbTUiUOerthyGhIpmxgV+GaUHesdPeL7YUcixWrkwnKy2BbjL09gs4gWipwoybcn3h7
DXqWxqrbRh2uVJDAAdvtec16gd/01axu/GsyKATaFjWYlh0Y4g1Ppgx9LBMZdKUGC/yDt0AZ0sci
kwkYEkSzTVizFSKpEF/0cUp0mxAOwemvkzGRqrMCiHawsnGj5x9IcnuRe+GSZyFwcrAy8K28d4lw
RE5iowUlHAyXZhpgJbmwtr5PvVCWaRMXtQYI8LtJmOK8f48zNWdEtI6ZIS71lk32/RJ16dDIpWpF
IgU2m0wBI23pBLEX8XOI7/b8rh6dvw6TAvd3v1aXZyfKaRfbKMHQfnphEb/GrtF/mJl7R+4dCA7h
LJHVBZyQBZ/bXQ6Oo7L/zoO9coxjhWpQVBAh3QjlIq0hfw92bKxbRwOS9Z7jCE9IW4eYW//f2ZaW
+SHKtO1TjMTz25Qte33KU0goPPc2KgzD4/9v93fZ24l1JwOCsVX7WqKmmFf/67nxSC+4Flw03i/l
jGtr+iy5lu2oKxHwxwxAJZLbPfMrZSBv36P97QTGGPNAyQ8Q9JAOeECuChLkT+ERgZXXDfuzQKo4
+cs2wvAfwSuyvSp+OJFyuAC4t8aijHo92sgskj6G2Rn3JPVA0AxpFGEIS46b4RFj2ndT/7l6hZyk
ii/AkPiQRy3ZIBU80TazOpBd9aOipC+lbSZeTR/ynHZNpLGXYFO/tLQvm0TRA7GXn8DaQ/Myyw86
m0jquYkw/RYx6LsyEyssmPVFC71qMFPhaMT0wWznjScaQQtUXQreHClr26qgCxXimBOrGiedawVZ
HLWLNqkpthXMPC0ABh1u8QJKXeyU1tAZS7opiBD3ksCr5GMDXAAwm4Q3FK3wHpUR3kHKXKXN7MAB
J5usgSmKiulEh1VNhN23KvtFarcO9ww/EMMj2Nt05rPw0Mt43jyeC1Nq/eEDHwSQgExow16pXpvt
8KhgoC5GeLWszUxLo/km4VBoRcta3e3Ku4JcMWr3/7+u5qOi5bjBNesTX9hOrfKZ1ZX7IKi7c22F
2C96o3v7egBHiCSzJYgHX0jXGd7thmxwT64Y5dlz+qc0Cgf4FHU13WINjvIKO/I+YHeXYX/nf8Lm
O5LatsZsFFPjE+BCP7vGxnZSTydKJr/Rg3LbrvI2gW8narr+3LOakLQ7/6y7qvSxg1uMzZYQiTnp
z3YRNplmcTVFrv3GVe+gi/78rRYWAsNJeHLwIGkRtQHhH/4BzIoRPGh91+ZuFUAkViUlJ6P7jPdz
KEggmIpn2zN2qR44d/9sKCnyxCYOFN8lLfZmr0ScE2unG4ie59IuLUKDGOMYnttGFrlU+mtWcHU7
paMlu91sHK/LlhdNMby2LWA9S9oZAm17TAo/nPHRIeVzPPnqf+oikyGg4JDK4Et0XStgRCe+kNLv
rOg/X4iB6vnH0LMy5c9SwCvqEsTRAdHr1bhdBzX4jagGhUPShBfPJxjd3hZdaublzLnHhnHxV6rJ
SRMTVVb4YvYQRk6ewc6ankWwdezkPfsLnq/i+DKdFKU+iy/0L1dQVUg7+6u1dxhOxJX5e28sEGiL
OxK2I4DCTOPodjp7UcxkcQUjFJr+sAWoaNmpnaUt+4N6/VjvD2WANcZEgK56RxbA9v+GW21zzxkb
Cf2ZS3OASO5ZPYGzSDhk2YWtWAfU23U0huiyQGnQe7Fa9CqkERipQZc1cszW05eQCmj2+KdfyF6R
ONi7g7/TjDwNWL1q5LoOZWkSlbFLjhQ1V35OqcBem1HWtnWqEYQDK4LMxvNVwPIFKMCcgGTAv1eh
g0zv9GCboe+7+nGtnk8doT3+znIT58WLTdfWNE/yFc+dmf20UahXOYaIKFM868DwiUOgO/C5LqFe
eMboQYo5XO/Bj67djwcAATVaoASS74ZK3YABE07hYaBx1wOQJFSebyHtQIzIe7HVuzuwk7P9y1G4
03SRKzpj0hhUzB8ZJAcSy6I7fALnlPaVLo32pqFxjX1tC3N4IAjf35O1omEDKnoRdKkAAfvAnnUh
L4PLwbyjlyAAN16FpHDh4gFWzdR6Rye/ZqPRUVEEg3TYzygCKOZtLx1/b1Spu7omnEG+9H5NgTk9
/lOhy7YP5ITssdgxvsqQdhQt1UTs2YODj8oROJTtjwXH1klgEp8mO2gzEwuNO5TV5OFdJW9/By7t
sT3Bx/nUqasLf9/JXGxhCurPXJGQW743KKX2V9Y+QBZtU0206DnxZhSUhlM7Azr8OCVzT8VGbgiD
jOtKCxxthXwGUXwIqixDpYMac/ruuRu2uxFVZZldjDYwWmz24DFR2HitSKywEJYgVnRN8C5c8z9N
z9rdF5Y1rfwxskh+o8z+IMx803hidjXTr7flal1gxw7kHqzLjTW1BE7JHuzkABwskT2QYCGvqSV4
zd2ejEN4zDufWUHvNuwU0Xml91L/kvpcsTRSCT6LZdD5cyRpARdWBZK+NMUPznvEtiXMjqwOPLDe
Fj8OGiRBPrABybKizB9xdIj9CXoaVcUAXxWJsn6XiOeu0EEYd3hAKj9bvGJ1oYnOX71rF6tsrHKj
kbDYrk7DXW8RipZQXETWw6U7dieg7mEcRu4Gjeaf+0zMq6us2/4J3qJMJ8W1NkLbGh0pTGkGzmSp
US3AGpM6YnawzNKN8mvQV8agtMyQAurV73RjpyNBRAY1/7DmixILKioniDECT73tYPoJ81V27CwI
Hndzj7M6RMWConobkOoUHBUMTl44+l9FncTQkVQU/ms4OZ0b9Eq/HEKg/Yg/qe5/THSrAq27bCAw
DEE1J4bRqF6tFPkqE5drLgQMoO11xrmO9jPIGcjaX+IPmMvYR0ynG1m9B86rxOxAItymTFJysZ1q
jlEY5abB1iZ7Ha+Fz1ijltvhV4dT4vH7rrfLkOHZLjM05k549tH2HqjLuP5h3Ww5OyGJ6l2KckW+
bNjZHwoJ2JCEx0dHvB3s4BMsmDP4p13ARNRowF6n7hQHAt/roFqq65eZA1+qr5c1LZ8nhF+wWbcn
2L2fl9mUtWRCDfox2/6Z+zxrS4nbAXd1l1E5t8YcjxAprMWOzKuUTN3o86+uTT2thTEmCc7RWTcT
Kqp5OmvT6+5TUUUl+yUWhey84q68ZICSJt6+ymYIM6FBJtq97e9RqhiEQHEmuj8tXuQCQS93Is2E
11FECcfkMCQEWraN/F6yVF5AkgDmq8gwsVTMq/NQxp8kF5IqvEXIWF8G/Rosi7CJX/ozIfHZ+IjN
Jg8slHVf59rwo0NB4KcgylQ2Vikq3O33DhAaEThYsSEjIsVU2UDl7WzhEzrgKEFETXCIwHVpcT0Z
jr//Qza7tf/87cZf1Yb/e/U19ZRorFry7wpbdlsQxTGCMzC+vCwtXQyyPML7tWyOXMOfkcIDYBzx
ehgzR7gkxWOjxQrKqkZWHWeZ5Y9AP6PcOXP357vGlGeaD93KtANK9NKXk5krcthdOPds5VJW4ArS
kiOS1cwwkRIKE+mTaNXQW/28ZaHsBaBoue/DO9HGw1OUEemP12at7Y+ygs2qK0Xrea8PjaA4PRcd
Ib/WFuVkUbbxCX+1GuHcy/HxcuxrbG4FYFOXAmoBEJjJoqhbaTOEp9VgVn3MEMiBMpgyZW/JFbak
PGCcO/bVPM26JJc6cOSU2QddgOZ3L0CBs0hkT6CQW5xFVqI2Saq5I9G2GdQx5/rj1/Hqonbq44A1
pu6OGC6ef4F6iY2TKJXa/1aJRJEldF2nf0sMFUxlFGJ0vwr0tPMTdhJulEiA2+/tn1aG2r/bsy+w
HPeMExzS9AMWGliUzeii/O3pYUHt8nvJ9O5Y6nG2sQFtKEDvA8TylL8XNI8nLp0L+AhOQXrSz8As
apwm5Ux1+RSWJKHI3VXj7a79mXyqJz7klhGj+9N20wVnSwyGtGVd9F4XolyRXgtXKaVhJ7JH2tLy
AFGttgtLkTRjSdiLvjkGTJVQU2+NDAFi3HdHqRoAZWjphsKALByY91y01h/EYNGIrc72DgPbEUbI
UDJrYu9wYT2E5PvmxZRCCpQuH8z8YVXBipOT4+KQtV0rHUC8UiET4zVT+SkIQNEQa0RCvUu6zjan
ZFXo+KGl79HDZ3HTSufnwr5UF7iXwq0pLBV3gJIdmFuPP3t4tI1QTcCnILCr+u71uoWeP6/hl/EI
gHiq7qCvkH77fkHo9+Q/XCAVTGGkqQ8IulGw+vhMVTFFWKyZp3fD3rAAYHx4BOKBb2kLf9+DEydI
vUYy2ZdHdBTQZ8R7/XH/USSBuKnPb3NBuEB4kcfD6XI3MC6o71psNGQSDANkvqwoMDHBHH4rdDsZ
MpXffAAeplUqSd4jF6nK9zYiwct423KGHtuL09keQLERjLmDcHyDdiL5IPrGNAPjYhzySFDymjD3
jVUFmd8E+Y2cSctzBIBz7+mjYm7qId4LJ/mkPbMHxYaTwg2UjVlB2ur7a2a48l8xto2UvHiJZmPX
+9xxYzakNDsFSB1XKXdfVlzVBuTMBrVIP+gTKON302ajxjgoi7FksKlhC1QiHeP0zz/s+TRzhdar
+ODR+Upc+yZFcMEotvD5eRZ6DS8LkWkjDlJNXZDs2df/HEYIGRx8LtnfCJ/SBmsy8uQwkRysJw3Q
FvqGoXoc3slobo2O2Yle55Ru9dnOlnGODkKDQtTjaMEzS7NFKFYfMsAemVDitM7AUSPgokapOa5X
TZfZBiiknddLXPxoFWQ+FU+S+u1F9kP+oznA/OZxvRPwIWImZ10RDMq7TprY/7v4uiDB1DPI91h2
JGf4PgeengCDtHYatqPcGKAmoaptnpOiCSp1iPJXFV/1pIiXoaFaX1B3WM7DIoqiPf4uJHveT6bY
18DGDGKfwxFmOdrsoKivh6M9hD1z4wntU3Q4WdvubE5CJNJChfiZ0Tvjrx9ut7CNs8WsrT3CknF+
zlkVKQ2P37NLWViJR4y2pV1HG5nadvpdfgyniZFoWN0IX3TCi2u2kyeiRnaZ60FmLk9G3v6KXmsu
QALi5ToyE5osqfqg1nhDzZxccQIe2uF8cDlljQqHgHgzz20JkoQjYqeM2NVzFhBSru44sG/pxIPT
N6WwdXZTtSlwdMDKo/+1wUq0TELTRPzVOMEHp+bICP4E2wQ5rQOOcGQwChWwMUV72nA0mEyozUg5
BDMmLJJXF5oT3i9E9RxhMe4IwJEAxcEMeaId1A4amSQyGHAC5BOQpkVzwUJ3sy9Ir52SqsdNTDgG
0obKoygb8b8Yznc/pJJhEzX3flHtnIu5B/yBTJkl/I4jqSg4wXiHBvfcgSNVhzr9R9XlosMzsTv/
R2PzGAgrmIX7S56GuwluyNwPZT4UNeFjiPScUX1d1opLccM0e1mqedpkNxl9GQ+dlBd+EuuX7zDJ
fVbH5l6BVESj+cfLPxkMqDXTGsljc9K2txGvVpeOGs+XX+MplIUMtVQ2ZRpt1IGNGcOYUh3TvXH9
zQGzf1xs4hKHTpA18M07gVX3hPMaQczenRZq+aTAZBEY25jO1DoYGCdhlYOxR8bDQFFMKPxtLkua
En00yaMXwL1+ymytL4Gjgyvb5KlFhxFWpGK0+RVZdxDiVUwCSaiDWr1Hm/ee5Ikv9sAxrOF2KNMT
WdzS5fDifksfawFRXuDusqzgWWV855uWMJqd/tUwjnloFWRtpJDGQCCgTec3GDeRGRZXC/qUNIao
kpk+qT7i9wehTXr6jC5rnpSsKB76hTOvtiI4RwQJs8L/oB2wTYUP+xE72AjQC6NVsNUza6Z3Wh1J
oH09cK+3FOY5HQPJ/UJ5cc2DwfynMjdziLx6gppPePxGWs4nDT3Kr+OOXbLIEGZEKtkLhwJjK2ua
Z7dPqn8cU7ztO3fn23wsKinq9dTV2+ZRRUNwB3v3W/hKi1xXjroMNmO/f+aMxuNtWEZ7ZO+f0jMF
h+wNb7s+OhUsI4HHj+sDrEa1vj9cWPmm0e95mCOoABL5LGaJ5FgHVOfQE2XaR1BuVDDmMA1dq9zA
DK0vXfv/GXMkdldHxuE20A5cHkblbsrt6U1BWO8iOyNQ4XOrQBI0Rx3IpZ9jZnxdUGs+gc/DDsfN
EfgdiOlvAy9AVGXnNM3q+uyCnuZ8+8Ahzys5IJfz0qwfmz5SzokeNjhOTrKRJu+7M0FVWtJ5I1YQ
4dckkrjr6UGIw71VZkKnZr0lPQeSP8WPBYsyfxWFDBffZdIpmgCWYFFvYeEUExCYNBR4r7QO70wq
p9SXuZcjVcDw5w/c5Tr5MA2EBDd78ecXJvkWWKGE0zNsimCSFh2oArFFV5yESJbTS0XsCrGoEW2G
qNaAuwQPPs2uR+ZdujXywyiH1xtPToZubhKHjcwgbbxOQ+Hnv7g3rZ+8QTbOTTW1NsR6EMLojaeX
4zm3KP5jR51IHwOQhA62X5b74nLFYmwiBW9Phqea7gSTek/uoxClOOzBgQzbNgxSxg3NGmuu2zEl
tzbaqs0VAKg5yzLu8DbosrZGjl27eKXBjva5fOHhGkGLpCD3C+4CERIaILngusJmFfumKz2hjdJO
T+PGlZDiZo/bY93Df/Q/6QxqGMKhQaSznvbweICYU/yLqxPU6tjBwLhvE1UBQaPTdSuM2TiPP3+t
kxvtb0tKERDW8X2u6yJ/HO8if8yC4hsbeMgiMEeDv5lbxLCoh/ZIZwoIStviEIiKn+ab9nJoxuG9
Y1WTHFRS0ryaxAEgPBKbKmy4rGoPY7JCnnvI04FpZS0zh/UiAhyHGnjbxDL+NAyT4dUjzbj5lSfF
rakeSh6bmsunTHp+wjUmgWrJuqikkpHRJzugJy+I5NW/EUm6aFn/trsA57fOAzqOkiMj2EpdcHeu
QJzHRKLjcuLO+m40p1wkcF/VN4Av6taFBAckll6/ZcOXXuVwpVvmc6t73TkLAWtc00bHdaxZpMZv
P9zLSSnLuV7lbZJdBZ/K6QViF9u/5WYUMOgxkIu33kC3l7h3/TOGyGUoIsobpof0eQHiDohdKwdd
b/l46D6aCd/LC6+axP7BCapyHvaHZjt3SlbT3zitXTuC8jPzQQfmWJjIbeMD3bghd6sxDwb4z483
iciufVlkZbMa8R1Dhbhlpp4HXnO4kHOqZN4mXo4yQUKj4gmfL/5fWfZxH9nzR4c/7gqTBQIYcOZc
HxW9U3vdYDuH8HPng+7tAxSpQH0ymLQlwC3A0EJ8y8J3ebskyqR6LhF04PSGDJ2dgjhAtZw2N4vl
81flpltl68y6bQKERKywOGISXPuXeYu4s9HcPB3g9Nw7w+Dhg20fUZrJPCHQaXnvyhmf1d/83uBw
c8O11N15Jm5X3ptEjB71ssg/ciu3TQX0ZFRMW6vZYJJSXaK0vfcEfVaIit6gRp6k9uT+dKJ8nqIZ
ymH+INdrwz7qDhzm4FQ89bBrwu1mvlJXu1oYQCnnJKzfmYAfgeaqGRky2jz5I1ODtQxmaBVE8FxS
scrKkDdwKPvGieiVWJioA99psLJl7J0taLMhZIJyX23W4G/e4lHD6P/MAL3of1ZTEGTS/P9Ig5RU
zEu1VyHoa259acoHZiaSv+o97O8JjSBfbxnMBrtg2ujKh5e8N5xxL6pdTCIa2r+4O5nHQuhS5R7D
S1fOfYFYmHWdyhyCNfU2O2EPc+9SdQvCebQrIpH9EIVrZldJhDyDOu+2Hp8nBJlaKLsm7SQbUuAQ
9prhWWe7bPGeSKeaHrCc1YCsq+uISKgk/JT7AY+ySvw7X1tiHXfRU03rUD3hI+dhhHIVThnv8BrZ
Moa0Kk17uLh9Qcbfjx8DW/Ms+hnPwFogMAep5qKFcv2PZkUMQ7mIAQd2EIeFQb0f8t+eCAaYK6Tm
0zGxe0c43HbNYiuRxboUodg1G0bpGs4Z0sPy+G5X2VGBNwDbHiiKXDxQiYKeotmYNEBqxJ8odNW2
PvHlFFSt/feAlQh3BvNCNy+f0E9nPPCdmf/GSaWzSk8JcgW+gV745fFVHnL2LsEQ2KCpCbeDdGvA
5CY+9vsdAS9uQ2m7s//0LFPlo1IntiPDgBInpottdzwC4nvPL7xe19JCiWMgy4bG+dtMmk0qleBL
ffKlZIbN4fYPV6rEITBaRh6nnfcnBtksVN21YD9RnmrRgJlR3eoZF2qdIgxY8Tfqq+Ixy66XNNyZ
QXhiQ3AEYxIs3W3Kbx2O+CiRVByRRq2fKOfjT4G4rGKNkxrN55BG868RNlb0GpFWYQSSij6Hq+ED
PDhzQ8HQHg7MAvcOOybV30eakva555HngG6ciBmIWMv/6Q5qKmnjF55n57jWH2cERlu9JvOasRz0
jzyoKeE6jR05I8JUCy+ndBMZsPJiK3f7CCoNvKBZ7dQIK7zsc/7XKbgWIm0jLAcy8udX6ptxa9/Z
exNtjDc2w9Y5IjCKwtX9oM3A/yV888PDu6Cn261JzmQjY5ziKGrAzi5SB71pVg9bSIk9xzldwggg
eOvh6ily47S0oCa8Qwix5TAMjR8tnyIYn3BElTraz9nBpTraETo2NAjvJTCtRO2MpkHPTvmMkUKQ
+4/wjq8/aoubYtOI/ppJfveRVcK89b0hTge0PRlnEKckTcdMzXEHLFmSE6kJe8+eSTmtFNSeXPId
O2S8SBdbeUOjFxT50s5qBRM7hZIZDr/xhvAna1cUAeV6vGixbRVaouUrJMQCUqb7FXtFqbZL1Y5z
nzGwcdFwJVRRVeRJEdoSSvax1eZuf2N5bo3j9lHYOulDWOuhXXXG30a6g291vaFs6h0Hk1FVt+Kd
xlIXqZFFlcwLBxeLvGnqIDfHGU3v1LSOcBy3JZjvgR91Mmwxi1vSKU8aKehmQM4YA6YLQxaupQNk
9ykoHwdQEEsgAPff9FV/iz7GCfIau8FUPbNsVBFnHSzNH3ezdYygAImbR4zQOSWSO2SI4ap1pbWm
b2Ws9aU+FrqYFw6q9IocP3RTeBYXZcKo1Qea4h7UuYRfFp9dsVA4aE1zwngMD0iGKDDDiy7AeYOq
uUfgx4N7I9pvf3Bx1efsarikRXulYG0BZgwoI22HQMlc+w91ZlxUSdr5d22B1bCpp5RANFZ18DAD
Rtal+6QLD7HEKxGdMruYdxcndYwNoh+turQi+13Z59xAFPXVt2M9Gi8eSVKsP+cJNgYfQtIDFLpq
8NzZchkspNxdb3pQEJKfNFjJzj1OuR10fMxNbhB/ap+0cIN0bdk0Iy2kHd8omv6rcwzYzkSewzcY
tk7IkiY+gYAozq9qtxXljmK5LdytGjRb36QUFj3+sZlPvIjOtiF/KVJK1yYqptSbyjIEZOytSvdp
hbZqlLTmDHkCI2NwjO/AOL8Av1M9yFQtOQElqtuSckWsZwB+LwztRkAeKw+tsS83mgDzbity/9WL
oeM9rs2mJgWKmEPdMv/u08FSxHA1dDsY06nDizi0SAN+50W5WJTUSQUXM62+BzX0vAsfHTQ2Jpxj
hqzlD5rkg71UmkemyHYDtwTzOUSorNfcfB9RZ8aoybRbwkyi9xdfoxdkm5cTjwFM+b2FvpoNc+Dn
o8GAxinx9oZzbRrPeuetOgd0em1s8kpwj8mZw0KMAtvaKb/02VXDfUfVRKbyYGXfVKh39MqKzPg0
m36DbAxa8fl0oOdHNhOQjA8PbEghLKxaB36m1HPZ0ESZQMI1zv1KMSJEC6MBEZKPUYH4wmcDIQiI
c+TPqEtKxdrK10zjvhqXLD2MQmvwOiPP6c00/Asj4FCVuc0OsAMw1Dqar3dbqckOts2C+3DvuVrH
gRKiDf1WaDIX8COFW99gNmunjT1Ep0JS4kJqLhXpBAbLLntvbgIo3X/hyQ6nkJKlY8u9QVsblZIo
0J77SFQKTMvR0ErYgho6PdopNC8OCUloXS0LIyWURKotCQuaAXrHp0jYvJlEDlqjeqZhxlupYZ8r
eZzC0NTFbfZ1pSOMSU7V4nvk9d8KTs3La7T50IqYsLcdikS9hmRGOXbbJnQ5Uvka7KkMDN/TEwJl
kKFMgU1lvB0EFZqaOv0FxZaDQgN3ljCCnZ59jB1OA3E3eK9gU7enXkqGxZww6zmDogw3iaJD2zm+
9EPhmWBR1uihN41yp8YmnMoswMRaVgMut8hc+OI08TTuFgk8lAi9PaPxCAj2V65OM0KLnHdNqIe1
YQBfejmUdq1IkkySpdsBODwwjg6K7Qkpto1ZJxUC5SrCsyNKIqMDrSMI8S16x1E9cupe8Di3T9lt
gzNOmFvip3AaaHNTOGi7TlW4jLyADv5bBBb8kBdU7gx/ujegy9hK02kQFTQhyqEU5pEKLZrvqKt/
UdZaZEVyyJOPOT/a0J5jeLMy+KOSy28/6+asgluNZqmTFuOVHTzgbNDadxguiAKcOnUB3XVsJQ3L
Sz2Vrc5ng7/U5NQJGAlNQc4k1Wb53h9Jal1uDhenRd8emcd0J7Xg5groR+pgI82QstmfL+mJYYfI
gVb4BUL2IWKhlC6wyIfA2808+62KGxRxcqq7qfPRypuYiwof8eWJHJRsWFkvvRauY/n5zStGMXVH
Wte5+xxwwCFZ4xXRe5bdFpLUGk5IVwvxIMK4L5qaMYVkFPf7+qG18ee0JIb8xCs2W0aHruqneZWP
0VjEnciy7W8Hs6DQ5watfRiN5LmBXdVa7Cl3La1N5AsZQFo4CAy+MHP79AOYp/JKmme7KH8P9CQn
6tk4Zgwa/p9/rdxDGl7fXbA3qYOGkKD8YVmLBBzhrKJvle/++HGNmDCj5mbdcrhA20zSkMVfBKv2
EHi/oIIhjuuOnZJkxUcd4u6VO4F0MZ1le+47kmZae6xGbSap/t21OrRGQ53bqBnPiDNgi3b34IHA
JftWSe0JTSYSYRRdpp7CyIqULHtaQP/te9gSSpwuriYVUso9wfgCD0LDh0UU7f8qb8TBnMgpB/H+
bImy3zYUQoSa9jti33YffB0XsxQpBZGo3/Y9sIZfA8np5PpNg7mWPwMsFe3XDq/xPdK2CxucaPAZ
hFyZTwnKPYv3wLRE+L9rqhd1AeOTLqj1ValkMJZMF3MXkmtzjTPmnTP7JH0hVTmXuFMTi3P1hcYT
uWEc9hw7fYoXkhW8ddhf6dUQVoI06lgsJ1plSX9Vs80lKXE+BF77y8F7ArYEYownhYyCq65BxQHz
gkcKejbIlNkmCv6k1xFKvnp/ibk1k0CpXTPF/4SzQWHYCG52YFyCMQyziA8YwVXbcJnvv1K8T2vb
yNOSGtNk04OQCff49JdVo6h+dOzNvILhR6tzYzF9eoBFiNwP7JiifqlJsJrPYkibzuRtjeN74a+C
NJi2VnGkY+9vKv4aWAkwk0tQk9+Nu6y4xL9urMblqQVL0uTG+h9SYGU1XPb0UujUzE6ctV5Em2xb
BM0BMpy4YRlrbtMxhJAa9ocD4hgAhFEmMStXiMFQg1mlvYYlh5Z1e2k+ANxlomcegqAw2P89lBLw
LIACHGmJRL1ML9ZxqZGK6Txe6ZHqwF5bOEFB0v8KBsuCwztQuWUspTM9j0XT9qAQ8mpV5tvXQkRW
EZjyiQyR9uBHzDwEEsoW9qkJWCf7gvOThcc+C+3x3BFyEkRe18mh2iy6OevE8HTyZifV6PvWf1TM
55SJOqhnkaJZdBgQa1WzoLxkEhNDoLMC3MtLBTcEu98mGyuQhBIJ9Pc3RCq3xoPBNpy5rqhx4EkW
msvw2LsLBKDYo6e5Xanoxv8ug3ewFBQFE2IhumhZjj7deFCJaFQBMBloDYH9YrP61UiUymaXyh8k
DYaGkfDklHu+BwBjjcxUruCsGVtuh4Fc6RGsQFMb09RghDnt0kTQccFwr4vnN1SDHCL/+t1jV8b6
V6vviioqwh1/gG8jv3ILXEDEGpXtjQzkbSOC9l7fYRkxfBIY0xLACQ/d9DZ1knhi4opwWA55ofbj
GG4ZwOsYJaWTx9z3fyfly9niGFaxAEv3WiAw8m11AlXBn2FDHMc+qRLd/0jEzfI59AST7TZ0E4kM
YoNrWbIdMTYyehnkb5MVvjmmlU8/ttV1RHaiWbOfmKVrLG1eoLyciS4DLoJBcBhyiefbHJBEgyIt
ICiD2NVUyl2U7g2e5s5DzzoINQY5nm+NUMua/O/KUnVnPizViZVC35zdG3S5h/R4f8FsVUHrd4E7
2GQ86huQsRZN9sU+M5A+9tvF9IOrR34nptVsmjZ+FTYu06PsniBgWREjGPcFOL7hIU8NVGfggSD/
NDqH9iuFDsFSw5kqe4sRtTb6CkLtQDS/5Q35aHzlmaGh6avZQqCZ4xfGmFVdrZamGBc3+XcXgk6b
3T5eK7OH9t0VdHgIQYku2u0E2Hwyhm5QFmE1gz14/7QTtdtfaiCywLudmdJsP2kfwoOEnn9Q+4oC
obUoKXeUNNRCXcyYufwuQJKLyJRm9aQyAqH5l7t1zbthix1JCgpCoqgsD6LmG05hU29U1MlzRYtP
FHuBwhaTKLzmEj8/OQMmc4j92sLilyIrbk/NdvRYRnPmQa6JiWoNPbAnxNbilpYAoKF8PvVQeKW8
wzJa+8YrsoRv9FiorXx6PB2GrIBzMIcPXFJmDas1SSWUBkXwBuoO1YzOnwvaaYhmMfnQRstWFixL
FqZcYqQDTzxtj7iqBI54nygprxog8xoOOqcgAg7HC3jOGiUDva2Ar2xauLNFGWKTQ3xuMRxRlqqu
sKkFcs9fsBsPxJgPugxnmcp/rQB4+1PmuJw/+dEtS/7Mnl4S3yFzRfHbe68Nz3hYfTMoTlKEJTeJ
C8NWWicmYP1BWAaNMvE6p79cgHnaSu4OMyOY0vRjAzmADz7t1ny0SVNZD1NkW4PWyXAsmKp/mNzd
OERh4klxy3bwosEcpggT9biw9LJoFDoOMUcq9ugDGNvE6cMAYT0x7R6SKIVpAIqdw7n/1ZthSHEm
+PDdHJWv338m/IQh7V83q/WAQ+g6NhGL4urepFnZeLLw/e1Ap+/tQd4f1v6iJlIZ7ObHumOodnte
6whlyRu3OgHNnpI89K7qZaLJnPbJBEsrVV+ktU6dn91KE49ODJwLw4uXyMw3qEIPzB0SCaVbLkzm
rQ4noU/hqhCf69+xvhVv63aFWrGkpb6uL0J77vGAknqgqMuIOm/OD8hmVb3H8yFECupcU/q9JgqS
gnSzRW0aWGujEJ5Aw98AteF405wY4PIXX9RaI344crHzCTrQu2W5KZLtuKzV9AD96B21ru3LtSJP
TWF+Pvs2ESVbzy0IVh/wsEHnlILu1/9wzLAbAizVmmNACm1V11dVlpeXX0jvAFC+hB9Mftp7rF/j
4Bj9HngRKFEtMmQXOhVgArCUt40I93UiTi7xb8jsQDPSGTpe/HRd1pQ3/9gJ6RYW5yU9KjvLLO52
aaqMylxuuSCOWTgrc5prB9Mgos3EUUwox4HGrGgNMJhqx98eJQEUYxX8NUNLNIv0QoPEgd2s+wDR
MZ+oY8TBK3+MCFSAYh8u2onUbJs/VhPKgDKtWupzIzauK0js1V6MoRqONWTgcMsTNIPuy5aYRBdF
4Mxgft9Bam+ebF9Ip+dCergH2JzXfdAaDbHdSEfehadSutvEEJGsFPnKbOjQ0r++W9VRITlzz/rW
9zk3mg78oYBt9EMyneaB5JiNdT/iM1XYFtOQ74d73yuqnf1OVpCEsviTlZw8gXWE3SJmg5oZtgXG
Nzf+X9znPBd6fvAdxbK5XY06i5/ZmVpSVNQQBaqZhfV0ysbU0e5SapNGIKaZ9JDdr7mwN06Am6k/
8ya3fWjmpnidEPO4ZXzBDzVFr8yHN6WWttXoPz4pTUrGj976PQxIJJNi0Tw5kOOWNzmyGGDkVk2i
7nciP/+9U8ZapePd6afKcd+q5GfMVQ8n23o7Kxgp3dALsdeLy8WqlOECHviKgahJ44boayHBaACc
ixvJju680fhZJ8IETmAqL01B3BO7/Ui//RTuLDRgMSBbR/7dgPOfNBOJz3bANbpD5JzxxaWgiS/c
6l+h+CYp0YlhBUnJW3c5M7dbLFuSfCJ6+K9h/v54W1ueQXdXLf6CeE3E3mdaZV23TYDcoL5FjV6o
zuN6mEiSEiQJ5OBbGEN+CIhbLyC/Q0iKaYcAb48AU5JrbIbkBy+IHDUZsrbt7y4mq5VOCSpSFnY5
X8gm+BYhVRub2Ur8AcBgPPJo4Zyteqova496umjMF07N0CwWZnaclYDEzc8L4+HON0JfyBPr3wif
6NpZsVOie6CLBphAauv4mPgcfDgh8gtyGMyrsm4tD9JuJio2+eMYBdvzfb7c0XJcjG79K4YB7nZ5
qYjRgBllvnizrRFSoRSwAtUHCcCNTqofyID3FozxEgya4kN7ZKIfMaPH0UQmiO6oKfVqNdo/uuO2
tjy1pN+a/gS+7jsZbfCfUJEwRvWgGznPHsVNYVFWtPu+pMT7sjmpBORLSkhRZstyvLbBmYOvOPJP
i6mKPiXTDzWyHeePsEZ6D2hbMQpxdVc4+g9I++VK9Q0O6PfrnYajGBQ9ZJFa5VdYnLgwCjmR+Fe8
CfvHr3JYucYPgY33dceOVVbUzD8AFbN+fYjOkHmtKGphclJxLmqrQHk15yEYbprHKXGT+NHLicjx
Ng7b8FctQvnLaMr297dDyP1evNTX321qksCr1FBWWasL4UjElaKwAo9ePZTNE1+bvQMaJ3q1Hk37
gFGKBmnYp+nYfENS2R/5x5MPONBuqFS/vknAKv+5zGEWKnlz2I9Ux+BKZCvvaVbhKO10SUUHex27
raqw/+x/fVvxbi72lUezAY/AWhy6ZHSjn4Cv8ecFOS4Ksue5dQKSmCu9pAtSTEmxajzkpvS9ulrx
UDDcNl7ZoYIzGttMmKbZ0PMisUICAtJwsRJWU0K/MM4mrD+wSdvuAOO8Rortj1nF7tOJHr9tPchH
Nt6RddBF0vSDWcmgwq5zE/3lrwvDiDOnhSojTeJio6kwSKbg9PXmW2eP0QeoTG02yIhFJDGO3t5+
fcgc74PZd86fxGfe6B/Yef7CgGHeNoWhkjzIJ45vK09bHSSqbfCZ82C4g6DofRmKHiC8gYdvFtfr
U/aX56ZjeLpHsVaeUVgYslB2kd2KRiGzHGDM2ZYLUePZtAKSGatzpB4u7a728INzb1Ce+xp+nrfA
OcFZRkv0Ogzdqv4CQqp5cCO8+/OODvYzM8kGDUZIUG975xHdhFTTvRC+pGMPO1iFjyrPnd4hOZGh
pgx78oovroDfOcDWPoitU2PmiuLB5x8SzlSH3zHCyDUYxsI0/wznLFOSZI0AZF0meQ3ArHZP3jP/
6pdxgULPlbcjloGepGkBwRDtmak/d55ebwl1Bl9p5gpBtPEuneQ18wz4QBI8LdWCgSP4qkYv9VpV
NA35ydNBn5FqRWvnMM88wtpLk97PXe2yDyUwgm+LgTs2ZumNpS7ZPIu12qJgi1GYRfY8rm9rF3ym
Rc3uAyusacTlwumeKQTmG0YZfNxSm7sUUIRIA0TZZh7tkqjt7Hb6PsTCoMke/laLZdmTbjIn5YB8
pb62esS/VHJT04XBvzzCwJkt0/hnmTmSJBINnAa3iFCz7PPHKY4kdkUw2/Q9Kra45BaSMP2RgEjC
AXbU/cgU/ZGL4vgb2gY9+urn/OZat6av5fBWJpi4vYl/UFvBVALKi1jkZ5WYLgproQi9h9dDt35v
HxZjsI95J3F08ZIdj0udN6eLzhziPHemxLITb1qgHH0SwVYouaedHw/wcEU6DUiBLeViye62RvoD
z4AwuHrDS2NlbxHK+ybLCR9OIgr9sJEP4xwXqdB+YZ/Ts5whUM0t+JXpuo5lgGorEPf/z+FeNVae
QPkXUaibtXRE2xQoqnZ2Uvw+M37mKLbcT1YRuwjaaZsa4cKXK4eLwuWS8SjnyAzTiZmLg0Z4C6Cy
A21eCA7HbGC4NrEGovu3TDtEmDZpCwIMfvYe7hYtHLXzXGMAjX7EWwtLEBOyuIQXoFBLoVQ2POAw
UJ1xQn7n0k/5/jEZ/2htQEkPwTlw0PtJ2gFzIMp0F9LR883GSG5aWHMgvr64l1rxWJkRdiVO7yhh
VxPFPk7wV7rQxmxwSHIUqLu7FgBDKmBEgOQ3SJkcuT1k5lailKhMPdmGIb4dMcyHMQAMZmIcdzv4
jxN9S87HHKBsq9coYHeQxAr/U6T3kGv46FPr6dcqn//ARFitccZgJuk1jvYk71c7DsJhXz4pDgt8
JZlAPF8KE1yj2yYLyUGnkHynsRWQB/vRhHL74siVAeX7wrywrJNzWOhA6j0zht1sT4Ih3WHhksGU
ocruFzZ9cYbVXfIu7xqRdPwoaviD2bClqwR9er39JGlab46eV9Stmu+3bHCIkUOCUov4n6l4nchu
cZlJT1NR9CtgSpOf9cQjRnUS8aOd7R18EZRBJY2PPx3FgWz0Ub98rxbxsbYSxsS6BPr+BmPoIbcv
AL7PbNkMJfAJtA0r9IUNXHevg51SiQaP1pgp9XcnT+PiIXrVyTDzvr0EiQdQmJjiH+W5hKADiBPD
/Gi/DPjIVby3xqXHCaIbFa1Ff/nM/gGy1WziMEtKJUj1m78Vp6z9XXGA9NC8dKYV0Mq5ID1cGOBg
DmiJC9YaJR3N0N8cvmFq7EGKUNZqcOklArfW62mYR0b+3rohMo4m6C4dCaoICbfeRyk9VeX0aee6
mcTH0QEClgivOi3zkRbkt7F0MdML0yVCA2W4oOg3xMvOJeOo5bEdEH6VgTdXlRRsIdqGL7QCe4/m
9JMtjwZsz5UTGyES70rhP2HvO/UVckmk8SSMlntE23XnfHllKM+AHWOWbaNj9cAzq6PXzVZ0F1hr
RF54/gN8y1JCAtJog10sxNlaJHbPjvR7pgYQFvvsPVYzS6uRwkoMZP/ebjSNXjp0Khq0oeO5WZ7R
MXL+hvA98dXrrS3BQ+NGg9U9CReX/DbB8+xpuv7rbnhdgGWckrMhyZOy97gevwjyvHO+CxC+/aK4
uu+yhNQ22H5phYsZPV0DPrPGNnxiw3dPIqpQN8EbrLaVfMyuLIIzq4+AmAkwTpRXxrUrkV/qPokZ
gcyP32LT71QHKF9koHFc9yD9coAnPVSxILHOttPcq445P4ZRE6LSLJb/1mFWKosbdmUVohzFI5GA
zM9Qb8nnaSbHCogJnN07jvCo+YwmYq83FqpJT+10NFTJQBrGuORz+PTabgY0IlgQtQK5oEdfXKHr
W5qxKkmJhL349IIco++WVXlI3/lTTjCQ8QmqrQGV5iqLg13vU3Gof9Zw3qsrQep0Vmk8D0DF6V7r
865n7CgEgJB0Yqlx6qEVjQez3c8/DmJsKYfd9VDKwspcVA2Hpwqv5B/xLlnvh+BAT32jIHjGRly4
AtkhOB7re9/YrzgO1qPyUikKpHATmgUMrC9zvKvgutQdbMjVUuhgMgdOMMRhGV+MUesMOO5d1tff
m4GczsjBpMaOp3I8/KcaMiC8J/YeJh/xSd54/o33kvXeqEDPuy1eXMFU/eEuO6CluBS3YoIni7pR
Jr6ebxbKYL2scmM6jZjfrCUOvNGoRGtNhrxB/PckTuVqDZa7rSkg538JnOWRiZOlP+xPNGYhW/bm
r4MNY5xrNSuzwdzeQ8MYgYUlPkWkFjEHKcenSc+WNTEfdEL5p68RYBpxv29vzAVdKztR9bhsTnqs
0m9I1N5QGNsxWsS1Z3JmwLQFWF8A36y8LoPBpHIWitoawZT8XK16Y9TuUkkfhHFrx9z/9YdSMWTI
TZM7o0xwjrbJNSrmbhQHE3q/YlKqef9xopRErEQn+pNAW/USeN6PA1yItHqfVa0z9euDri4SRHt6
ilUec7LRFCFBxZsTNj0l+U1clGptAM2S1FSdcZsUCLv3m69U2iQwK15AgBqOaT4seS5DnGvcK36l
P0WfY3xH83IOYII9GZf0BQoorHf3WG66pT5hg0RdHg563kufJgzR56+YUGZ88VjuQccK/1cKmvpJ
Jyj/6afkBmCbi4HK/cvTag6C3G/qODx921kLTHC0AUMNDtXg3h04l0bMugr81FQy2Q83CVopQl7C
wafI1GcB6ocVjAKjYRBUG71REnZXcCulP2yy5aNzHNU+Izx7J3AKk1MRGkDkyZ/9XJ53+z4IzObP
g6D73HIGHJuJSH15fnIcshAdf44lBuet/tGicPt6gJz7xAhgFi0kqsrH6M3nIFWosX7Lklym+bwV
xE3JIaOIyWFkIPQINNLCxmN3Ra51YY5mp/VF4tK0nPtzVE2lkXM6e53FEtaYqyhyU2xZNbxi76XT
e2jFgDi/aRBQdyQ+CFwnyI2jZoJF1fR0O8QWhtTq72cMJq+GIWMSWcXqIH9VIRAhyd68/3aEavMg
o5k52SN0qdjficiCrJuXkOVOoBDkW7cFbfbzJKsYgFfVuFTVcxgcVMqjxmKzbJf3cBfTTe1bWWa+
VTNqBGbxqNuTkejQNWl2usQ4Jk2x8BYjOFin21N2qxqxhTtMZvYl84zh5UyT+bCg86shzjhpu5eV
badrhRzuKKxSpm90xUsoLVBBjJoyYJbkKoblIV8TglIEaY5dJ2m42x0vvG7OwKEO/3nW9x6AgIvs
vFYOkOj2vejn5n5DrqYYhaB7VMpk7EiFsK51J34wP/5X84nB47o1zU1jtgsIxze6GNLsRXt8wOCN
bRYueCvCT3S5k1lDLwqGBlNessp7cifwElDc13+ARnZWcgxKDAtBSvK3CrLaEJNGQhPOcAOo07NL
XmWgyxJ9O6M4DT3v4PzjAZFtPK2GgPXceeGcDrXcFcglF/pWG4giIbzjTXtKjy3PH6Mbuudu3WRo
nKw523ccgJweMjOh9zbzjG/Two3qh6SwuDaHPl7DtX3N2S6pXaBr7tnyas1Zung9fQFydmYsA2MI
GauGhZjhwbgRgZZNSdmmbF7v3TjfCgkgI4XzeXUrnoDqvUAS2lWgClNHjYuNTO5DFbmy1YY9L3t6
ccRwB477sUUpEO0SBg7c6ZeAkURwDw2SuJ3XAeCqoH884LUTCAtBcZlwf/h0Jxoi9iLEcC9VXl3I
xuzo68PlibMLZuwWNnkkUymeo+/BmLrLxblz54Ys6UYUcoqJHc+/uRKCGQq39NPPQvHPin/Zo/tj
N+DuE/phkufLO0ttfRPoLKggkFrB0YMnB6DbC6BAAPJztTjNgUh6FHbVBfVXf/1J99KazbLFRpMT
97JkeRUq2ZaOHJJ/GzoE+hUpKt/o6mG1tCdM9WtHVDenFyRxF/GJFEcl+euMIr0rmNKM0a5Ko1Ls
TQ0taUy/N3aYaeAEtNcXWi5lUsc67ymSA1+0v4ZVdhIZgYFYvMDCA+MsdDmpeYJWnYK1rPgnENS6
+tnuUfir6ouBwiOq0UAxvFUY5IGkBMFVV2SDSBehGkJMUSqgTyexQh0GFDB4yaNWWA3mBqCgsESG
Uj0YYQqD66quX1vrYueeCNouw5cSx8K8pDRJZVRCbTBqMpdxyRbLmLmMgf+vwQLbTedSzY+Bp3t0
BiZK1SaG6FLLEpvrTqfurKY7JROWPCBZ5R7QF5pvP+V4abSiDstWP4t/CCvo87KChOsaanM8NswQ
jHzZx+XIT/j7jy/7fbEoPrDQQjE9w5DVgs0mA35/GIEwnQ7M9Iv3rd4sPLQVIDWbRe7HZ/0NShjm
iO2W0Cw7070Oys1GOkTQ9wp4yEbe6TZlR4hG8oUcnNuQA/nqVky18g11wmqqSFMr61/olf8s87hN
sNLO6pF8ATmiztlWZ8ZrL/+zhoqVqjWi4HsLZyeTMlkRzRbYBaC72d0OCo1c7qJGFX4/WnGA/83t
cI6u5vOeu2+vbZ5OGnpICPgVdHgRRGZdOqrmP80y1k4nQGUQ2nh3JMjlhbsLmGp23gf0C8dwjqwA
cF2MPVUwnXtADW1N1dARPvgR8sBau7qysFVJIXFktSe36o/nR3bdJbvrkTc0IVmhwoW/7F1uajoB
oyDJlMcah/9WvVqlarAte7nD+xxxcTi8/2vJa2i4k4b+F5yEl/68pCCoOw2Ifkuo3FWkuIllRSni
RT9L+tOfiHAbf/nLGC6YxkLOr+6nvJEfMu28WkU9nudZI/AhOVGPOy4qTyJB2Rkaj2SoKdounRbs
1Exemt7EbMlP6CKx5xg1zluCwAvbLQ7Qee26UNVK7WvoV7VJwsJ3ibLG1qEXKRaGi0iLtKijtK1V
zfK3iGCGOBdA3ZiPMMO5Tx6ESQopQPn86RS04CPYTovUubjVziMoM+aBwf9Q9l8EzBSovIbmGd9v
Gf4eZslf6SeF6QSwkPP7Z2XP67BT74s7uIQ4G/4dPQQ+udWdtLmJ6zIiEjzbNayC1pzkn+WBZK0+
VlYfsZz1n3FWuk/XhmVe5kuaN5fOHI2G2mck8nrjtW/DlwbtIXdyYLCAHCaiYuAY1WrW8IcouOsn
All2u0kUe6Dor+ypRj0Uc0l8dQFK1OlwKG2IuWThk8oRomFYKu3NbqDl+DpE3LbsPyt8Bs2ponBd
gQAJqCcYGHQ0HdDpaNQoNHgkSpVKQVxyJ0cXd+TJFPNBDt+aT2Egr0TctoVBUeQkwEkCMeGkbvIc
wH/qf3wMbUOAivXqW4jIs+5J1mmRoMzn7WySPvyPwM9RRsnoJYMeZxPBXsut1nc2PRZzkoIZ+Dbp
1TvaLgL9nQVQLdyreTXBwww2yZWVHdAKvGvQCZ6nlax42APQ76ZJScd/k06ExZsvDwer3NaSPqXZ
yR2nMmhHKHJjmoWKkrzmajWRwrPO0LiadkyTpfHfP776Nyo+oo2ABQfDBpUkzZmV9WrMJ7GRpTqr
d85XCnEI/DrUInCSsNZy7SaxLO8KQxGXA4HDRFtAu4+6bLlqL0HgQVmCri1R57phGnrGi/pGbBjV
CxOioV2R4IsMAorMEvcRMOFxPsBYWoultOO8373J1xT36Jyt8kRzdJj4hCw6f8SHzG0HVUgcP2hH
eBKcI5d7lst4n4SZAScVFM5cyfVamEjJ7kxcdqk9KOArPD1kItWz9/8ai4lN9ZzKzhbo9AXpcdS7
0V2vA0uj0QLddpxgVIV9HfZ2Dd0UbclZopqtCYV4nliC1nEQm+2kRK16/YQzqcVm2FKLjS+C27kd
9zpfEWbKpbNSJDBNbJRGdp7D5WSoCJfOSs4HkAn7ESQpHwpmfW8xDPQR20jxdlyPPf+bXN8K4l9u
3M8u3jDVymeFnXFvwzQLSLgr2PO8DgJRZsM7Y4y3DR3f6F9pDynEQVIBNqxuk7t8yurNR34WZqTN
MBadZhEwDQy8O0RTRisX9qwrugNjlD0CXyBLc+SQ0rPZ0gljBGm0+cSoN//iG6LsFX8Q9qgJKBlV
VDQAhbgUViPiiVxlYEBjFpjRVC6xA2+79CppUQ0XJmHU4ufP1e/u9bhYg75wmkdbmQGlORgBTStq
D7EiorZUt6aXP6UeMc8W4HqKnBzVMugrWX9tIJOcMwveH18hNyTftN8P/gdWPP0Rj6qMJwjhgh8d
ExVFD6oDTjafht9mLhq2wSzvl+DHDsguajSvA6uviALs3ZOaAHqjG6jtwDV/6ryEe3BTiEcSfveh
bRZxbb5ME3Z16V5F2g35B8XuJEGA02ch82g2BzkGhbmlGPg1HOygXbZ5ydgxaqzm4IOLsVyB0Xim
pDLhWLoKgFqGfyUen1oL20Hf0Y1t13owI6e6JULlzPQWGhUb/JkQ9kLTH09bz/zBFcY0vxmOz34B
pmNqxGbaRdzLfS2jUvifAPaxfXvQcI/QBlV/NUJlwsbvs9nXAthhzJoSx6XaWZ+a96DiTQOpdkX4
ReACJrZApxiSel1HOs8cc6mXmnTFV/C1S1w2Jr2u3/dTeHuhvcuXSCDDi/30lIs4lr7lPzXQxzrR
35PmK/KBGqjvtHlFRz1HWvsDqMlxWFisLUMbA5vkpunksLbxg/zYyLMs+wrKHds2qyT5JwoXeL5R
t7HirA6SyffVdarZpqTmCzFpU8KgOHVDp2NM7BlqFfFTwjfnasb8u9JQU7D/lS9Ou1P6FvIBntm7
FVS8Af0mXvqmvxQPge2H7O/1I6AIc9kFnz7el1OD2jAIxRi24RSW1Dcg92gBpAIRhrOwOdsuWOSR
A++KFji6ZpnzGCZ9o58xwUFfv8F5ZRf/NbYYLG8xq0ZuVVMiV1rCkXG+r7yhPCvYfDl5bSxltODr
r4BCd8D3l+WmdmjDs7vvE1V7VGT+iLlET+gADAH8qF0rVc+5fOmGHHDcu+jwh+NUrpPGTwJJfPw3
/+ffPk35pupRe5TKTxkfIXvykHnjRsJ6t9dn4LL4E1Ezt9T6+dhpZmIOePdmk9QUBtHcTm5mfti3
UyzeBqvJx/8tpaOugIWig3QESLAlYA01Vc5gFzCLeuIwaWFR5l7q16tbkJ/LYru4d5hZDVz6OydE
eK/cBDG+nJvuTbwrgTvhyl6FhhOa0orh7pJ87afllU8BZWwIFVFhVu4tYzVErq6wDBf6DKaBnnpp
HWgHXE+hi9QHlTk8qxwfT5/m/3dJeiwPNrsSRKE1+BZ591KRK5fc4ZKJi7kFckTDNhw7bVU1rqJX
P643z7x/Ibh3i4uMNkv1+G4oEe1LfzPq2TrMF2mBG9D6GsoHNQCZErezuyiHq//ueS0fCmqJ5VJQ
MIGtQ6VhRlm7JEJdIwmX/sJaTmO3UnmMygWfPEPqV4noRxXTHm1290oSKCmn+DqXTruj4RztUG29
RHQyl/aIrw+gtNFVyEmXOeMaN1SZdqyCHa4Kj4XIqHYEa2DeNCkaxy4ihkJhuyS9heLWKMWIBt7C
Gkihpzbcw3aMFWhOM8B1Fo4QpjXBBAc3bk9AzthZFoU+0NESfvJmtRwLt/zhzFsx3xDKlMK/VmJZ
9TKgPW9RRB570U4aX+odQk03xIO7fBb8GDoxjJwNJ4WDYSMgiVha9LeEu10vPh0ph7WtV8HmwIOK
MKfsnEwRQsNQGJpfU47vSIrfvmldtMyPcG6TkjEL0pn46bVFUZfa1bcoXzHfDbbsNBrYXQC6MfH4
HNjtNNy75FloKcN8PfpAN/rBRmR8g8d40tqyq0qIvRwlneTZaHDCBKLCBAaoxdADGJHRgEPn8i3S
cEMwb5a4LDMxDa1vy+o4ZZldncqFFsWPeAuZElp4+SAlMhJW8u8NkcfytI5m/Ep5/VyXtkMnprH+
yqh52x43m4pENe0jiBnj1ueFAETI/M8D5HIGoVr4tiKeTCQITKnF4ENJ0+enVMAgUPAVvtYdSw1p
5Qx24nNHI6+HIzYMpbqdTexRdYZEMauLHHgM80TpspWFwsuVNI/Z7gk0tXstKk8Vvy36UE0qzExO
j1n2DN+GHexAP9BEfSkdRKdndA1vOXtuZQS+c7zB0WHHPM/2XnCyS+C1A2EnQdL9HqgaJp3ugOba
etQvAYqrd0t/2OHAsrpyA9m0gKZo52V7J07gMhknJiDS3qEvAUIR/zv7LMTC8ho0VOvAn+yUzeVo
zSXdk+sOb4UbL0P4Z5xb14N4BplKMNnjAAFuWpUNv8TA9Kk/VRVCiX48UryRXpKoe0IcMgOSv9EP
G1TK4YyxHtdZWINLLl8w9yYUE2vc5VSwLGLnjgIidhZWqRxDR4G6L/1PlB71v0JRMJnx8lRb1fQl
pGJAPooYjOwqdDLKFTcglvBx8KF+l/BH2SyJ9grbBeFXuyP6O+V95eAYLVYZuijHkStnP0Dki+Ku
B1TR6iPqoUhNTjG3ih57W7yFsx/6v6XHvOnPqTfLp3/79SomAKY7kj97gZbMviJcruuzDbvgvt5d
n+NZH7JvhlTh/2Y3jIOGmLmFpiZBOHCb3XiUe7MsJx6hhcR6EbGDkuwlwW1oPam0so7S6TZ8q/Gw
CZ0+M75lwt01gF5/cTZPP7eMLrSMNQRx3WzFEIKUFyaAuOufJHo5KQMEPyehwZN2bmouDj4PXMSB
qISXVXVW+4Ko5Z78SOt242RASCEEIakTIMFfV2nA7TwkX1l9P6DvZWFyd798W+tYMkJVAG+qaCg9
2O4+9RHQ35tcgDs4wTLdGo9gV7Wcm/F4QhYzJjlZxNBwfEs66LTyYPDPWIUoyTQQ98uhU04Unsxi
Y8L3d/KXkGOLrQZHCMyvQLl5oN4MsWH/aOUGGdiIbaa2khfvLoSHTIazgETxTt5HsU9DX2z383S6
r7pJXgThbsm1V1hoPO2CkwhSwamRKhGhTh9viTFVtMcA2XfvhdwT9AlIrGf9fGkbSPV+CJF2vtIM
pLFXVN+V9iQNNggBVaqEB84Tm1fefwmXI7F7fSU1dpY+qRRYVnRmoBHEuyBSiteJOrIGoVMRkLgb
IyTE3MYH9XNvh25GRtisQYNBPo4nyHKrKD/MFUCT+4Wss2bd7rRcjsvGui7DVIBcEa0C6/Ij09u7
smmWcMewnMFYy1+5xj2Wc4vdpxX6ZhGaYD/uJBTSs3k63gcEH3aCHG8kay1nZqKubNSyxc0Lqpgj
HCxOK2xRvN4Bb0qrq57GehILZUi597GmImjDGI2l0gW+n8bI+ZErxA4OZwIYFqGUvoHZeZLrRSLg
S3yve3V3kg2/LehXMPQ6i1J48RPu98uG1In3k19GG4Ek8hVVBtG54/XmEJkmJYetufTkjFsaMVSJ
EhnAR/N8NMprne8e2q5+EdDTm9/ke1aK0WVye33lz0ETAwh2jvK6X1kJzknFJ0IIS6M5xuexZFin
3xu3IT3JlPAia+ABovVeV69aW6fu8jWGLhJyd65gZp55CJg9PVmxIWJDq646LxBXLqr38rPHFNSx
QolDXs42U6GUNZ5o/dgip0MfiVQ/h30n9/k3Y1CXdrhWkgD4a++nH+zN2URLu6NjEIWu8cvZo3Ev
SRNEO3mSTDV54EpA3S9rPI9Zv2qcfha3DvRwvadIqmrnhsTt/V/L9JmAj4w86B2vCDtpVwluIM9Q
7OM5bcSgcIQCdntpBR5bIXBuDa49v2J6qY/z/wlYuVnNU5qNq22s3OQSFFk7IQdJLBWqwCdMEXeN
CTA4EwI6XSVytlDCnmaP785JZLWJpbgwWeKk4fS5pUwIWfobB38x7nL2hcDNWJsLQjXCbzo7NH2L
VGaf3i7g9mfk6nGPvfaii4V80X+0Z/d4M+jZMwbRt7AaV6xMZkxbQ0DnTAekZH6CrpiIrCkG+hZf
QuIJhMzbAt9Sd1wx0pzjfSmxXEXUxE1JlIsv0NpeB1xemq12CdZfCRycsnu9gPKR0zvAmS75eJWv
fFKzNDTgR6r/8/RTh4L9fmCAiRErxAyuu+FgIj9JWsBXN+yLiqqTS9ttPwBWdOZ6JWz9rBG2iNs9
J04T8+GDaUP8PWK8Lo0gqEAXsjzgVnSC+CvW4l8TQnf5AcYV276o+W3YWrQQeqTkdKx2httOtmmi
uAkyENFtA+cSNr6PTnrW70EFzC/nDx0u9N/HJ65QJipMEfh9yRzroJEE70P0SBj3PYmOvWRNGxAt
pTae2yeL4v26WGXCtnGmqE2lnnNU8mFa5kRp9uXxKefYNaFrKzmJC9YvZ6nuY6tRj6Bq7YIezpgo
e5TxFg7lZQEz4BNZNakVPPb9n/FqOaHM5r6pWLA/AIAz51EbYN4TvHqqIzBREO7e9ubw5Ss8GPSP
UKHoJJzqXnCzQm2sVja+1oc74L0u9IH0p/kyg3qhZ8x1mlWCyVpKDW00e5SmkC5Q5kkcgqtaICaV
vtayotoJ8ZDGueYQ2CwdcvIZqjb/SeNK4Zp0gTMMXRz7KXvXXlP09zVSASsUR4ffljXVvkILYA3Y
nvGXL+PUjWlY7YtL/HwXHMErUO2FSIDMGP1WXWk9wt4Pk7dhjReUqX1ohiRe+5C1we/WMD/VLmqL
PgSrA7NykRMd52oDlCQK0W4sD76IQw9hQVEk3fXjjOKNvd72pYc9p+HDSfdzvgMaGFALqccVHqKY
z6qOXOtyDIeixgOqlMmOlpHRnPjw9QIJ7bJwLk3+kD4SiJ3xPOA8oZhmTssfqbTX2DrsaJpVHZDh
YPM2OXsCMwJrV/pcHZfzrLgJnju7/8eNyfO0yM3v3ZfNyYCg5Ij66R7W4O7Ya9N9a5yjbayIO3Eg
6O79ImWjw6Mn4u+lNXOr3sRtdSbSsR6Sk6xdKr5FMDTq5OYmNQl9PmzwqK3+TdtKv32PYMMcqnSc
JWvAtuYt+aBuG0O4Kf9AUD+aV1hkO6LeqfW69UpxQoQqmnUgKN+WbfEOqUKG9FKhRp1p+h4m8m3k
933760/yPvRxSP39tksUOyzNLfpowqXUM51QzMBd9lAQgUA109/Wpz5cjBhVZlQEt4QXfIubknlU
rC0QdS+pPPYuDdt7YrxVmZMEwWRxtm9HPA3cMmkl/GzAZGgP95nrfj53w5/XAx8O7x8SE1qaB65c
VhO9wt9hB/n1NhtWNvblE1V4S7LxFydt6qNAviGXUq9lj+yPGtIxOIFpQhKSVLBP0Paj8/9WE4r2
D/eEJ6HMH1ndVMiMf4xsdL4ohIbvYBLxXgdaWb2KI5mLlZCPSMfEPJdGA8kztv0/7lvcDo78Gguq
w310lTYk7F3nU0F3Hc+kJF/i4N1GwHsk3F5dsQwYhz/13dhW4zo7WY+/tzqk6KNbH8jXfaj5sHwl
E9cwashda7bSz3SriSETUf2LuS7LhkSVwpB+TnRtpPg/HtipO7DwbOAGmbB6gKWCZXkevvT1iSvB
NsXZP24V/gEU0qlqCGIItat6f+9hyyuPpdIPF83utYduMx9QojQLDdXQSOdqR4MxZHn9j8yV/g5V
qLnnWZysl+6vHqYguLs7vCMzJ8RWk2pjrNI02Pu6RmeVUD6mshElqKG2JhzexaeYItXOSOxAhM1b
9PoKi2tH6MyRWO4aRfxXzazYI/76tXMxQIpMUuOFsTnaEn4azTPt8H4zyVvVnClYdZyz/mBdenvS
7DhW32x7vJpzpn9jKbD7682c1FaccVK+22pp1TjqndCu/5iO5AJA54rOniuroQV8oeo8Xh7UMqYc
GdCHM76qxcgM75ExHiIHFSu6IGkWFk6CkJrjiG/GDbJywscxUAabnFqOY7a+VXYeHsHtWIYJXCww
Ywl+XzdjzV+B7oipghtndtgzSDng5EyOiJU9pp09ibKYDYshd2bUGNlxEWhIp+Ak/84gxMplUMHX
akqc0ctHOi34bb7sHwDwoQ1mxS7LxM2sse/ANttseA00ibq0sne0t77KEGKrsdgJVZ9OiuPxWIq1
+HNE3Ogf7G0AC++JIU3qIyhpGFJxaeULOz8Lr89YyMtUFeeJJrFq6AMT250H+r+s4cmHMLde9j9p
eT9FWjpKl1GqzHKNMid8TbgU7YtrLuIn8CobiBUC6rcigaXmpbEuZqFJqMIaEegKmVijM9AcxTCS
YZOB1OIh6BqwTLnx67c3er6qcN4olBsxDwRVeiN+/IvuFEVES9sSSbKgjPdJkr/ZeFgc7OVxnpu/
uGGlrhOmxop83x5lQYzLmWSgSZ/tmwB4Y5sAIt8RqQOhCpL6m0goIse04uFJgz45HFjZ6JaojPhA
ZMBO7cQPlhFWD/rWhcPm+Z2T9KNM+PmdMINfKElwxjaMS+pE18vWWiEF9cao8W59FrMQ829CYza6
zc5N8suwd2fR8Au8e+Ylq3DqLz5FzXXYAbNby4x+axOnM6E69KBTTWevinYVdnXcNcldMQK1+x9C
o6K5afLhY+ptcqoKCU3uUfzdkK/uqEejSNvJR7YyBPVtv3S4/BDGEHflUAzqv8N6rXxd+GNmVI6W
UwibBJ/nylGEnSJ7dEgt1u/Tk0SvioW9gLRGzHZMFkyR8D2KUg2bk5leXS3Kvh9Ktwlwam/6psOU
IYygXpzn6w7kYg52FuL3C3KWzfX85fR8O6Rp+eTU/oZwERMeBZpmwQDdX7bDefdzAMqYlkfTNckS
HJpVgDZoclErVwGTelPNQ9REEJnMsrk6o3rGznOsBt9Fq5X0+zPEDa7Kd9ubjWfeHxM9+OYGszf7
9Uv7IKT52TFy50rcEtYaSyDiEhyzzROGKrUeBjGD5cGziH0sObDlXUyaZv2lT1g35qfiNxOfTTaY
PBaFQZCWt0ryoxP/oiwbWjIWlCiRfqREHFNT4K0prK2S5P0NG9GkELwSpFdJp2KfJVq4ddVgAd2P
b1LAn/DBEamqjNqNC+VhWrEy7+NH7eokOWVvMm4VFUPr5KwX2coQfm6l6UIoQmi3loQbNrLE5oou
pjPnLksyoY5JfiBwYniRjagc++aTELv1wa1oHWb81dFMqXaoK/vcxYkY7SBYksLJyriW6bpVyYmB
SVPax5auC6I4dIZQ1gxJt8UrjfnoF9AR8kThzdukpwMd6T9exx8godca1bu3c+h1COvccsBedMaa
ZmuPpCFJeVTm6G6hf+TLa447AjV/wjndOc+ZOR/k6PqDc6Q6umY8kGqNKBQBu7qHnRWh4UKZjphb
sVcIMvxPlXe0TmlNTHAuSXRj1g0M7vvyeqgnuzwws6F2myT2jEgw73K+yfIK85LqOTkgvDRraFmp
Nqk1oCi5RN4obXVtMYDIMuyyeBuyEonHuud5Q6nl9kmRZ4y85l8YxAUET/t94+EGxY0tDlHiSc8S
wlifDTTFMuV/SzVwSJDbDO5jOcv+xovva9UWlRJMXiDncqqJHDS4Ha8HvuJGhfXbVB6TiekhDQKB
j6ycnYXW/Jvs0AkHf8gvmsXnd9vcZ3sjLuiUjJyktPsVcx5WVTeMtJeEqt/VNwWP2lKfo7aIrqPC
K7EqFip20nW8EyNUcKC9LiCir0IfYJBYGWpFUxrYq+uhL7IIWGWTVTbiJgiNtVjfAjyfXeBa7oA1
zZ3pQuiZo6IzalaP3sECtv3aMOnida3Izj286DKC4FfpiCxUMc90ZOTphNtY1Ij+cikzNY7nT25/
vLOCIliMILY3yUm1lEBDTlFSihswOPjCNqAASR/hSJ54zSxO7T5jufmwhNlfl7AsuWK62DfnzuMU
5L5sMcOdp9kv5HmyFMqih3IuuVMr4lY1JncglXm6grqGTcSpn7w2jy5JrKne2Z+qZEs2VlQzxFdT
y6L/oLPvHzD1Tc6jRkEFRvg97z7tMQQIKVr5cRnAnAuobM/duQmxHVP7pm/zlX4E0oEJ8wQHiwwG
LeFEhuzocr0cjvj8OmpRW+u2iqwvqk5n29aa77mrm1Zro2OWDOe2YuaAqnILiD9G7+1APodrB7PP
h4p3Ivqu/zUO+gj88N4hRj+scp+jrQphq9CRanmwBJso/JGjsvyFUruZK4a8441q/ra/yawtC0IH
pwackKXLdBZXVy+NuTTwPLFos53SWweygmXfAWYTJcQ5LEbmc5Lscd7DW4QFLNdJXreFTuQ2fV4v
3WbiF2uFvSUfd0kG5IGJtp8KGkDt4cpyF3HLc+W/mgU8I1jqhdRipMvK5UXBraQdlo3x8K3sUesO
RLRFgw+I0rcYa7vWL8H0vQe6lmOc0st8eN3L93o9Y/MS5jG0f6lstBiYMNseF/XX8bfBqJPdbUcZ
bVnDtDmEtITA9zra9fZaLYzHdLQuOvjpQXWP4EsyvHCbOslcJLdYgphc0DYJpUdkuoq3vDaZfgeh
NFIdOOFdFkpazenzXZwnfHSPQerBTvUUNGX5WkiRgArR8UYx8nLNkEkfSrciLgBktMLZVSBXujmu
mW12H6BT4ii8R2xwCB5GQ7xR5I3AgavWLqnmVzr9vq40N7eBcEV7SUVH0ut0YmaM+olNEaOJIiXr
BWEqqkq3dQJaeVcWhojqXQyUT3W6BaYu3kZX2Y8SVIiNWvxK97RjnZTfufTG7WvFLVTY9fs7tX7D
Ty2ZmOWfgmXg2BmHf3GMHVH6pksa5+mEcIPqkQI6h1BAN+SwTGqT62cmkK52BfznqQ+JC2hc5krj
3vn7Y/oZesw/XyWDRKM7GEBzImPjIYY0mw4RA9HXTWJejrZ/j2XGoLnmCyqsG5f1w54KYnZ24+FM
YWF++ntl+Vsc4E3pxZLQudWThufLWWK9XFT0p7cB0Na23rOKx9DZz7ML/If/hWCOm0oUVWKHb3CM
U2Wp1CZI2G8S7Obui8usjezruoWCVccnybLMrLaFk3RbHHV1yCBd0tJh0TwoEeh1+k02Tk55Ad+D
tDJlKhmQCuSezVwktvw7QtdWe0FuIhfZgHYGQ3OGpSg02e+3vcicgYeB1iSYLzuSmdt9ojeymmdF
QP3Pms4p6hHo/sIO2YAHMpjG/V2Q73b8ojb4eYD02RkeKc7E87y6vp3S0kbFXoAlTAe/xfzvI8Yt
HByygDJThM2ggl6VlusZx6choxgUiIujYFuOS6ACQdde8RLLHvzqWxBmEH33Wxr09888fDHBy4bl
/Knatted2ksxqoC6yr9DGjkfS2eQA4IVQAzTmPZoX+ATqKXHyNv1YMSn2x6wUb5uXYW3NUSAbn4C
0r24fFzYGAvDSCFzJBdVRCEg6NZuuCbTwpumvgLYyEGMrG8vqljXs/56QkT3ZP9g63DQS/12+fdE
PnAtjv+bn+L2g8sbw+sIRvY/YQO+/dXR8Bui8Usm2igJpO/6NuKYQZa6OmHQcHDu4XeH8FlBYBMN
rmAs16o8Ic1ekgVVpyDv6QWl8IR/rcgvsxA/uRBf+W3FIdbG5QbnnTzZHOpLNKZkYdZyeXep3Zwx
TzCoOIlxo+JFUXlHfDS9w4owV2vCF7NadoGOVgpVHyyRPt12C2sFpG2B26DOuN8StWUiTCEXWuIc
gWHV7Lks3prcFZ1E5pP4zYfi3ZYdEBETnkFyPZxqWjX2QM0C5a8326PV7IQ2NT37GpIQpS5fUwGa
36wGCLicG9fyp6ZjqowepiqnQKnZhr6SxyHeLXLC24fedKvMOAB2DY3TmydcH6W08hSeTvDoS/u2
Te3tStVeNl7P4dvZGzyYl0FrHcx1bx7KzaVxKl/XvNxBiE+M+gQtPiQyBZO9+LjQCjwZ6OjuCrbs
Uo8MHzbp0IT+PiHMn+dJRz58Xz6lKcAMG4d66AjOyqFf0exnDFLdHGMeZKkFB59R4ClLYdM0gTUV
IHqoxXeXWrCIV6puWQztSSMn4P33t4kT/WiIG+NPngdYkg29jWdRtj8cYfNUzlwMCDGzgg38jWEL
47GyjUH9LjS0CurSuu+rDpfrb9QnWI/eRSaSloFACWE3nHTodY3hHrewlU6w8uvuVsL2gqqVrCrQ
qiStIKNQmApgOuxvGTd9eOhjfsQ+wUEPEb0gO3LHsZEkUachd2symUY0ukoZgh5wsGCjMnd5AE1L
0oVETZWF/VAj2sJC55UjFhiuCuB78j1w0QX2f/AR6qnzql3E+0xqy4YQsJsQN5YHCbneSB+HpCKa
LG5EWh86aXueiCzPFeOQFYQ813O4hLYNXck/+RV0d/kJkfnhdRSN6XZPNdkrvqT/R1RYu0F7MPKw
yndSSauUw7e8LKwnSroIsE4aVdP+0aZ5Eq2lgqp5kEGWWoGmWzoy7tdBCHgc76iCX6fn4GMOSfTW
rox6og5MjjMVKtroN5x5vt4a+yxkMS66cFWK4HErZ4tLxjUJudhVlWS41IYi4vK7KmTtQgy2M4qz
l3GFglTHJ5Srawl+GjnG8W4XDHDTlatp65czUVnteH+tfISiJLcsG39GFFrmaxXFDe+Hpg9a42CS
YYNsS4wJ/7/wpe9NwTHQqlvL8sk10n8uX5HE55/4LBQUXlwK8lJb+ygAN9dMh6uq5scjdzE+vL0t
VgmUYXDCXxLTeUlV+rnWHx80RDmcTl/cF1avakfEz/VlwCNMNzOaIiQRDuA+wae2U7iLJfdxdstr
YLjAEVZEikk2/KcBUdwhXkXNEmzs9dvlIQ2NF364vxNluhgtvz6fP3Qq6HchX/ptdSHpV99ylNIk
eBX/kWtbWU6+/y/YzQaVP/djJAgERgJPvJr7+HGFU5xreHojNMFMnqusCs+YREfwKpFpJsqKBM/Y
ZmmUD5UsnksK3QycX9Kmj/5EKAGtQlQlfVPSHo/+9i27R78tWavkxKVomImJdWa3b8+1t/BKfsvK
VR6vWLLfx3B+MeUdH17Hu4cKGOn4jlu9b0D9dHluzRz9mxpE6o4hirCQ8wYxmQL93OqPRaQLJxQe
//v+bmCQFzbKjeFW02DRiKSMayuK/+37Hw1a5IXu6GWS+dTkA6m0uf3qaz2h4po7CegQRutCR5BC
SdegaGCBUsSG3KlmRjISN+kytU9O1Mh+inzApXxcSZfyPE/dy8+U8u697c3gVHhKec8RYPVmso86
bMBesFNGObIXQC76WXk5j/8MDVgajsF0upl7ziudw76neUyXxTV4fDNnCs4bB0+h2Gb+MmAKQlQl
Wiq25ASJ0rPaIJMCP6h4OAPLhNpiaf0CIygbU3Rrt78OliSHYDs52kivcRl7fOYb5+DGSOMhlxex
NdDuc9iAaB1kthnd9sr3U3Uzo5cZN6UgcZYsOaPhjqCd76xrLu8VS9ekAvO+mklGFZggIfdmW0s+
ZD0y/AnAOmHRpXhfSnGw7Tx/5Av5SNSfD82fyYOcBagBdsbL9OLrYTvwi7qGUHtrnB+P7NyquS7g
BIoCK9w6nsfVktiFz71YQICV6C9Wdd6+CLQPhgCAv/cfkvxb3yDOe1NMY5AnA+HKNv81Ml8JtaSW
wcx4UNwZJPXA3T9lxys/f9TJaKUHwBL33UAw54bpef1UPlTaSSz+BQ7axu4C2k5sUOJgqDznidse
ba4bT5suUVGOjupu8gZJOOHsw1i8PDhGsM1PiisrM44wDJYbG1HBRp/gF8v25DpoYlEJYQUXI4jY
i/f5fckoi4fiz2hFlT8SJZtrJp4WgEG7nol039Z+Iqtwpp1HJEvro/EVkNGUeJd4XOE3gnqqJ8YW
83SR6N4GWbW3MEYNIMJgnCvwDOt73nC7v3Z03DAifZiBH3momnRl2jDv5Eo5WWGb19Ynt7yKQr25
Y+wNTQArFywMiZRszrTCIBpxta92Emm2IkIquPDx0JCuXE1N7cD7R5cigyBN3ZAUzZCjZ3M4ryXV
WlkQkQTwr4ZuMAu0kwlhC2sjbjDHZbIg9Ny2lcVd3BlPP7WZ1dxTkb5SZXZSGPyToioAnqEaIaF1
c4J19nlskPZ5qAEvLh3r9OO5eaIZVz9qTSIxj0Ih0MZPi3k7C6Jkmp4FhX1CBpVXyzTuDJFX1qVR
GTMkgIgV0O5SuR0cwVyvHtwXcR4b3GYWvAgwJi7Ok0MD5sc0PRntMbAvFodeHSAPLhMYED8nXQPe
HlNSfas7/jFGbpCQAHnAafRgYVBEFO3/51uN16VhBW8xyQKxiF30YHrhJSXosRz3Du1ZeP6Eooil
Hc/PWzygTSk3s8xBjdv8+cA2qMGe15rWpsu7SXIL1Ejh6KQKaPLroTpvvZf34m2klMLSSMnJwjKF
n4WBbd5UTeMN8+TcD3vPkRbTh+w028sMw50fk2mpjCFT4jsQFXg3xGno2vEw9FNkpxSjpdAkO+uX
B4ZxyfwQ3B6Pu81gbky4qqe6XOl/dRZm35TsF502PcYuOp4JpDHflxdRkQhRIEVGIP+XCJelOKtS
hv7KPpjDDVYtPKDDTyXNHkby/fqbvgQRyQ5DSAAbbU6e64LadMwGaHcJdNASergOYhRpAiCAlMLl
cslwz/4wSzuYfQVj08PZ59crLOUe/86E7YsunNmWlmy8l5hylsqVlkll8r0VL7K4QtH+eSUXDoMu
pgclVBjzoU0Z93rjidSMQxKNDe+jqZzv45/0fJNX3+XP1nLSX1vVDS8Bf4JPOgjFu4q6Ycb0uCC6
CvE3ghYGyn1AXAA4Q56GeTntPEe2geRCj8CgI7ltrHFGrCUV8VgaVKoWZ5aWvFv1y4q15WQRi7X/
lMoKlBuuKyP5BRSCEl/SE/Kd9FbuTYVSuIig9F69qyWDeFfzqJ6VWS5+2Q1/+dai3Bgz+BXC+mRM
iTNHf28sBGW5+CNynLxA/kwcQlgDQcdPvW6fFkPoe87QuEHDyMZFxv64QrJRZ5kApp98jt9f3mYx
L+d27i4HlxeYO+2IxuaU/mwygC1cnpeDyS9um2y1x9kwdPx4sFE+KL/QeHO07/hZ1NHM4Zr6/Bnb
M4Jb7l4Hv2YyDcv6rPIbIqsOTgIw75HPRIjy84fjXn7aue0tRv2VuRMnFW7Tm7MQ0zpYlNKbz5X1
Jc+JDx/dVEpIu5Fw0fX/aEIPyrHxeewulCaUviUaXbcCBTOiY0AdGOwnkRF6bmUXQ9ax9p7RGI5X
4wLvVudwH6U7vp3EiJT1b4SqTCmennaDWPp6EjyClFUEvdnpAG9DWUHOfoLJiM84IRz+kf8l7Kfq
SZhTmlLpaKtSJdidPkc7dXLcWvL+uoX47LFYJgGsjwXLgeGN5j+5RLC2JOgVlEQGr7zJumOMILje
tjpoiF3NJYX3q84O0iBdstKYdeDVKKBLa/FVw6U8reCE83Xg8B0bAUjAJEozBjz69xGDjaJsGmeI
K6eRgSVXuXtC01+rC4BTl2mvBG21H8O6ggRFtyoS6kZlGqIhuLcXDvogECwB3ueO+6ULf/K9A/fk
5EqedVWZ+jppELbImPI4CCs5rmE4h7CEDckdWBzvnSWuvZoSORN3g4sWyCTRaT5CPtdLdigPziyx
x3Yebv16KkdyCUl8NYnwFs/f9ZM7x3lxR9RzLOYuPg0HZdf/H3G1LAP1mDIlWbmarz+WNPTk0SxY
pwT1maTGOlGb51yBnTTxUaNUt9zS5PEMn6y6aYoihMYZA39ENNlwHOY7dn8VBGmwrtO6X1ehyH5P
HyMdz27wGySA/JEWeSWDn6ufNohTd0ObaG34+5ME10ah0PEfpYdsruCEIN1Q1vaP7GDzrLGEIXB0
vAg2m+7Tw/V9o5pBQ/C9n35yXhvLH22dBxMwqgFB0lKOomywshUzvjW6gDAfWLDnBlgzCW6wKyoM
0wmXvKXRVrg81h3Jptso3BDH84AgvGzCl/PosX7wF3AhVMfkiCgRzBsoJLgfzA5D6vVF3dADVK1m
5tnqqDLRHkD0YjLFWDDqm7TQw0Uaay0EuvKhpyW4nRG8+KK+gHsHfxF3C6Ywk+EroPM5Pb4ArN3J
mw6WnBoQfYsqEDecCxntDDuLzxQa/mQw8cvJ6hcCYwjpA0xvW+ZzZNYhDm56vD1Exrb8/Q4tSCd7
CpNXh/6XpCukui0x7RME+D/8QQqHSvppUERinA8e8sDVXaLS1QBuOn2Q5VGV4Mau0nKe+jBtLmx1
wluTwbtlDUxTgLbV2e6Frz2Fh7U5Yf5a/aJahNnIJdF6twtdDAcTHiFgI76RstB/UGboIQUXpA3V
tUQEgWX0Xdyl6HjrsIqaDVhgjp0OE5xoAtUQpqIYfJdCiLfcZKDdDaqHXCUywmD/C0R0+8qnesG3
ikhZ+y/ILpxJQOsb/kSoSwlCWfNLGGq5TujHGbrEz5gq2/5cZnoF/8OydaEw+IkU0nY/p5VUJDnH
IEyNWkWsRdlbgH67gGQ5GsV86CdJtR1zdGGWUuBVVDutHGJs8O13+qmVu0oKEmfMtz+VLhTuhhth
LA3aUlKzQUwwwh2qFTWNyaRCP4kpULEcERLlw51Vgxw5P9trtA5xFJOh+RvmxNSSkgpBGrZBokH7
gz2Ch3XTUfOyLeE8m3EU0ayWvnel9VG4h2WR2zItnzZPAqh2YHz6pXpdRZLS2HNdO7mwx8770QaP
QQweTkcjtXBMYJZ6D54pI5r+InyAZRkKXXpV5dBd9rjfmb+AavhkvF+LtaRzLGRlA0mZFNmvM5J2
2rSDZeNoeMgZ351Nh/z2w1Fo9irriyf+7Vy2ODhx4rJUe6BgTz02AbVrHbzzs9nabvQaZcZ/OoST
PBF4punlWJnGXOYPQnTItq6rQrXbGAqWG0FuNKNoKzyTjgOCOy+tCY6/wkP+gUrDFkR2I6bTK55i
NysOzp+2WxXh7Vujjp16omFsmVlp1wdonSIimoKH+tQfGN+i2IHaHfuTwXlHq4+u9XhXkk8Frt8Q
F6Yht10xc7OQEqoJ+xM/WLhu2D/O7+2mYnqwcyqdkf10oep/maHdEBc9s4YWGS/XGl/CgNNxEA+q
SCphc1wtyCWJZ00uw73vzUPv6OGkbL/Ma7sPhlh1LE7KRh9k8vSRDdk4aZpTPSq2TtSKbneg5Lgu
94pgKwAjWyhmclLBD17nMVYnAwZbCYJZO9NWeyKJ4+Blc6Fd9Zlq/MBc69xEY1O9Nisw670D7wZp
yedd4S1hkw8ZFmta31AHgPqJpzG0FqIcATqRt7MM/h2jijzOyzT2gMGAtrKOAHQn0XUPeUwUgmr6
bLPHpIjNln14rKd5mUqkXHBoMph93Cc7zrm8lvc5iOUQrHHrAJLFECKHbnBugsQjOnilXWt+z4IL
U0PRfDS8qz1bGi8Dl2YzySur7Y/oE4CdE/U0tmCUJSl7Nnqr/X03KTxaVxh6tntZHq7dT+tCEw8n
Yg/rDuCch96//Icn+XSEKjy7uHPoKs99t3YcWeZ98bieAVN0U6jjC0+BqO5wGHOo4zfZmCpeazST
9hFl/JEQF0ZKr3hjzjfEaJBfGX5S76RvAqclvqyug1aR2sE8dUoxiJImBQRTJnUvxUuopeXcx/8A
EhEAhCOAPqQ/cDL4OpUK4hJLUn/1otfHYrwp5wjcHE48W1qKk/48BuEsRD9IaJBgQwd6ywHhXjYE
xVOqU4s1ko7jOckIfVbesMHzJOQWGb1zWgOP5R1lJrS8tadVEYKHAxkPB9g0+8PHwKglGVuAU8US
RS5PMviE+A4e1CeNwgrYX56uTb68eQBh1QxDtu9FscPYU2m2NZdjltbyFl7cQuRxz/8F9dRd5xtI
Plb3G+jJatqE15gt4I8qioolREYhxCTGFKFkMdSknbjAeXLF0nxJgKtOaz5BAL68vdUjBWdqBGbA
IuNeRb9QJic0xu2MUYTOHeKdHKqR1vB6gsGqq2UkfgnzUqlPKJAa+FQrpA8bxrwJDx1OkcgBcqss
ylG9IJxWnKWaI1BH5hvbGpQbsKF3X+rrbC+pCpZCmn4ZOKPC9KF0Rd0elaHK1Buhm99I9r0/ZD10
rnv+jsKtbrfnCqmQSTLW+vcqRLfNj+ojKYaMQb+cZ0KXxvJW9cvt+dLDvfBqdTnuHhdCaL2URVOh
rSj03vQnYujA0YwYX7EaRHlr2wBTkva7BWS9wx/EsMuA+knYA73qUN2u26jPTpklOzYkl18nKWeO
4UL3nRq7TTb1eBl1I3qKr27UDgIh0Yi4+Oj4jNgNtqikc3ckx4gufRT8fza5495Pcm9gWJhdUAki
ruLPgZCx+BUpSERa/oyDSGy/RUYFBLiMYlqKrElNCjyathQHWcd54pO8CF/JAVAu9l3tloIU4M9V
JOU1mgjiy+jAmQY5lR9NNzPIOlZPk7zLHMX2qY+Q+2g5MYDTvhCjPok62yzN9sznSJhBCpusCDoh
ibr1v75R/DIguDEaeJ9fbQEpf/JeXIY5fo1GcgG/RjS8CO6OrPAC0sKKkmCystoEGsQLUNbeXA3c
YT/QlMYoc7T/Bd53dadue7jYydHr3B23iCwPfl1cTpDQgWLkwOSLVGiC3BljQsUzNTy86q9rxkaH
yqjcMj0pGDJ8XJtnqHfiJ/aOOPmeb+9pK7mOnvYTJKESJJuKaODLhrZlOgncoITb6CyeYaFK+ZBc
XYqxc0qURYybu+vBZMiZ2jyvqoORtAFTWtjyCC/Lqy6EIHcB9jvbjcErvrfjz4d4JUtHLspPQj77
Ap8cozYQzQ5LLiIaiH/v99z7C7wcrTdRFt0Z3/ZfaT4ST1LsL2ZzjwGb4Zy5NKL7+bHUZnaoKpou
Ji6cXVJmPvOgVSou9aN/wrlerJHCq8HiP/l/0BdNNy6B30yW25SusC63P6yJfREjVvaP34h6Abmd
9WUARUJ4QKStkU8y04aNcL+91scQVLAvX47+zPnkMUF7kqmQuAcUKPnRJ0dVIRp8BmrP+kKy03lH
66XtuUygaHE1s3KIoqaUdd3Yjagy0ktdKNmgiUJzd64Jeb3ASQ9RxFaaU0iG6v0hjhAjC2xg7QTj
tuPbH3j36Oj+sAvIM8hUflLWGTRMO6OjrA5WijPxHPRbA3u9oumhkLFq1s/o4o1Ke6dCBsMtedm/
tqOXbanQeSt4EYP3kIWFlYWG7zXg/qnRglaAcSvUHTRTjQRy6B8dRqYFqjPk1NvIB5ESReJM3Wax
kFxOTxmHinjpmY82hp4kYV89kfxEuYuvUL8+DB8ZuWoH+ubg9S8+I4XJ2NYvDO0q9PuxuG5fPnOe
8UmKRVEyOMIq8LuhtiiDvF0oHDhgUWPL8BaVX+02mx9Q43N+cjF5SlugDJpE/dUdk4QNTXWqLi91
Zduy1NlbFAcAKfyhSQ4p9LWaO9VXeerCOfUpbcgP4YLa2XjfgEdSaFeZA7pVcBC/ygtMt2K5g60D
NsHSiiyO/zWtIr/JGid15Hiytr6TZsSRUP4iTLTRRAM3K2O8tArTqIUoQC6+79U/U4TNlNjduABr
YQXTOtvRiOB7tBTVYYDlG1KEm+6aOo2/J6hrnLMzW+Q5a4cUewgTcR6+IuzveHPhoDBkQ4iUYD0D
SHAh6pfaU/M67UnL0MJzq0YnkCEeemU3IXAjQIV4oZdcrFNHmHQQqrDm/978j+FdndbuRMiAmN9q
lh/Yhw2x+BqspDxh/gEeqhuytWK29fQTagJohF3/sMQtNlhbdsw6gBdFLCGESeYoAMYeLYpVz85G
nzDYfy+TPAqdctyoPZmt1VttrXywYnHUPsnojBG6O4zz7Wl/xi0ii/LGxVFP7WkvLLT3eivuDimO
1Nk8BAgfvzO4biW69J7CFotirPHZ5YtM5mHXTiq7NXjmN/qpbl6okVdMWz2lc6iRPJZrGTE2YCmR
sK/sN9qElS+czXqfAZXZ9fHulJIIIfEagU3AXFHNfwfeTOy1Rd6+WulzCwqJwnQsRVhgakOAeaQz
Y9SJQkDceqpTfgP3yz2ySE00EFw5CWlH/KOjR5weow4780tHluX+CPHUe/MBD+gXZzluU2lk2Rdf
iw/aZfKbyaGV4BxF7pPJ0llY6cLJHmVsRnewnoCLey9iyI/ePZWYdiNWUPvGH6Wb1G/4y9tcy7qu
c99BFk4+gnhLo/yqLmNjOr2TLkoVZPR9ReAT48DqDLSVs319WuCs13FP0B9EYXiYqX4XYbOmmquU
Ui/9BJK4E7w2wBaZeVXOajFIIUejh9ZJ1m+tn6AeXyRjwJ+1qZQ6gBNOCq/rKsatAdKNG1stgLH/
Hw3XCKgFYi7ego+07iXA7ufVFG3FUL7lLiXLQtg2x5/8a/n2aZhT7F1HlcbwT3kzTiYUhZy9rmY4
mbPuxdhRt2hreWm+cD0Ayto+sUpJs8tjIe9LuVMNDgN1ROIA/u8CfWIr04F0/+LFBQtye7bTCym3
qrElEmva3VbfOzi83P0CPVfQssGolYL8gz7YRfPkiXcO6PoHtk8rLqZPjFJ+bkkf7CUq+pN3r1oT
2jsdk+pRaKahoVdVQNH5bRsjYGjhsUla5uKbDm3kkuA6s677I7zFIbqEYhWnBqd7IYQCNmmy0PrT
HQ0CQ3v0HOdVLY0p8WC+E+YCLUQgycrGBSABd0otLFL+BI//qx6RKg0kZ8MAleXWEP0T0tNBF0Yq
4uzRwm8Xmp7+2Mm6gK6qPfufximfU3/Ykoii81pYMEIP9j8kIxKL1paQ2zD2JNAXHuDLl0i0p8By
yItfGKC4VUQUpKOiMqzBXeWtwlhUy2DYkOJ8yPpm+IGkNzQe9Z4dJvCzhX0cu9XluFBERZMb61V+
vcSJVrOD/9TSqZxvN/evm09IXNM2Kt/3fs+B+AcG/B8hD8fm+zMM0WGnRFWcivihThtbOeC4yDYw
YB6t1msuJO1VA9+cJJoxnNFx0Bg0TYoInBNawPgMHpNHAStExtNibP64IhJippAsYwzC7j2yLx4x
KDHYgPZdHlzucX5PicxsEQ/mJwI1qij4wWLs6CGL3EAF2bSZpl0hKmXu6CygDh5RZwHs2x7jrlKK
LKByqfD10oh6Vq6OxAXf6goqVyoLH2sdYLQzp6ncH2/BoYY8vdDgra+1n+YUgV0vZi/zQyrIU4Gk
ogX7RduX3ozc6+bZvIkufzMkWcBYHxTtsTRd5yRxNFXDS1GaR4RRQ8w5h2V9IktrhPrD/+Aden1Q
U2BcBvacmPUEwss5ZE0QIgZrgSfkBvhcFprdvdz4pd6ZqVCbnIU+v+jLOlB1onBXJI0iYxFm1hKR
nGUeyvCygGD6DgI+JtXMIsCIe8YeGgakvMj8PiuzJ7f9aTtjO+R08fEKDgnGbWDME0sslfMUdN9A
6nSglRfVEB/7t6aRpSL7izbhgSzkrZ+1JKLyNrbL+KaqXwpgXClwrnctkxgqf5UNU2J5IOintnz9
15ue4cOTx1p5Hj9SF3s3z/bEWWvCnixpSMlLzfxr2vrWu4F2xRLRkSWlUVGJMNJvSMgXEjAPzLSH
x66Mx46J3gmzezXCOyU/sDix613PIK/J2xG543IORI6QdEfh65K2Q1X7BrhzmmIIXWooTUdIQ70K
MQskIebBEPWihN+TdYs1SuDf4/4fHH/mKm8hokRiqmhgbNGdOmxuJiNYXaGDdIEB5icB4/t6fbVM
cceq2rvmDjX9fPU/4K48WK68GeXC9LT+yWfmL7aad0YiiIvcmBrKJ1koEUKOZJ4cDDWxXMHKWf3p
GqsZqWg/JHyt2dvcET2SZcaEViVWXqVvUweAzQ21D2xZi4lRqcJmqNgnfqkKf3MWQNvyEBu8YcAA
/NZaR96hb+pCyhwAapMasleCiMxRpDeIUS9p1L5CpYgm8C/5J+/uVjuvSkJTn5y003kOsI+b6MuW
EKi2sUvvUi1ZC2dxOOTBgYrvwPgPF3uBLaKjRp6TmTVu+E8/xnEuNzV88vUMaf6eDnRggskcioZ7
jnB4GRtzjRf9qSuKAgmOyh+PUqgBc96EB4dhTTKqEYaMYYFCH4xlF/L/LZejgfH3gPGn0o7djMfW
SBOgZ+aHPkfBHpZK8DvhMBz/ZUbed+eCo4qgClAp5vLaTvi87k6KuOlHxBkcdYmO/sp6dyyN7dQu
94y3ZUffa1Iw62M/OYPMGe9TvRFdm/4FIrK8fYhC5L2ywPH+RU3w2xSG7fmdvBkM3ifGnlq9jCSn
z0Bh3RYnf/fUKPNUlDiFkcyuplp0ee/Y4g3Acyz3nx6BVieGISthidYhbs4bmCl2qOK40BAJFw6c
VnktopVhjVRzdN0KHafWK5MPzhe87bYCb/EPv5BT0AI9Z9nahkBDIIfQvRyL5HQhQZVt6ENJBcz6
AzsNRVDyhQTgRrXDs4gttZBmCj1VxWcybGfwD+gyGCkUqDU5w6H6oyHZ0vx2Xpdo6K5QhqdY98gb
OnhxIroPfmBzHnAaFSmoR369TvrPwmIX1Q5kg19PYajrMSUx1Ui3Qmra3TCeXk3/fIG1UpdpVE9j
Mmi5JCBlM9HgjJw6hCf7CVRW8XIEMEXAPiChnsKlc7jZNLLRrFjmkEX7lerVAeAKDmwTKk4xoXld
0iUCgEswYwQbNVxN80KWKZMcx6IcH4rJYH49BiBkK0t9Kp7UcCojTe6REcIcjy7It4T5/77s+vaO
YYX/jiYbJOSMEI7TMvFYWMLADcgIJxsQGyTf/i6YF4XHc+vgMT7fKYRKjFeQtx20NnlOP1kJzeHt
gAH5Qb/1vxIj+Dpvw+j+7KkXVuDeJz2jvFcNrD/HXxE16tqCph0xzkor901+/4wlBksPMBgGhdcI
xiREqHtsi9qp1AHtWdd04cF38kokZRfPHfcUKw8iexnWTAme5gGCMaBHhLwEPNQa1e/QuEqNFHGD
U4y9BNTD60Owo0hKf1aoSakWY3qtiIaymDwa0Q54jAWv52FYeIENMrHrOqMIxcG/bCJhmxHr2gLb
FHRM7HEC2QCTAZna2x1hyXedMGTA9wTytJoPz/klTKz9cy+5vvl9MaOLm25ozdTVOa3rIGaK39cr
QiUWhgMt0vPJsfK0si/upnni3OIq7RFgTVnftqfhHKGoqbx4d0FOA4z7TuEfuLyUB5oyN4eaH9k/
ORPoAOIHBERJw7UZwBAFdP9vPcIryB600JtWRAI37lCXKGMdLCghlYI8z6zk20VlKE4Z6eJBuHU2
ewCb2827EQSCv+p2HX24UsPBEhWz2B1+WsOL4vUTIRlFxdlQvQor1EMBfkKXi8YniDmiIzqsDCX9
0EWwFS6LD6pUwwLOYuTr5XuaE71qTNpIeF6C0olBFA1L/oMaAi4znOZyA1guuIbtW13CALwtTY6R
5Vcyr58VB6U40XCMpZ40S3/mXbuvlnc3Sb1woZRA9wxjnIWoDukEU382f4POu4yBoJXlWZivhPjN
6EqJ1QCOf10nONls53vR4cQgBHcmdL5+07q+pVASXsTcrALQg9wBYXy9IRzEsnmQPor0zQYG6sh7
mmh8a+161kD1HlABDSUw67wdYFUYyIMupuEt/dhdNSXKh0LPukisMPrjlS9NaDdhJrSyH9pou2fk
ZgVjCRm+Ore2itYDOkrIpOxiJt3M8TIYY9JQ5TfJYV3rP5YlQT5e8nJZOajNtphAzjH3GMQ8D6Ks
Bp3e6qVGdV5N3DvbTT4+2F4q/JlI79TITBt9CQ5/9e3b6QW5pDpCLg1n1Osd40ko8ls123FeSlZ5
FN0GiRj9QRFZF1llQsnwdMNurEFMmn9pOGhFlM4X540OJdb7LyksOz4ovnnIEni0ESOJMzxWEiDy
ROkzd+/QPOb1mHvqcT262dAb95InsnjErQmpB6448y3EPVJqvHgV43ggsIe4Eb+wpyy4z+s/jvXB
XVorFujpaBbalnOUveOUEejaUVZuzu0g+81bcmtnUNzk3UlWN1/V4g9sXEccoCB24X5WHU/EhIdY
e0+JLvCNrkS6bwOqtOSWSDMAydxY1xyQdJ9Uf7FLCxk4t3lgf0J1uD/XyJz0AYExH2BBvTZo+GYN
C6OldQ4jImPP2RvaVsVIO8fn3At3TVNTko3niOEnxRN/UxCGIeJYOC7Vya+oDXo5l10jhs0101Rb
LJjJB2atZnp/UvqzGSXih0Rc8v8iUMOQhyYgsVEh0MAdzg7gCw/3NQDAyt4ivsW1vQdC4L38Gksg
sGmkiw/qlHR3us5IX4BeDGwkJJM+FzfQQzU2U2Kb4OcJ4z8ik239c4yBV1hUQZfnvrsjeNS+m2Ww
O8Rw7CTLc1Yk9NhI7sZeElWxwoLMdi47t56jNuY4oUHxa0nA8d05NVDSabaXyj2B9XtMbeWRQakz
JXQSJt6Mcdxy0vKmvxNgeYr1TAtxGmWWJD1ammfUPJsgmEKNi/cSpjfH2cqhCEskWvc01RCWDcLI
h7MoymBdfHnZNxxmsjatXPLqmeM3uT0kF3doJtKOYQeA9qIRSIi5w414H6u85IygsCX6+W73aUJg
g/miWvbaFfKoEv8Wf2rqUAUUk9JcS3Wd6q4d9sN5ZQ/oIpqkEUAOLQu3tCCWbacp/Jui9u0MyHZE
7bx3qN1RnJonyoQOZpGls5Nd7OXg2WA5q2EiErO5vx/dfXVNh2A6T/XLoQcF2xLAzhwV4KCeFcqe
2GD1zLUJnCk7jWadOG/uGTtWQyXEuf+jb4FaHKEWDoZ5OpNlQmz2eyPssjPEESjA5I2bvJxhFLZt
zel9sreDBXnEHc+Q4brVLkKPDLZ9hNoJQIKcEE+YTLlEzgH0jdd5ue7j7Gkfgtf04pFdp2Ob4/GB
RxJ9LbEU0zngYcQcen6iJpQ7+AfJPV51PFcXqwjOp+RPvvceZSlcrvTiirdGpM6qgQzGvG0FPbhn
QPq1qP8Jl+BmblASL4YiSkqDkyR0BK69GWUhgI7Gs8mhaqcQNNJZbk61+RCyFyN4k3Lbv2rwC8Sr
XOs8l88cbFnr76YXls23zuMuS2N2R/3gom/UUYnDdOhXBM2op39c+tAYMbbaotPYqtwn1OAE90dJ
0n3iC/gaINl0iC3uDk7Jj2sbrq8lka+vxuJzRhvfy6ZfDWjaWb5v9GJeNgUflfev9216NGlE0oDo
1j6bMPU/T/Cph07s3H4adbEbCMNEJpCa48/bkHI29WJ6oiXfPPoK6TjO6J2rOwJt1nWLUZbxVpKl
IGvU8mH2CTF/QMSiCWZDEkUSbVHlTH6P1LUAQAEIwRIYGhfOKNLqeTV16BiHl4o3VKLK/FAqJBCQ
vJ4fBGTKJtOngAxn2RG7oUapw9w/PeQh6RCRaJd3rBlzm9DZaphWaScER0UhlwZsTNHryaODQJ8T
ws/G0TYWvZBm3iHXN1E3kAy0jLdre8D3kNruT/n+xrdU0/KQPxhX7mkk+dvX1bXrdIGikHIHlhF8
Qwxu0vCO7WXvtOVvj3mxuVQY3i3w99kaxQFEyp2DlHbrAbDPqoz2Ws0o/FgyVns0oPNLxvmTtwca
fmpHJfV2hB+4kb1OEXrMFDrWM3pCX5D9RVMBqmFH8A4FZWumRDsECl9qPqTjCuNU61QTWmwOhjh5
C2sqAnQmndRz2E8nHNS/M4xxKKmI89crEECyiEB1Dy3GXSGRNeBINw2ZZQARL+x1Krk+oTTSNW7e
ed7CeQC5wzjDjZWvdtnDPt/TY0nRazRQPnvSPTY59bnstt32FSMGVpd/JKOPVIsJvJ2XtJvcXFd/
UYYRyToHNUE7ySPV/WGqptlxI/Y6nVFYugfCBfaRDHWMdg93Wg2Qw7MQJOoCrmYMK3pwbHpCp0OD
XMKg7nUQsBVc4xQ7QqJczAkKP4t7fwRUMWRzD156PoDrlMP2CsOFDUdARk4f2Ws1Il6Slgoyfwr9
RyK02x9KmtVx3iWuofLls5k94lobjqiZ72gcbr7eJouFPBbJOLsk96P4K9PdRk0i/DKI71I2ZbGi
IdTyQgy2wTM2rWiIERRwG3Hf/qBOZE6Gxs7rvS+gLBz5+/ju6CWETn16h5Hq8KpCrT5YAJWUI+4e
GKCNEveNyOCZCIU9GgwE3QKnVEeJYorKSweqtkPrrjPDvNSLNKKF1EBw7umcakiDz9eQPviS5S9V
8fgRqhSCFgNJTmt/0DpSW9fxAmiobIaQQbMJcSqAJcrMg1hiuGCPUNaRGNmZx9JHY3+J4EkD2XPm
Q1Jctwb9LlSXNDR4EnyHzcaxV9YnSQuxh5yKRvFqtCe6iD0gCqokkehoL/Nj3f+ED1P9S3+/Dksw
3hD67z7yYwqoEuxzFHuSNYaTYsa5VDwvo/ZfUuQ8MHwqydUYUlsZE6EQq9loZB3BiDncRGyNCYXC
akw7psOZRhDA8HysbwZtQRD+axy2Sgmdb978V/B/jTFpPL19KlHaYMkm7J8CpJqSZH4XyaivlOe0
nkdvpxwdSHKnH8Wqa2W94ytfZiiL4/ttbQMz+KLhme6Rz4utRbJNlYN+fquWULqdp3johc5+p6jb
6XA8Rcjg5gWorcavmwDcJ6og3cTI4D88P35uPLlAhmvdMdniroFu8awAjxfQl0w6eTscRZfQM6TJ
lKHadsdFyP3priJzHjS62knQP/5pdFmMatnJU2UPYxb4qzCsuImIJXwKeUWDs6DsIDIqEG8yIyCV
74Qmm9duTM4eqa4oarryvhBmWKyv04p4ONcgD43TR3bh+Zan+jpvSFmM4hyMR0jp2xKP8oHjfZgt
CYWP2f9uWNf/1lXaeKOC+Nh0lXPQn2PpHMxVz1pm3A6dCtF5U00x47a8NTV2asWDva4wMreSV6/w
NUKMcA9Uy7/gSbcUzAE8cc0IZ6V3Ma2o86wIkUsHRrDzNdKhYohBJ31YXi816MRCHYLE1o//skio
nkjgfoth1fwie6nAovkg34QbUE6PNr6N5UASGieiDVVFm6sTjLXT4HGHqtS1iwr55tvn0ueLwggp
+RqhnXAN/klh8UvTBv0L9MoxkHJrvwYGbn8bQGV3/9LMqgdQ3GweO4rIFZSNohmQQ0XrTkUoX57d
mJqZK1FdrcAzoZ4zG2AWiu2VzvVhSeajL7qKrdMNBlrHwhRKD4uvi6Sde+oB0TAXpIP3Ybusqwr5
hTMD47K+wgwcBJGQBUjHo9mtjUXIg1wwaxV8lB2Ank4QFBkn1ojbhkTx5HPpve/Y9RtLVEc1lzAu
PnRy5Re/NWkmP5DBj3YumllgdtrYmyekXVyul866wHskkh+LhSqi/fi6wkrFC2csxl+f0STQrMQI
sCNWm2ZkZaP1/VFS3D6RfYUApyHYuxl6yLSr7BZ09lXelllrppUSjtTbuHnexSxwXqiqEZivlIuM
cX06p4vl5a/Kc/QKt6444OUh5nBGzVs/Wen0PexClblz7opAQzDw7P5taBXFJi1xIOJyXqY5Agis
TDAe+rTkTzJQpdmqvIOhtDGEnJLTNq57YNAkzp7KQrmSewOFxfFb8DgPbrlIT+qwfVYmaaeN0X5U
7cTQLFta4T4VNTfthsCM1DPyzI9+eGowtMpJLKyg4IT7xxmuLuJK8Yg6voc9OKUsskeOlSj7dbVm
WBoCB9+8+Uy41A+K1O1WLuVGQsVIFUX+4ZGZ8SXqiwR8mimgK2qJ2M8PTiurDamm/lL3a7wQXuE8
FJHhOW+gMQPtCC/b/KWXl0iiaCKHvwxl4mDQ0mlR4vW+sLMM0L4eqbpaG7UoHH/5pKQjUTGFnAaa
PJbywcOEXmTY52EdbRf+BYYVV4pxcMmgPM5XgzAI6nGr977UnTxrsOHHTIlDA08i+bV7yDp+7+oC
UFZiU2HOeR5DcXnGoqEV9IQ5mG9kZjx6gvHkX70v5XF4yr1Lhl9S+Rx1ftXC8MvrTLymZTncIsNh
19vlFJbsA7ojr9pypWTq33PAXJqdBKwOmkeWiUNNY6ba38aPV3EoYjmeRC6zZ4T7JcJiB4+gH3OY
G05N/xxkSGg9cCqnl0Q4Gll5CREEV7tV7wZdum5dyySMHWxb4GYmUFebhoa36NfwEYXGHw4dOj3J
4OnZ0z+BTkSF68IGypgxA5UfEWCzI9bRTORujE49EcCYJbP5QiEPmHXKV7zvdjG7ZIisWAmsjxJ2
cVnBkvTriGgovKL92DQbEsrray0wUNkuJfkFFLNd+MX7H6utNNJnw/9yUfXLrjJxGFPEvucchRYr
UgOHXAXZpLrz6jU5lX1m8nhtaj/n+K3HrzuukwBU/5ooqZ2hG4Dx99GM1YrDTrklhRo5ShT3Yz3E
Mse3B1PwtX7OCWrWuWmvifdq4KaLI7c/orqdGQ7XYVX2MEiUSjkRCvNO+7u4TmL2OIyj06A2b9f0
VHiTN4ZqHS3QMzta/JVR18R7c5bWaxI859zzDF5dVErU7bF9DeSoo6AZ23rtfGmgERpo95ANVMFo
azl3T9WC/PkdHL32hlhNZFys9SrOQfET6fbh99KEAcSIPBiQ6h9n8hHoFAQUFVDLtwFnKWtf50ib
UmjWDpl3mZURN2viXkOM1uaI+A6y70570wjx/HGh9T4PhhR1K26LPH8HAxKbdVQmFpeIsREXNDPT
CyMq+DvfLU/JSglxEYPVxrdJcrQ9x86/BlVFwFWv0uviP8+RITR/rbOz9N9N2bEXpmwl5qTqfNPx
t+lfS/CE9pOvDdwLL22N0oI69b7vVouuPUiT11tqU+TTZM+hmlyPXwSG+2+VoUyLCyGzV0q7BXdg
c67pd3nQBbO9+W2wDXDBM+m1nIprAhn6aCo6vVB5UxT7KYDph2XEdHnV9EYhC09C9BWeVHJU3Jyq
0drg9YvjbdZuwycZ92/lROzDrZtnfZr49eWwsQ7Wkyx1joaXcqwvkjpwMY3Tjpl/p2oFeNmNjELT
gdgLGDRL75oHZOB4vUeWkMQCe4jVvPr8ZFPoOncJb4SpJVpsmITBTVO8kVjrxVJS2ZMKlcb+DgIq
7/XRbSpv1Y+804GuoAOyertzL0lpt7H/5H6yFrGCscWGaL5dJfA3la2+lxWYSHIZUFDiUFopRC0x
josA1hxqmNIOM8L8g/ZOD6edFMWh4UmkW0KyBXUNj7nhGDhwkceeyIiuV1TF9iUJUp6KJXUdNhIj
E3pbYys3+4NdpY01v0v08CvXi8q62uPrSf3Z+icoQN7Dl6tgbvhnL/HjNosPVDqRe0g45L7o9RLs
wfN/LH0zjOc0MEFahzU4TLwGR3N5upr0FQMN8T+hfmnElPzr3EsdQXrlrdIO+uyWWFNaykgZhAUT
BMIZw1msRFwssj0O1W9Bn4S0T8IlbiH6+hVD87itcr572fR3xM9sg8DcHZGhjbLlpoFLhK9VxdOA
LJD4Hrc1M7r6qFmPVvPVfo3LmaR7i+lxqhFP9TNOuRntmUcMjNX+LFt5Zqq6EmHnDDJ+n77+W2mX
zu5jf5HdDOk2MNCdmcRvmcjXIW/nY4g8k7y2uqjMvMguNGUaOU99CxZh+cXo3FUbkaB8P1/QGw5L
stJhq7FzDsAiYQ0r3ThZGyJn+bIaKym/EEYk58UReudxDy0F+hkTq17JTvSL60Ig1V2Ba6MsMpV+
qioY6h118KGVogIyW9y1uTbYQ/fhIPgM1SABvgQd5EAJYhrJeWEPqsuh5JIHxHyl1MSYmexUAhwG
3tOzS15n67iht9xH3bjspQ2/TnZRHFHiH4pId3zLG6A3OQPK6VRSvPgZ009c8cb9qn0Xw9CPplrs
5Uvc9aRSciDfczj1bAJx/EbvU0VS8qvtbVOwIbmG6/ZK9L1FO/TgPTaiLtvK60dJDJ2AtGst5OTR
dOQZ65/gEXZaiyBqnWaHFm0Lik3ZfP0KCav5VLr54GgmS89dCpyfBiC/5vEAWfBWDS4/qPqVNmVI
owo9YAjzzjaR6OkclvdH3Rz1R4UP3MpG72TK2jSxjdQp+Y4ZenObAPdfYfKvsuDV5Vtu1Eq/Nyh7
CdjXrT3nciI8OAUY+BKGgP2N2Klpv3ZgQczxY7y8kpH4mfR57+j9icELt9S3xZ/tKjFe7U5F5C6J
uuWjUNWHq3/6WqZmVFz1BwWfLy+iH4Svp0RZQAQJxwpi3fUG7UkW93aP9186osq3Sh0m0n8ZqXoM
B4mNe2Wlutccfmu8I1gLbF0Xt0J2J2s8ct/MjyP91xypA1lqJKBkllccHw+2M7Y9yxdnmWnea9rF
Jl4ZJXxEvSIkfwKEZzav1dQe73N9KgkXMM9mnA+QlMqgnWN7kTwfffK1T5INfSZnmTzHIfLfNRpZ
L9v6YUOVJ+xQl/jpaTusZjFcx/P7oW5Gr55m4zBZtQKY1E9MiqITGwI9XTX2wdidktY5+36bG/7G
xtAGul/1eV5PWhzjAa5a/RecFbqktz9fiY4W3zCP0OLcEDtETMImCGgHioN5jiiWHcqgjEqUKIBL
JCW3XmmaDqM8lfPUzJWUaEWHasIjHuApCdqCya0WlJ6RIPYUYr7Gw0TBnlh2JRfRzwigybaB4QKd
EvnztSBjrP87BwuhNZP4Tr5FR9wQ+GBMgoL9IFHssUNMUR5ZmXfZQ+bBcrZSZe6Gp6QpjaON2+hY
xDSGg0Ex9ZiJFr9f3QplszPnp4IzWLyNofa0iPfgcM0Jxk+6+cD26xbC1awAcswb2yBlraDAvskv
1H3fRM7D6MFIT8A60YF7J5dz80Ylpp68Lz0YHEBqt0eh4XhafuvFfeoBtHYQ/Dy8IQyavLtslx0l
vuH/H7xhCXLj+nFErHaDwdxyBH9s9rxJ6OJb3JgaVrcJ7R9SxpwkJG3eFzPhw8XIjlvrA29VXT1s
5JRuUda5LHPhv7xa9vNY7CdqKFWBON1Od5EdnGkYcaGHs1L59hkZAIyQ+EFLjwv62IwpUqb4DMSs
AHJShsk+hXNpmZ1IuTYSVf7wgMJNz35qJGLLY9KgWmfT56VdAqwkz5uUtGO65IAQ3SKz6Up39ekE
sTh/x/I/IYzuD65xsE0Ru7q9REGvg7mJVjspKUl/AeO+dmmrNZ3mYhpS1GobylyNW/BHM1MoU84q
oqtPmjZhC0CkgL8NkncAdcT3Ah0pNCCLDGm2SbaUYONJ8oTL17t/5s3wKdA+fNXlRN4mjLVxg6Ds
stLYp0KZOeMRz74xIfY9koRBiSf+OboQiybN6C7t+KOSRLDwhbRcr0v2QtjgWat7AND7ztkRn75E
EBBYmpejOFXSaFt6ePBu5fYcKgC2m9NefD4HA4j44m4WpRa8n1ovW3i6Q63ycJ+qDzpgOC6PuXIo
I97gyTEeq4sVtH4ovvusZxEOIu4sgaZY3lrSYexVsOLZW/4LU6BNALdTjDmGFEkk71VbtQXssGNa
CyNj7MEfbhLve0EOl0xtpBV4F3TTsnFQpKs1qcimcm4tnR/WRWj68w7u7qookXSbSatlSEttDv/V
jKIiTI+aRa8H8S2VedsdlMptvNzJ14m/bhMsZCo+dKH57CZoDXC/UK2zxl9JeiQ0ct8ubwN8G5v0
3V5JBbQeO11HPl/MGVVyFtdU6N/djB3BnvXYX/hR+YZlY951JTqw6p78Kh0kWxTd4v7P/NC8e7ju
QOq4rs3iqZmGRPDueSKB4iOXcmUhvJYk7mrSt1C7YOfDAeP7QeDe+bU4rJD05CD2oOZcFUPNaKfq
9Vu0mhxxeqj4AjbvFg/YM/bPyJK0AFKSEBQk4chuQlAFOvMyNcTpPPqOgCm4/Q6TOrQ8yi4E1lBG
1AV0gMYPIMmuWsZ0IioGUfKf629W0jgM4mHUf9dU0/GUV4CYqwMAhgMWv9aYFOwvxXttyO1VUKoz
sIFLDZZ7UTALpNJ3G/Fx0w5QpOBq94mSEKnnSleoN79i9spHTeCa8kJHIuN/hxu5x5AKhtJhZ1Ng
zLDH94itCkyREzd8YURA4ONFhIk3IsD6wjSV6AUGVt0351ncIkqKTqTCY/JnEefHEqE4fczFWUj0
m5IKuvFqnTdCgXgWZa/4stI7PHEzOXc6ebHnfkeZyaJlUef2TyKo4yqAzchmbB/hLqPoFwpDa0b7
xbPYH2YjgGEYMJ0KVC7L62g7RV+w86w1TbdEavES/H5xiFnhwFEafkaxgYgvMfcsgWRYDKqHiYdz
gmzzJRDWW4luc8YrfeIoqGJXqSAmeO1bq98lCEKhNWg2p3zHyuB2Uk78G1mQycumzyV2JtrDbUk6
BVmzBhQbEDXJI7Wjh5BLW4gaPzvlhFoKihKXQ9rRxE7qFrr9Nv14tqKS+pvcuAe7SjuAbDLNbMat
xk2I4Gc/0JJTik4U8d6Wv8pPEcVNU202M6PM+6JtwoeagHQmzIweyJWn7yzjOk84oZ1oe4QpQHHN
GGfKjOdY3+CcHWimXVp7cBDvtQUNSXu60rBWA/PSXZJdoloRRVweTJ68aCZitfzZ2T04/YcXAsNi
pJ+irigzM3B1FjSuGDf5fyCOtPrmnuoh2cb6tUxclV3Yl3PbQLAPIpzRKlRLW6rLnIYT7jQqhZPS
zx99DPbqdoC/omjDGRCEbyGBL6cqL1oXrocm/QYdJ9vsMH7gHfcswWCl/pQhSs7ueYGdLwZdmedj
9gpUi+iMH6eBn9gIMmi5xboaxOfC0LnW/JiE76T4AyRWZc5A7nz/Ej2Z/LUQBtEraF7DMnCpC60D
dYy+QJV3ao6Ru01BbOePy3TRJ655v+4aF2ecaUuveyPDm1C1SBtXq8TRt9qRAxWMZtNMysE1Dosy
15uCx65rhpO6zCUP/GvN/SAjjnkicMtFvU7QqLgplyT2/Ur+XVPvcCy47rGjVXt14MeGORMj0vok
YhFxMSsfLXJ6u8xo8cys3m3PTFy35ualwmrydEewb42oxirc9ELAJq45a7h7KByDbkOOeKjyKciE
acBnF/ATAaK4slmWL1shSJYApuBAxnYUSe4O5uxa2X8RhirKit+39yLuUY01azRKQiw4UibQeDKB
4nNacdITwzTNSw6ndy5nK+qUSmBX24xAv7QDL8ehICMD95z2ovKFNKigUVA4a8Ufg+MHOKiS0L/7
x7TBOlIH5mgx7oCsGtyzD0uVmVO1cAzxRM4Jwjsy/YvdikG2JJ2SRoqA0noRKl1FpyGvAxKZ7gt5
O4ChFxGW41a3f2JZWx278PjkUsM8AkhfEWRaDQ+JaIxQ8ObMHU/WxgxuhdjoSQBTjBLYLXGcOuIk
7yQOS1MiA14zWm/HQtjrVDpkYmz8a0j+OSpwuBtXxNWTuHiq8P0uX0pp3OZCID/imQESKo1ThziF
LETsM0W/EUnqVcbyFR47P0fth08wdnUEwFBE7+Q56SwLaZMqFGWprpRo8F+ZpRcVQ8ycDIYxbpWk
MLMwOrPFiEHQntR0BTIXEjL3d0MRk2N4SIVbESOll38qdZKCXk9ot+V4HVn3QfIKX1Ss0PJ+nEUL
5dgyHY4XF1Jvqz/4anNaTE7d+vHvSo01mYIArr7jsf2KKFqCOcaNdTgciVBKzaPn8F5UbWZGZsLb
sGEd0drcJ262hDUWX0LxoIojhX/2hPr82YfwRJ0WTHdftH7R2tIfSvhJFFFV4QAf9WKTt001goWA
QMQELtMDSM+LSNvHeCg0W2iZwPWe4f/KVnOOPRuu+yD3XcsjL+8fAX06pxS6ov3grFgjZm8tgBD3
q6tp7MAVE/YlHMsNbESlia4AfueoK6FEqLduSrgAY6F/XCAQu5oSKHXGRx1RM+yPFK8r9sUT9AOX
yx7vKL5wgTm7PlyFQxQqDisUH/mH17Ei2a0/WiEQ+rQiYqkBCUsuvnWfEFaXkeyFUZL0/THfoxqg
EVJ03nMMuZ96rp4mTrE+L4Pw4oKef3MqNUYoLdnEC/k2d+hQEzdG4P4XBdTsV6vRxSaQ3/U1vvS6
29LcHJ/ewzb0ksBCBV8l/t6rOvJBVVvPfrG8vAYOjeAQ+nT9XglKKJ3KNJB5nCQR52LPdUSi3YOh
0W6QjwK5sJUBCg8SpvMJdvCDvEs92CvoPrRASZqXRM/BUYF7AtSvtkOOUuE5BiohwF5HXU1c3m5a
t7Bi4F3/yOCIWkMtYkmRxI3uCIbaHxgi6QAGz1OIQjdDCtUCzCNU4eyd5ZzKgs0Sy3EMv9vDT7jg
DFLh0H8d28gv0IZQluYOBf+9DAmksAVWj6Q/njohQyrVD/X7SEPZ1oAPfcV610TrRenvMBZAwL/O
MepqOTC/oORFp8/PQrVvl0ThYNT4qIBZdR8m299N5GLUcELvUfio3wTguWqG1IocLsRfhEeqkmZV
xzr9U8qvVmvDpdP3ex9rcCTddP7mwgYO6baFe1SDe96xj40W2EsTVJ8nj33DKbNCyR90/g+IPevO
1tc2vHUJBdVvbq0yjVc3MT0rk4gPX883LYjSl3i2bxVdBdFkTL6Hw0nJCCfGrqDyMP/MSIoZHPHu
weLeHq515PTluQaSDVEDHHbNqiVvx/9NFZo0S94zdngD6AjmJpTdRJtEJuq95JqLI3mLbjK/FEjO
tWwOOGyvQP+evXDkEvZoEuALC3SkyYQ5Mr6Wv50KJFR1uy9FE/7VubsXTgATRP9gkOtOyrJEtELs
Oh5eWolwvZhHsYYEOAWb8zjLMcCTzB5ojCgOr1A41f8P7m5RWb1IB8CnoOSaY80VS6yfTpL7M59n
QApRgErkld0emr+T58ExGwgcla3ytxLQT0r4fZ4L1piR8UrTUpuURx6etVSseO4wYals76y9A2r0
06FQ37Bac6poXitEx/sE0eeV9+MWzgFX3j7QjXRxv6m8rhI99qMUlvpT05Hnti9KUnnZM/RdyWgz
5ebhxYuU8tIRhroUqXdNhiAZwvl52QF8Cr/K23TooXHyb0EvMSx1CuLv2RedgBmzpICkPkID9Uh1
unyg5/yxyqleeD+RV2Z9fr5tmspXZxuCrNRoAXl3yRqDY7pf5ViE50Vt4eWyefxuba+kokf4zkZG
qU7EPBe+Q3s8VJBwAUbg/Uq3RTfp0IWCeWUArnMX4BT58yyPHCgutaxlAD+7TvwwOkpmoPQhPJuw
Ddkz6lWea8ALObA2JUq89j5rMXoXnumxz42Hzt3YXj7xJWd0N9SyBm4kbyPAq2qOrmc85ta+B71E
RMMFbxGoU+jozQdgJGtZyagKfxDcMpzcvU2e6gWmwC0RQ0d250VC4v5Mxt53iBAgUMhNK1VsyZud
9ACC62kMj2/C+POiUErbAmHxWSjsCraBDtpKInCXHdNfofQ4+CDGVv5BTJ5y0L0s7IwD3aDz9a/A
7j8a4Rx3nbAjelx+6W+l8bFYCpYJxBwxhAhDt/uFcn+bvXLc1Lf8/S3hYvOohPJJtqCLrRaURdko
xFRHo+b8PdXl57Smbx3CvDRcHd3U5r2p8NpoW7v4AzoW6eNb9W3cRebCvjaJscA8J56xw6cG8jq9
+GOIYlQmiFMLOYPfZDlU4nZZYe9SIow2NF+fY6qFDhWDBSq2alCzAweDVF6utpLk5mLozGKR28cU
+pn/GNm+USK7/7LP/QOtz2ezSuHVNMJiUqnQey+HKQe3XiRDnPH7dg6Getlr6Rw6FbqfN9FpxjMV
CH+JDgE+iTuZKP81Q1vz8zddBXV78SvLWAR2JxRFffa/HZh2YOmmuwTUoQkHHwNM7r0uMi8YZmki
pKvX95bu3bG4F7k1gZHbWBxrigQWVXzIQL7S/9jvzARuv17f+Xapnxf/aeowU9jb83d09hEBz5Hv
SZAxu0PQumZllYE1zNwWd6Hz1RGVE1S+C1edI1yzGzv+ESy0ODeCQn1NzNFhjImIPFQgzr/k69IO
R90uZK3gj5gwJt7iqNouL6qbqybMp6CTD8urdT2dBe+/EtmRwuJq9dm1/GUD1J73PANgjIyugPKG
2aDumjZUmUegtY6sW3+11VPjHzsLBVi0r4vyB57gp7OPah33ic1FvjQHlNxAC3DpwHjr4mSpQQmq
XWl5EC8Eb4WuB8HoA9um8ezWCRx4CwlkQF9gZN3GUSCilNyw57AR29IU77Fk/BxhE8IzQxDUmG1f
9QXdbYXFCtum0IAoXz8/Pe/+ysRH7oOlX1b/qBxrlXYgbKZ140qAqDeC1IuAflKT/WbFLKNtW65Z
w+jwxb4wnKQOi7f7wmwxJrEEqHCEEUEIWNZvXmgAPcZ5IqE4A9BAX/XwXSZZxUx42+NBN/tgQrjx
qiWuQ5OS6DdG9wF6jYICJpy4lxziq9FiWCdd99VGOlVqO8Ut+zTYiY568l36eJ7xf01UqHz6tyS4
6KA2jzcb9mgxzsP9yllYE7s34OeJxFB3WAI9wiobWP4G3u1e+CQBq89qU+32/GCxZFNJEnz+/8Px
Ej8LVqwpwpWavEk2ATKNa4ls0hxd5CmzOpN7NMVXSpSwJAYro/ibBUryVNwVOcj4xNNmK6atGhJY
HZS5K3AlOdC8ODM1w052GAVl3GF8CGZje6evEAYCEdJ10DCmWdhTVXirObz8j7iDi8/9d2OvYuir
5sAy1ydbxnth+lh76iMIbVgSjhBfru3JwiYlfyDOE/w6+x7oe1+7maIk5T3ZzaXUpceofPQaj3sv
IlKcedyIdluzNThV2qbf/fx1wbQsG3ZBRxu3hSINGq/kvvY5WsLUtfZ84km7M/vXLYEePmAR0D6V
4fI5nypeW4x0B1IVmTE51N82V/h3Nc80V+h7iA6s/BQt86YS/1AyA4BoevirXxpcGG6JkKJ4/229
bciViqoZ7EmyJWrYbtYuT3gQa31edv1gexqsHdANV0ZyUDbN+rKkgDgzsYpZY/LtlwQrmVWbRMsF
RFjTlx4oX0KOXuigAMqbkY0KV1+7RNudzbJ7GKOJBg7CCu5u9sgmuH0LAoUgS+60N/z83OsPY7Ql
+V3S2YTM6MTTbJUp2qiTohxUKFiy7NZo0EhxotjIhHtxikEpCeT9m55StKITdjXIl13QDRR2wiOs
zQIimCt7+sBhZJiU/1qhIw+78wbRzM5ZMPp/p/YlyN8qO372Ai+SdiaPm5XXLAtQ07KUy/wiR3gz
HOLIuJq6HEAoJoHZNyatHN60R+Giw7CytSHXs6ENvuZi8+WyvqG5EAsN6FcHpyJf+sHzks3hCfEo
UNMcyPNktEWpOWF9qpwS/jB0Q5h0DGnINNMj0XPdQgAugctHE2BQo4eJ3w2BcO/c9RswNybwSfzZ
qWQy+sL2hTuFyqhLuyLafhiDrObY9mdKMWQYI9kuNLLszYBbeasQhmmXsF4EQKMU0r9l5/7hSiAz
YI11/5mvXIT+CPLLXfL1mh3d+VtEiYcmV4cnxNcbkp7Cco7WLhLwMgPmLzZ6fMYHF+NIPCD3rbi9
dN5VySdbuBPwtO0Qc6kmjzVVIY3X4fd+64jQ2P82IHKHsQv+Mjv+ZJ+Ejk7RHpXq+oubTbAY10r1
CqI+43mD9gHmSuwzEj+vAg2VnvT4rk+n91l7/c8rpfm8dLIbfu7q8wCP3PnoEp015pNJaeAgpWtd
TaBQP6szb3XQjiLNt+1jp8nGj7j/74wHrKWc3mXkqNi14rdRuE5NmFTzmcIlfw+qNJkfdNfpqpRW
I6yJtkznzbuyoDsCVwzogiFQARx9Br71mFWjdc6qEOo8F3M97KRn1nX22RSPToOzYUsfXsZp96oO
VIEmYvfcx64QC+nUNsC94iH5k6uhgghdPYC18qzoiaishkLp8eqtoPM2WrE1SOCELGvpBUyD3ENW
Ww+ty7ZDDLAOf+fl0Va1CB206PcrZPgiwOC2GwWNhjk1TIOJOjZ/7mxzjLgxB4C0qImKla3X1W1d
sVW3cLMHPOcVLujx5Pp3p91abaGZ4IHXzcylcuhdAg5nOnHyfLenHsknV82rvUvTfsHFDjPEjige
fFJ3i6te3s0/D4Fh3/TVd0RESbI0ATX+h3pFFJwXYPhgndeQqDa9qR0aUYppQ4GEY+GuX2w4sDTA
i2BWS1jDnf9O8ahWjgqNOZQk/FgnhCE9fRL87m3UNrYK48ND4+NKiAVojEq2Qfj1McgVKYQlEmyH
ZyrOaj6u/nEq9PT5ZgEtOQY+uz3XHLMINCYg8kkoroN1UXb1iWed9dlMby5XSI9Z588/iIX5brIR
FkJlirHffzfNLar3mCRY5hZOuD803JCXxqDUVlMVTZ9FP5OvamaE+29D+SSdGZoFzeP8BZUTzpNw
ZNpXSHY3bwG+hb6DM4Vz2kw8tTl3JLD3oI5rLe6vKJQZnfVoqBf6d+GjKZIs6QyHf1euJfa9Rfk8
FQ2ZuA041lEjI92Xj2mDAvQn8GJAr6N1seDicdJ/keKz4LIgCgltMpgy4rdhwLwan864MNpy+Pp/
ooY212dQhJMrK0wJfeFEPdJXVfbAZacAE9YdiCKjgF7qHfAkC/eDQtU2OcSOgLVJFOFs5BviU+XB
HPBOrPFewWwr2LHqH+a0rAvwG7nP3rNK+ZZckZ5MKBg+VFffut8KXfYowUE3mM5SK0ngS4VG9KSj
iq0VecioiZtaOmAOE3lm5OkWqMtwoCgV/s+4ihAq2riWfrj//V2nUkxA8uuudpWiXZPpa2JnO9Tk
Vizi5tWe6LqMxN2/EcCj6bhDH2Ujok9nDEncVnvsQVe0yVGAIIcwoMPT1rs1RSYYtCh9ZZTljLs+
CInsG6sxJVlcjrpkkhFaWOHeZYcgIzhMLrubJ9D+v+ywKOV8esvzEK4IKFU/lP+Y7rV59lfWRdZl
Rp7gg2G3/RCcLsC8+lxeWHPGgya9qAqk7TVuwiBqqgUhkgV4jI0jPp+/QyzkFGWZfaBNFGFGp2zl
XX2Ey4DDTuLI8w5Cu3OwyL4Oa+Cc7hp89tXbjQE85yKFFOBju3+uwAvRTHA2lhKokGpBd6uFFo+M
yb2y+ssoIJnQRh33VMBD/u036UMJnDuR1bq9QueIVcl/GB1ysOvIXPl7LWJKwHzLjPMH8V2hzk/f
Tl+ar8z52d5dvIO8enarbZXAvA/KgsMSLEmI/7niL8sDsnQeiqpffm34d7BSnqmq9klaKz1SVrMB
ZbRgUDK1eTSvmyWjF9ZDA85xFkMJnk4dWdN1CTb7gmeyf4UN4As/D/SWguw7+DUM5ofWuHl/54K6
OjbXRBxXxISmp8f9oj9Gl1LezRep7XoFNx4vpC/OaqiKu+PawSmA2QxIT470RlZKUYAZ2g1GMEpr
YU3ZuBfEQzZBdTGRFd1Qy7awJ2a6ZnsljOdybkZwUxKmSzHGPr3swfhnTmP704XE+oLfrSIBCwSD
WfIszhuc1qLT8MpEhit1lWQYIk+vLFV1Mv49aZvaAGnm8NOd1Ig4l9iMvJqSQNowYEDhSG/34ZuD
+szniqc8qlavCBZo1Hf9yNf9MpASzoLBbHjXK7qSVCdKy7wftTddFCrMNdAgyAESELzmAwYf/61C
izNsM39CL8Apb6k4nvsu/3U8kdGbY15QGsd6RHcCul3NUVKCAQVTRoK6ghBYr/utn+Fkl9+XAOkP
izM4TIgsc8qHtaUWiluqlFFqsZK6JixGUk4K/sW96Mbbl2gqqx+Wj+hYVJzn4x0SZWhC0Lyq+W4J
2wxbPx3nQJIcZ4eQSJE8LMddDyqb4UTf7PS5DukqIMiAEkj/T5L6oaP3aNGVjU0fNRF+NYmXIHy9
VCSbf/Z9kO8u0rCuBdZ3DC0vNRLt+X51NvDq0vdAQ6ORbyTPHb9o+lloWq6SqKZx7qHakLKOSypF
eU4LLXKGy6DAwJFyK7PpfBsIhN60iWc98tX94gagnDXdeurqyRUraRceHyeWjLsr81q3XFx6fyjA
86HMid56aNt/bpZPSHsK9fhc7FkwtqyICFd2nxTbKfPU8KbWHf9QFsw97KM2RUsU/b0tI03jyGlx
SQKv77+dtPeEF/RlNklu+8kdODFxQBA9ib9oICrDEGgkM43upgLF14EyfJT3q5kboxTrGD8n5ips
Z49pJ8atynJ0sPhbR6nWMxwx05T/ckNlfMzfPpIAeaIjyU87k8leTD2nI6Y9KjY16VUYlUlkLiXE
Jh/O6j1EKh4Owl9VCI2uFUSKvWevftvuCoWaNOjKZ08su0mXniogASmbToUsaRtpL0ClerwJLofH
7WANo+2MFnNZ/5G0wvMzrBVMJZQ2hRT6rR5BW6l5ZT/TG7tYiPa3I+bEjWsIeF2xToBTHKKItUUP
tSok6Vg++qQ8jdtShXbyjUEgdoScgcUlN6JFq7yLZvcwh+rHA21OJ/zgNzyq+KR+OZfowgPKggb1
J1ReK4wc+WEaBbwvTTcC6Qv3wwLYmLAwXu5hkucpZxzmN6nemYpDne/lpr0FIj6A40ibqQAEuFgl
oTWOu8TX0cpbAqKEKT48qqVO1+DM3bJ3m8728QZDafcUSL5OBw2MF5nZgZkwY46/cG/KZ3T4Rhpq
jc7hEtpz1p8rXUDVOOew84zn0+JR8lz8jtMJ4JhahFMjN54WjT35w84UVOesW9Qy0xlccQ3BCJNt
QJH6oDxxyCpwx3R5IDPijsxEbLJk/A3LTiJV+/6WBmaDMLcdf7zEuGoPNr0vQyRt31sr+mD23zB7
SgqZMt/tOc+yLsZzx+2EbHKdrHWb4/zeL3+CaFzssPqTGGbfS8XKZTrQsHNHzNlR6intyu5DmsS9
OvsEjVnqJegyJzHUHxaPeD7i6grXWSFfZwDtIPqsBZp1frZCvR5fdEV52X+HjiyWhXpVZMDxrHWi
x46OfqjtfQ+tAIfpLzasTR2J0c47ViVxk2KCjF2M9HOsFVenJB77Hvl5KsRcBvzA8E1dNZmN8qPp
7wH9djqYDw8PvTuKTrdPxsP4CzSOcc9dYk7+r4fFzXns13Tl0LA1UVS1Hqkm6CGuD/IpZ5KVkAZ9
+SzcMwCNfOvvU38oLhSBdjROWuarAOAvXhIn+Cg/lflUgltRG0rVhqcAI/jtsvq4qNDkC5ykkMbw
VFPxHqgJ78FqnHMzqw7QyGSeVToHcblXwwxnLbSbSfx/xl0IciX+sGDht9BsbmVB/1IiSUrUGsOC
O4TSnWrqickIpj15OFovMe/Yu1bOTikIV63ZvFUWJqSDs+mkmND0Kl+8aos4KuwUyREmAEWfrva4
iLjXIubsYN9s9djjjvIBUMIMGcVD0td7h1IqVxDwYNC4VVLbWHItMPC3BjkJtLxsRqrKkPFhk0BN
iVi9tAHhe8FZVe9dF3N9iGJVKLkfDUxbOU5zb1o5F3S423SuPG57lV/DyF0XcpeG9Hn8MJH4x8cZ
m7YMbR73skcuvczn7G7U5bMccJltqdU7dKUPtY35dqCk2HrzDQJ4W8MDN2k/qlX4MpjGRfn62cUx
LmE15zmSfvTB3AHFJViJUo9SYfGTetCzwGb+NHjaSOofM3eDyRsMsrHOKTXYiJqlFmGA7u/G9pcV
EUiLfBZAUjTOPguj070Hbf0pyOs3lHjD0CqVtGCp5wKodzJ8BmSVgqQXsT3TniHf9WKAVKr5aAan
IBFn7QCW+uLKkhPOClr+XOUuEv7rLVcpuwDNvUtRynypYUIZY16or0DyDGp0tumSOOHN3w0YYl5m
CEP9e5PJVg0pfjVPNgNfTd8Men2KZqFZn1N3TGUcz3010IhK4oRwZSdt9pi7Q/qtIjyg9dxGiXdu
RvauVRb3pxsmTBZZP20PVC001/g1TlcZq6TyZ8kqRjncb2FD7BNiIXkTBmIt5Onu1EeqIlh8zYWX
hfJLAxMOqHOA3Ogsx3HGh1SxBlBlHopx+TFD3h6Mj6jrvamU8BaqJNcv7zaRlm0aEKBfPwmynl+/
VAfSCb0ufAd5dAiCCx/RJaBhfffEOOmukAnh+9io55jBJuuHijUJ98Z2BJqv5YEfhPYAlxL9tc/j
12QZhv8znBijSby/MrepLzQ4tVHzIMptxXRDYfxQ+y4oW0QdywANZg1vWkBXuHuVUZLp7Av1l/JY
Jm6FgNUISIVJkEN5hLVcs87Yf+vmAwbTqEZ1VO909HaNtI+3/rqGxA98G/m/S7odHAOMGd2Ef4du
3ebefQ/yluiSoOlz2efHSo8y61YS1Ps54iA0SARF8zEKUETVLc2v1+g1rlDzdR4mxBtw39ltvtND
tm9G4vRCq214hBcBS4DRzjBNfwxeBRNXq38FPz0Uh5ebRUFYGyE8S5pt/2nI76uQtRAL03I92xdA
0OmNxR9He3o2S4dKwe8nuoR1T5Y/xf7rCmcpQ++obL0tHl6S91d/RD19vkJUmxfi4+f6xUx9bNRs
o4uHriUfgXqYz82YP+LVKcFDdf1x5ePOcQ4fjY3EuK6lNtgnqWIINm8MLokiuycd8AJcq47TbSK2
D6o3iKDOWUTf1zxzQUKP7u2DLrD3BnM4J+y1tx6W+TwANYEWOxwbZSATUcR0MoMK2TD0LDym5HeX
RJJ9WJ5BSF4siZUwVwccGq589tcg7C3qKfUb9FUFV/ei0jiswx7uzmn94vrsBmGMcAms5OMnnlxK
Y4VGViSX01YJ4HNLJAAZ3CfqA5+20G/pW/Z899U7V3Zitin/ccTiDHEUZkd3cbrPPrZdUTBijrv/
Y2tN7ALjU9GZ/FMIXm0ZZejZNRR/f/gi0ijg8Yc+TMvFTw9nBuDSLH2twgv0wwYIQ+/ECWnIG7AG
9UUSQVRw4ITVHiDKIGrN6cGsaMZQQk9hYbTrwfF12exZsPyuSotnMbhFirVyanlsGcP2Q5XIyZQQ
afo4meinG2jRsB53MIV7q6w62HpMtEOjY+3r2BkEv3fYqunlomOaYw3fKUeukKyvFEyYJywXkY4M
RGg+EcdIHwkretB4ABDzMS/+5iPocT21TwgX0obBgqP+cyaeR9Ax5StfOWvnXvPfwMaEglCW8/ep
0YbuuZsqRv9QcDh4pP/JHZp/+iTifnVhSIPNKGmXNpoeA1f3AYtc5JN8lAci00mKngneWJQA/bCN
ODRkvD34B1Kx6axb0lyHTssyOAxN9bqIpFWXPgLsIw5joTKl7M/eWA1IO2B9ECi5q8s9U1kSmyZq
3E/TB6EtkQMl0SOVHTEXPdu1UrYFdZQpQXa0g0VUWYF6oOuoPMr5/m35EPMfVxfrT0HsNj9DnsRH
pIvN0H9rRs4pMM2adMqblv6H5Rt9glVQMbPhwJIGwPadOPTFKK9gVh34g/0IGqNPBhiUms9YIgZI
Ht1fbZpg8mdduhFwwD742PMpeIflI3bWBIkmdVobKwL4DUqIBBVklMEyDEXgkFXR0H6qok7WTVrL
FYcwWxpN9aV9v7BIX5JbpsZG6uAsfVMrtuF5fMuK179mE8QuKjYwp7BryrrDiJVEvijkXqShFG47
fOpiz3MbUgvPkBiNQ5M5+6vSnBNbMHQDcfjc0AuhXFyYk/qcAWBPrDw2GcJXdjCT1mxbL8Qu28UT
Kx8AM6m9MxDY/zfurNXK2Ss+OgV9gHa42WpLLT/D7fKqjHbVSO8sDfyDUCC2m/T6A31V3KlOxaRh
yb98Mn35K7dpnYFfCPdZ8iKfsqmlmNISao8A5rFS+0a6kvqp4yXUoS6j0qKcUR0KbKbifgdjul/l
EfqPyXJGg/6GljKK6PSuRhbpZ9RmYE2i8uc19K6ShgI9kqAaJ5Pe16jb6w8wRKvZVPnGpHFVFTMl
VB4tqoSZAlj+DRNPJBoNsg8s5rh2fbGbUPjmu6n9tnXDcEFqPv6HbP2tx0wzzQ99ng1S6MINMWbF
oQkX35/xwNOFuadsj+/+xK/4XWF+0S6QvqRO6nFIWzcDcn8Mmd7WVL5opnMxW+kU038EVwIlQwEJ
eOjHD2XBVLNqimIGLdZSBMBgx9EbO7067ye/nWiZ/sLed2n5YCjB/hvQrdfoACNQOF0+4tZSKsuv
9PMSFboGfTXPRREABQL9iz4lHFj1hCMK/dkHNxryJqCeXCtYAP0k1gVcmmxnsnfo8Bp0dmDRrdSH
Ar/gHnBSgCm8N74jndT+jHnwU2YQ5f+P/2ulFRHVZwAY73boyEUzbqOeSV0ZgiNSurLj2qi3KGCL
qqyDbqXfImrZupSbVkjnlMgGJAp01nX2phSlBrEF1RD56uzV+/BLejOiIQRWc+BYFK9bvwgQ983R
AFxLqxiCeRkDRQU3d391o/4dxgigFA4tNhf+DZ4bnxZeARz4qAuE+ggnwU51Y7os+BtJfgWp9CKR
TZXlcbiMOoSXEKNaIXGtpl53ISr+GhzInbe7f5wM5VxeEOsG6tpe0s+RJzMq2MIBUONP7HvF9p6A
XY2EdenbW6vhPNIH78EEN+YewBKLte048fGucsfa/waVZix9f4nZ2BILrFhF9CdpMTrjkxcJU2SH
dvFC+5y7VIBPrXhUftRsJ0wuRPGzWl2pYhMAn3OMS8NRVGPD/5Ck6sUChwmPH2bSn1bmmGvZ1V2j
8aayK0AGktDR/BdvWgwUk1M70PqJvEsSUs6Dd/jvzt5z02qMN43mX+IBG+QSWYHRguSW29bSvLdf
XS/dhy26SaiehRGTTxoE027RarINfg6KB83imyKL9BottRs1YcSoSwNyseeIRSoang4q3lw1U0+X
q8YKscgwdSmFSweTc5B4qUTP0lvUGtYU4cX6cj0+jz6aUv8ODPGxwn2G2FzLacLUVwKjxGr/+W8O
sfbnUDkm5jop1GWTYpviAaWhdN7Buq1y/xV57CWTOrGX7/YXqbjFiuw7gOkXjaCwdaqJuja8Vh+i
fvY25miByg0TZbEMoZOy3HCsnaJj7FXuLEgdYZm6S+5H2uNzFpsHI7GgS0uZLf91X3B3EaceiN6J
pv5GEb6cDMwK+Yxpt9UDOJd3SXfrRJB3dh0/jDF5AU1Q9hD2iljGwM3DMoQwS+rE3UO8kcX/It6q
8/0RVx9/1idCgTHMkWXDb3ffgcDFOELbREm1c+4s8aXt3NVTQxmUuSUe5V7Fho9upzG09s/enMUv
HHQ1YJxyvKq2HmLWBEDhZQaEpSLUhgaPWg2ivXqyEGQfymfNT09EcaEcPGR3btecHoetCkuxAZnX
1hr5VAHuQqqcC6YduksdGGAZyFY/H86pPq+rFdDMat4mJ+4MXjGaLAhlKFsg18m5J2JO/vKgLxxj
OyhOokLthcjdB1iCWG2qpazEC5aB4ZD+zBFKjlwwWgSJDDdy4uy5p7F/Y5OHWSdqm9RCb58roIe+
lfKvoWP8NLVkJ/7tLs7HY7gfTQfW5z28iwbUQNkrTgXnZ3Te+2QlDGbGDousud3y6P36Kbg/fxbw
wvI6bOdecnRpbeod6JihqnD6oZ0cWGXCtRGboKT3G8PlJytGJrne2wJ2uukgQK3dWiNN/Jb/4xnk
sczUsdnY+kKI2Wvd95C7SE4NrwOGK3dx5G4kclIhvfFUO8nYpYSPEa5NRDWKUgbE3dUCeIbuPDph
kGHbO0n2Nv2NFcaYUMwXJkwjcVIkun/lH1BAIDEs1X5uJIxIvhJgUlVvKPitJDXxQ4V+/Zy9zhGd
EEbid3cThuUIgM5kbxEOI7DVj1M70nLHnMA1rOPs/6r0Yn0dT4EHwuaNZK1vaHH2z/5XhJ0TPK0k
n5iA7ZTNOR9Mkydj+SB65HImaus//FgZ6X5F8HVoG/syK6ZsRoqI4CNqVCLWcsbZAitsVq7qpQ3B
xlg76nGUt4AX5QtXgex5UZtRO3L42lfJ79DJ3Myv/opbKctuwtoM9dDMtS+wB3aJot9E/q+E246w
aABFFw/GuYkNY3qwA8hMlk/6wnnRzbWd1fjNoMYWcb+z4ezL+rZZ4SMlsdE5z7IZKrk1tuSu1qQs
SLk+aZFWFXR/ahGr5VBYnf0CirJHmcendWZV38PmcLAlNdA1yM5nqmLXSy32tw2dTkZ3Hro7vEHf
ExtJX16jeOb9Zip2B5kh6+RqHYzy540J3JlvguIhF39KgJ3zMAf/QCcPj7j4d8fK4CEd8k7e6E9H
7Uyi5n1FNU/7HvkGjB7pOT/O8QgSNDWtFRiwSxJXsUMPCnmlzgDkmx/BPwkPYE5DfJL1rRtZI52O
XJ7poGiMEq/iih3e58az2uhLtyw4hcYv0k/zRGlwbueOp8/nSBbvRhhQa2mP1eVuF64Ey6rtH2St
EPT1x4DsffFGR44o5PhMQ9CeYoxo3GKj8GDbaqHDQNckGAMccayB43XxCdq+q/x7ep4sQ1WJ/SlY
Y15A6by8N3DQ145WN4NB1CnMscE1Jnb63AFrZUzH33vPfJmbXvAKqDT6Oo4kERzAuQAzXNVjxEuH
4si5UOWKq7xGs2muQhSmFl5WuIbcpTOm1EHnL0otFePZPwr2HaLGdcFMIx3t6mpkFG009ant3vis
OCmHpG+DS4d2W5K62g2hTPBttbmLNkTprhL8KZlwz19hxZLcYoFjOgoTGO9u/7Xp7up/3vccS1le
1azEKcWyyt8cW8/lr+NncB0o/NT5cluPlxHRtmeEeQQ00pE512o1SncsTFmuxZyktJ+d4+vmPH1M
PrNs8CJyuwSs+KdB3X2XwN5bj19nJuW5G1T8UieLyDibgzpAaM9+RmGBf+X3JR+zGJA5X5awPHcY
ymXYE19OI5KVLL8BVuEoqzsp9xBGL9D6eEPcxHpXaCzQq/jGN2k5w73WF2+0Ck3Yd+EBrkyqryhg
drm5eV2HtYdKksaEicF4Rl1DoMwh74oek7tINi0wrEGjhnB7OjtSpi/KRfsvqpVvXwP5r2MWL4Ms
ICLEMPvpI3LUDTDpIec3k6ZMHp1sfXs6YckyTydpxCqdSUBZhrM3zAZFVEP4dzdLjwvZ3Ljv4pLl
Sb5Q08GmJ/Uo0/7rYH/D/STTU2f2xSx29fsn/verwfAQcZiyfBhgUfhtAIHBsRuquda9tO2iVMbx
r30d2DkAw5NDsW9PIgnp+0gNx1Bz/oa4v2b6KIwK5vinjwLjJENsD6HG4yDPeV61VbCyUcvwG8/m
/8TsXp9PmCxuCxCpfNpIlPMmmYDRmoG8WVtRizFRomyGuWrRxIpyNoLLYWTcNKRvRpLgzTumrUIz
3k6vW0nuXcdgYcfgoXkozWPPgzqbMRc9B4Sjya3UGkBnOwSCw0S9Ja1IRPmlUD9pH7EG6ZXUQupy
zEYpGwwI0KR6ipsm54bEX59vrgi7asZ+5mWZDjogMcWGU27vk58Nqm7TPg9ZVZ/Al4oDjjtkmQiJ
STT8NPISWTV2T4/PLbhcR7Z9rRnV5VNGXDFL1oFi4LNkRhITaxdbQQuuYp0Zdy+Yj9rc3CAsZNi7
NfzOxUPZ++BYGxyK3Qk02P33Kob3UUtZpUkbSaIIgutJ8UKxicApwdzUOJz/L3XpHX2Yi0uNiZIU
xijcQK5TBVo6wm00XIepq7MwHl7qOtgB4MtcUliUqcdVxHZOhPyuA/SGalwlT/wtd43rX1GRPxIp
lxFhzZ+hUupyVLLIDT+pDr3yLFbXhWBg21k86JPs/9rPkOblqRFO4T8AgAnt2VilwaEa3EXLHFcP
5YXfdao7cJG9jFNR5M4rUajoLH3QzPxQ715hJsZKSV7WpFdhe0YnP6i7TnNQBSc4TgM0KC5rXmKS
zPW/IkYguMrjngquQfog2NgLo+nV1wxAUy9azaZ3oWGmdTgotdZItiMRPSFaBCpBJkJtjuST08bv
ETwkw3WeHABQXvy+2qegnZpsD5TXV6/j2I22GghbjcR5/9bEgMVDjYNo4XpM1HqvzFJpJHZj+D1b
dc/h9EvJa4exNvQq9W9Jip5WxS2Sb/75etRRVmEVgAJNWy5d4woh9WXuyRdoFX9r2t6YLh9RJ+yD
K4SEH2iWYuvv7sBMnQ7ruepaZaQFnBF+qUIvhYg2mEpsJ4llyVBNblHx7WFO/JwXaHJ49jXUXAe/
cQUTLt7vRJ5lsTrqAugseqFd5Gl/zXLMUdoOPDdbzGSsc7m/w3fDN9fYIEYoaDeAWwQqAwb7V5Bv
vj7l8ydDkFqznXqVFQ2nH6coQT4P6fBX6WcG4WJwlgtFS/O2AgMV+0lovDZTAOw19Nr9krjz79vN
yrQHrJpiBI5abFilhalUiZBv58QIBdhE3DramU9sKju4LP+H1+jwGaJqT9AsJ9dtWSzq5ssYIJLi
SBMKbyoyz0Em/lkAMy1DeG5qGGhUrawP+UsqTNI4fXGTfVy1ntGTX3L0SwKLOKBVwCW4xOb0cbOi
jOXVhihJa9EzEmcvwJagpzysDpsk0Efl9wFl7dUcKzb3Vlt6mJhKlfycEFp0yPCUfMkjaQRQy55u
xaW/fkwwNbpauG4S7nfgh0qEqeJh/JxoRLBVlqh4c0Rbx7reFP1Be7Gb6eQLlvQfIb735MEyycmu
tqfprzbGVNzo8bJYG9ZiH+j3OK0Vf6f23K/XVRm4biK/D9pH/k03hd5cEzw/0OVXkKnuHjmEgHrD
fC+FqUW2ZHxSY+irC/OLKgiOYlEx+gIWoSSbmiFkZn04EI0ywY5+xoq2lQoB5LPqZT8AQHDeufSN
y5t3a3Qv75ws4wh1sAEInC1vDL9QjT/GM3v7k7r0SVbGRcRj3pTxKuUe+diaevXMdL7P4ScY3fHU
2UN3ef5qlrq459o7Te2au0pn5iFt/3R07BhPa54qYHtk6TJTWHMHRQnEyYwYfQaxUvcrNzZo/qul
OfGd9KGi8I0gMsXnHA1uPgWdiTbIjt0gsKfX7hycMj/0Qa6RAshAFQC76gs2k2kTZ5+QMJ2duhaA
VyO9OTJj8oUAZQo8RHR28bcujIbM9ZvnMK/Uq9yYfVqaEd1hS3SL8bUUUjLV8C2UyP8OQ6/LE+xk
C5kaWAT63mYZrDSjCbEVAB690FzBfAkPt6D2kOS5/KyownwJ9Hj2XCIWJ8WVtWnl5Z+vnoASLv2v
vD5oLSUYKqcCL6rOya65LMnsI8DewdBfKqVsVxyn2Yige4Y1lXrAThFvGOMrT6WhTBt6MhXF4ZkJ
ALi0thqsP1d/7GCeKfVMzsqtuZPaHmRKmCryjLduzRPvAp0CvZEe1U2L/pYoLFTT2YcNGuZ4YEeQ
DmRIq5OxiqgGZ4LHaLLxdGugVPK9JkHIGuQoC0TlA+AMUgv3NYNEVicyLQTBYy4o7pq3mN6eEclo
paIkFaLukmRfImbR2fSk4yZMThDdpVFi43k6zs46HNf3MNwaDfakEhOyvSn1kJ2scrOZKXwI2h4R
cGZuASqKEs+5DE/xumZEVv0et4Q4hnN+fg2t/Z9ebB+B0HMim+q1LMGJwr30Z8IdSNGQaCArQHSo
1+Tg2LX/5MHIAHMGfiAgKJa2CDIwCYx5mVFtWPDjAUONa4wGPJ0hO6e8woRi5LAzIDVJ1CseBs9Z
6UkElNcvs27X0q4LiEeVJK6A7dafYsDRFL6rFqOXzhbn3bVkVj21zk4cuDMBNE9zUTzvRytuKP4B
NLLMdEZqgCb0OZxNAtGGW6iM/M36SqdR19p1pJ7WhxiE7mS+jGEmRErTwpiLUCt+Fw3wsUzkJ3fW
34PL5px2l1SiJSqhAjFT+p/xax/bg6dWPDwyMJlgCDUdpyb+xo27f8m6KCSOGMAxf9zEMGF9Uw1O
Q9qxfaI+Puz5UXL+e1f9jEU3Yp+bJ/eNSEG/2diJwYgyDA+TfRQiUkSYMZKolt9ogyPQnNf8MzMC
sNeajKwYMLYK8shZAKvLHbTiS8PSxyb3102li+aHzfy4YABTQtokWAEtjgYiqmSqUfKq7+LvsWKL
gr2Cl7f2fsBNWcteEB4JhbSV/Wc+KB7qbn6wMu1Vn9cLvJbSgYvDl9hJDprZVYnDwVgD0BYOasLP
qQhI+YjM0rAhqqb/EQvkxXyyVVc5GsyxfSMj5Zpae6SMj2hsp2Ckt9Nuyyydx5K7dGPEhtl2NL9X
YM29tgxnvFe93SAQ+k2D+TTVcejTTZtEwfnTaFCY18n6J69oKh/Z/tdUInFULCMgWyzTeIncbXku
gwgExagO71J31kPpjNdc/bYNaF0jMUyhBvZQlF+y3BXHiVnUUzjBlktJzot3pPgYJbmqO/DfW3RP
yCiLhDZZq4rOPSejGsYLhAvwtfL2qw33+A5mkdKyI/GOhyYjfRKpPfmfIEC3Po6DJdEATcq1vzw8
u1YpOaSMqK/eSx7VY2+n4uKX5yoI1zFQQB6ktIrvqeOW37OHd/2hFHbt6VKEBiL3vOV6V8LxyynS
4Eeyisy2PXh8npEUqg4DipFo9IPTXVwZq+F4MvhS62q1rtQDAcSemdKqwFfpGtKzRSu7/dr/1q12
X4x8Jii4859qN3CPlxaal9YOsjG/8OiO6XVKhgX0EdQdKo/vju1BlqTShRlDpB23EDZAjTUDohKR
/+buRZkFdc00G/CLLugEqvwaTCebBARvNhzxn4J/RJKVJXuI/IDE74cAFUuI48qlbKT8I2iR9GUN
+DVrpHzeIiFYpnAOsMbJTwZfgQl1M8Ev30bi/eGPwJ3pGVgwOTb38+eFm+hmx/VThNvRyB7Q6Gxj
lLba9Dwpz1JO4tlftEYH1BrljjGOuZXvnVJSr+YVPEfrlgXWsGzB3xBvICevAgsWobsyl7AP8G2g
VrpP3CIWZgQarHPNZn88j92MNcY97agV3vXpE1j0Aw7x+OOLmpirdlrBIkWN1+vbGsIJFL8Gz1Aw
okTvwmdrFNBQG8SSrIhaNdF5E27q4QEzdOAcqQmgLlYd5pvAdfexewNoXhAmZ3RyNwkFvBUCIft8
Zv4sffQCwGg54XLBOTsR8CkFQJf2CPS2fIPkTb0JMRPiGFD1fduuSX0JLt3nANfJbwW6wq774hYJ
YaeG1pdzY+VvF3cmsXkkGuEpqk2RxcmjmoSWUp9Z8B9SYUfyolT1fjc25din48v2EdtTeH8WJrPB
k/hY2O9qAWPLpeUG4jF6eV98chzxROUjcIuqOH0Mudn5woe/ToVM/OLl26BFMj6DhWReGjDKX/Qq
2JXrzmwQLTQ5m9k+sfc4nRYrowkCFAgf9y6fu1JATMjm6yBOEKin+gAIlKwPq1gojbm5NnrXTVuJ
CzgcUo0XDna4hzLxg5V3oC7+HXp5Wq1wqsgEV0axL+k8rh2uFJ0zyZrzPFtpR6y7DQX0Yh0UdO5+
YoyBKhC+0DbZdjaQuDky0fUjDaU3ldxCOnCkz+f5Yiyn+z9i/KR0rI1TcD/YZ68HZPMFSUOVhEPk
vXdwu4n7nB/9rinbhx9C4tJ8Ax8lENtVhku4s8eoqx+02gj6UNFqytoBt8p8YSaS2lGg0xRD1ub6
6xLqzTWhL+pWzrg/D3f8wbX9Wj+PTMXBknNTXpwxG9N0fxu6x1LCJy+NnNLZXn6PoctpYbl+GHDM
NC4mW027dE/JcRNWDY+fDN+buD0WiALvwzkos7kkukXs7eR7naQHvFpjxYbabsIikz9gLmHEeldc
6GHI49VF6IyLnEEIClV+rpMWhDYdsYfMGYVd/MRrmN5hAr6hojWd0sw+/RNkMQ+scnYobfnOTCTH
IawCWe9zGdUgv4CUG7X3Z60PntJblMqoh35su4GYlC6OJewCUkoUlduiCHFvLippc/HTi0LUA+b4
jzQ01eqI21ZFax/W8ICW15cxF3+9hPDc2imS9r3ejr69A3hjgBVLdO3xYI90NOReucWV3p6t7NlS
952aPFf6l9OvRhoGnzkcnpOcfFQBrx5IlfXqJm0CYhAV69R2pDmle+BBREKCdMezUnWqeMxLU1Ay
+U3yr+eYHdIg88NN1Y+ejOblE311laHUteHh/XTJJM1RWyAGoHqNb+IJAa9oG1E29Y/sjAoVgacg
pFSsJW5PMn6y5AvbNQtctAAyhMq8GQe1wOwMKOlQ6kLjpjeJvP6CiqHtWx8UibLPRyu63uk60sYS
cNJCW7aMJG7tkK8ezLhIHuSOgGNqn/jJ9AswGtOuN9gUZnDGasHtMqSB8wG9wi5h4WwjYXd8xmCd
BudAG6DrSfSPn56QGeEYnjHdZfbIT+0uj+Fi7TWyjQXR0E7pbNuek+M4WpVpwzArb+vNIVkmUTXU
ddHwWe1dSStrapvCUhbDhEeQ19IUqeJ0HFfKg3a/reTdF3RLMfBtCPBKmjTXMsCmYORSiwIufQaR
auMYdkdZvHQSjqNg59tVkjpIfBc0jQErLOqo9XJ38o+EevW9CyHrvV4bg8k0+d2p/Umu0teWzZAf
BI5O8ukOhBSy9RI+UHEbGlUOXXeyfG9FIFw/HqsUsyBowDLQDilcNlKxDYIsB4iLe4cYSJGqFG1c
DJrJXmh/mMJs/pu0S2DQv9kOVSVKl0CNzLsPm24dq9elJ6LNqFvyTg1Sb2Oaa+ZiLPsPzsWmDyfl
fWt8kXFhiKc+DDCe73lCFeiY0KgEr2ZmxV54PAUnexVra6a89Z734zal1wddJkgMHWbqJSSv4Te7
3BQ0GZOZHAgcwogL4pWD/qutNDg5k1r9/ovAIK1WDbpYa3mj1vDE80gXfOnurtLpUjp00K1Ssuf4
e5MT6mh77rBA7gVvqfJysB0nFyg47k2BoIIhBValuukHYix21s+hqUzGzoP/PrY9mLiGDcczM7h6
zxRGvesy87ADPOSfdVLWsqBIL8BZmPqKFtKUYxccZpJ1gP+oj2IUYxM9XRh7cbSf9WUlJ4lG7Bsi
ZZJHQ5Y+KWRPSRSboVjBd8EeLBZGIKJ2MylS2b16LdqmesFOvCnUzfEdbS9TGXO/KdicVHUzlx3z
CzatlxecSogt0GwUuT/EgxKT3bvfDUpy56PB5vK0/mmJnlKD7aTsIvSYOTNoTm5l7/VLi+wtxATQ
OY9XNBHCDOxcl9auB52XDr5/ZZYQT9SdpEgrMIF07KRlWMRx/9wq7/60nopxsAufoXIYEV1AJptv
RPsCDJLgnBd5sR2dTJGZXRlkDcXUF/O5/oL5MspqDNdppHbICWfCF8l/juJk7xvvzRGdRVybqhOp
87HhSX5nvzxb9Kwjig4elDXLwxDfouIdp/ohJoOaWzFrWbyNeOw2s3lJNM6v5Vowtj2WNFid9IyQ
bG82qTFgesyAlX6VeZYLxT5GriYpzi6kndSWn9yd2jx68FtxZOV1CkPK/Y9j2nvGQEUf2SY0GNDy
GP6Ve68PA3B/2nOjnbfhO7XcAStUrx2Q7dFnriiUD1fVZ2Ijohw/TK0y/vj1nHWPq+DpjTEFwliq
qJgDRHWn/EWV0GuuKKfTrPawr06KsoNa3PbsnbAT5dISQaZ2wCjlMmTxzaS8OrbkH0tCL/QSp8tB
/rdcaPz1+8bwObcGAszIKBJ82T7J3+DqvmrucDUDE6YzT3/12cDetpMy/uzsKJpJiun5oeYLR/Hc
qfc5w2U45Gz8zW+leINPZNS2HXmtuiiLfoZAwJJbBOLjcKdMsxK+6QT77TEU1VuU/t+xOTqu/JM4
GY/mjnhabI5YxQZJnynSLgl76iNIY4/R4siMF4SrMT5nSwAcbTSsp0y25b3pKS6GdhUharAoiMZn
i8vsu/j1wKXLXPu6GVEZR8GF80S4st3CGiLDRngiGpV2PWuwCws9NQaA8DBiNk7w6q2PBDcBTOgz
qM8bSS57y8UVVqNVRKRY7COm930WGySEFYoZWXg4ms/7sszoRZQyBUu7XdA/XesrUhkgSZhj0ko+
k/+otGIYC6mOW16J9NriW2KivrttH0j0Fu4xBkxuV5taSAzFizDZ9vmSoWPWd/qSfKzfhFiFnrvH
cdrFrAvQ9RkfxTlh6zRlJmxfYkp+g71tollL+ZtgoDPempe6jqnxtb7ZG2qunoat+zIaXFgM+4j8
ycs36AfharPT260wu8pO17Otg8BP1CkF7IaradgjCpf38kUZJm9P4+nu7vub4BHI7wLdW5PyY/FU
nFiz+Wjg5Jrr/VKPhsR+ZWVIhTXM6YDur8KX3SxARnU13Ut9BniVZaHyB9YI8z3jGEAtGkS22FUe
Jp5KTXLBOtQxnw+yX3MeQLboUcruyctdDCkuzc3Foofh3XgriTXqX0uVyX3OAgbRkD03bHwwBjwM
yu+d1HPREvTLuz+2qSlQzbSEoiIGLfX7/bh1Ev9S6A0SoCIpOY2GXRXGRdsFUhyRjPoWfPfg4r6E
KRgrdFktUPvFxpuxodj3833NPMEqbTl/sMR0BI6KWnzu9rqxYR6f2WyuZhz51DstrIt5h0eJsYG7
6BSRUOCI+FZZVw5ZusmJRFdU9WgaQFpIdN4aX+WSG500pkVaKj0CQLedGVFqm8akpIoA7GflthIG
e8LIEwqpUSOySiQcFy8RZp7LRIOC8qudXtu6PErhgDTA0p+SZDvQTEBkHbLCiFlZoMjxM+b8jEqy
dXHR9z0FNQC8m9fgPZiqXC3NgGUYGlk2DuANsmpVW/rYwdJadoDbv8kWEIQnD1impB8KpieQ09z1
dFAO5QFX6GIYN7CiivHF882iy2vLBpnaFWx3jDp97Z4+ERQMJxV+qorztJzitTKvymhnAo8+Ej77
GEBIre5p62mYzuvjkG3zkqxjiGhnvrJuoW9KawaLsepBl945H39agBZ3OnzZWQ6Pf/mXQoONx+rj
j17c6pL5Ds1H8tTMbck3cWsEdpVaFR15Pl/+rpM4WBa4vTioG2iJQD0rIhsv9FdvvJcHABHr1GWc
65lzUdNxkI+Qj00Wjoaf1jE1JFsWEmGz9SkxERvje1otbiBFcBpK+NoGRPDZmkn74dG9X++8Pl6e
CPIO6FcHQ/kDIYfGxHBsef6LWgMk24EhJePxoZLicLACPf4jcKjQH1ycUIFz6AZ8sgEuWW0i52Ui
f7eftOXxb0Xc/ko3SaMjHyTNMyWhfPsAK2+XyoLKjHsNzP5TrXqx9iCRF0xPq1gblA+fePXvRfG5
DIBlDRRgwaoj1TGM2UjtVG149g6oukaOl0MA7x4Wp4rCc1RsfNlTJM0oZxAy94+lPqeiyfylgkj4
AV/i9s05FeWLkZX3yNJ34+651sV6/cBShDjKZdZVzoev1m6bxa0wpXxIDRhTQYt09AXWrfv07icl
iWWIkv8SzL07dVJmmzuqdyAh4MqawauqJVe5pro42glPZK/2PVXa/tipLGE6GbeEDmUGejjBPjYs
2BgPyZSijWnPueGuTPb8DuDTpWpbXF2eLOJdkoeAtKeMbhWGxNW+ORmN9WTlsBZbYfh6+FUSJYFp
mkEWh1nNcKcGyFdJD2IwyfPq3EhQfnKzv9vxKbDAzVsyqi5RPEiM3EWWOORsS2pXFBvMX61FCXeI
8YNbbRgkhfvQ4fFGJIqvh+2Ylx4ybldZxJx6ZuIQRTmnQtcBfUYp/RDqFf10ZdhXxdVG7BTLTqfz
WLk+drt38RgJ+9h05ZYiH8VbRaC0MZXOQk4VV4otbD3zgQ/Tkx+V9xykkTUBBylvBXBba2Yj+1Mq
OTzKG62/BOlsr1f2onh+YICgR0RCBWbLWVkoP2kyz4Xoy2MaRO9L+CKjcCR7+azlqM6abP/kVBnm
7G/A36G7yKjM+eOvZ0Rnr3nZaZaMQQnNjW2PQrKpFCea3YGv6TKdM9VxmvHu7EZlPINuUyU3m0oN
SfjrJCc5EdrZVWjqcYs8Jj0H44uLhwNFNpf2KSCiXAr4kwcFsrYQaLnkQnnMBNDPAxJHDuwBXMuG
TwtyIwxQqFDf7hSnlySOnMycaVUo8qORLTgcmgog8g1LGv/dOpO8MKPXMTJU8T7WNeimwyB+1bzG
LI1rGXebPcE3XkjdIrrV8D08Uv3gc+xGNPHzttQSN4hmOKFf/lzrIu29uMbg3PRmrOIRoe2xg8Rz
tsRyUrIDW+c+0zzOaNebk+YBz68JN9A7oOYonbedB8rG4LdHB3W2zYinXiMpvAcYyvm0sOfPHPv7
mxFjVqns2auislsRW8hjQTz/EvcqpeMS4cAyOpXMsNJlyADuegHbCZJMrkDjMTlRgoXOr3I2vwsY
LeWJphds2ATTrRbKTwRwuxhiuWhReL6OXW2vu5IWEqfHQVJtbGYyNuvoKOr5w/LwgeOXcfyoDADf
CNVKE4gIOdRaqyI9HS14hBzPgUnCYe4KGcrk6pH/sX4Sng1yh5tGOp4RFxLPszM3ZKssm81pWiOh
5Kl5fk3hs1dghyV/4IdQEQkxmDcvMCpK0i+U0IpVkZhGScEa6ZsrUTxkyTBVT0c4akfgDnjnSsEZ
r2N+L21vyEiR5ZNH98BxpQrtt4QaWCMBhZkfbrSMkX4SZFW9DgIc4yPlmZfAu1XbkJ1JRYnFLKk4
kneMVxRYZjbhUFwWk+1Ws2zTXcPDECzeFLfohW7rxJNM3mUC6zGQMsfX0GYCaCYG16b6JaGAjvCH
fHIYYfRIEm3+ffFA5LlqO/AE/37fuZ+j5BNTnOEtz7nvFos/ucQuJ5QSgKWSF6wVmjXCFlvV/+9C
JkxCQdou2eEBwCgO/5ccIwfb1+JC6O1XPxpYz2zE+eNsIcG9qOQh+FZwzuhTNkcXFzoD+BCF2WRd
XPM/FHpHgU3FUaZgEKIJwcp3uycTrCnhGb3lCvZ0tZvOZA4/TCaG4K/2i/8wSA2sPv4+eKUfB+5w
/+CxucH8YZZ9G/kHsr/yglRJgsUgbV5eeZ0InQkw4rZ8pd91rml8bpcsj70TmHfPYYXLU4hJfYSk
z8HOEx3acweQL7eV6QvpbgYGrcnGpXJgOn19vniQFocKx3gv6ZvZXEh9AVC2KSj4K1ZPz0nG6dIs
esae8LypfASr2wPu7GpykFss/esTyCe5hgHvQyUypAX5+MRtfNCyEvxGVfWOE2kCneghPz6GQZDd
uTL85fHJSyIUMc6ds53uq72WAeOQ5Gwlvik1zdmLsfzNe/prYOHwVTL5paBMpxUBmdMu//rageRS
nBQuEZ1vTRmmyPXWxE1OLiD7OYTHkGvDONKQ/ZYSFgJHkhWNWoMf0eG0hz+GDNTmJj2N64bTe3yy
Y1xwKM/geo1XGbuXJyiXMvmL5+YQOaFfLJSYVN3AXBgcDwwhAJPAWSIjljaW8QiYdmZycNico4ll
Y1CwJPjNPzpiOh7J1agB2keOqD/dPweoYecEIwCQjQ7IjxZm6nuQES1PBr//5pP9mX80axDFzSRi
yRBXUwSxdYmHkYqKzKjxMgkzQsr9Mb6H6BYKUPWhlH+iJU8AUL2CkE8o9gqFbiH8o7Y4h1QJWEw1
H/WwDMvX3oEoQBULdG24DXdC3bhejbf0vWhLQxPD9E21oAhXCnze7YuRUZQUZTZNu4sYkcxsiSdS
VT/hEc00CLS0kO3AOlWdCekRDv0URH9lGMossBhIN3I0PdnyR8bfLKEcKgW9ZRT2pOFuHNe0oxYZ
Fti1y2mAXbC1PAecs419+2auAzfAfoUM/DQe3CHb1m62G1xnMfo0wiZS+oTzerkBIcz2oMYgH7fQ
lbcNosyKzD/rxJqcuMCX/ICSl5XNhNadSjgEzSHlR0f30Jsq6qwB1t8XRzYIaFLWGXiWeDsUvcfH
FVRJiWE95cFWQBggpeLxFPE22qr3a2JCtClnT2YSbyCUd5MxffSKBpEyH8RpL8NED+lVwGzhI6Ck
lT9wY6rZhnvJVIFI8G/XnteRy6dj16HzB4mC1t8BrBqwrQOQXvN6+MzjJOmfIILzy/ywNdf52ZQ8
eyS3YWOijNQXhpwWrTdO+w1p01bvaD+PAHqeBtN/RO6qBTrVXaEJJPwP9XwQW8hma9EkcazSYFdr
87ltI+K+5SN9meYHfGE/fxMeaywf0xw6gIVz8DeVl4wojE7QG4AydgAdlmfp1km4hgouJeI+E3lt
L0FvPApzJqqdr9SwncNoI74JfnvEm0tVIIGOWTCLxFh5Z20fg3dhcL9G/qqdViai1SSl5S8hGkVU
Ma75mq8BBFPy/Vstzh8wncOiWBqnFciotRM3Q7SmL/DNT2/kjqAmpkafn/Pu1ExDo66o9KthsDai
8KU3QdGIbnSsfZ0RY8EclFtGJdQrAurlx6Bmt58A07hq+kIqeg3fDr0bEc0SRjdZUT3EQStZDAUW
jFpNTRQ8wg1PdMCWPWfpSek66v28WSMTVW7HuXyujJyUKp7vZ+47/KDQ26wMZVgBmJMTwEayYgoT
zud1Rscv9id8a18u0A2v0acMXZcqlx6V1wODjpEw4Mowh4gc8xOZxwUC0j8438dbqr0hyUySiS7E
+YSd9hpFj5sT1KVcv7bH1kq8CHgcLSv2AFjK4ARgTwxMiqp2fwJhp3ir3a1fnjH31q146xROSwVF
GkyzoSeduOQUfevie3t7JSJFcxDzPveBZni1F4UqxNcBUXT+ducLNoLQ+/aOntgvDWum+/B1+uEX
Xo58gFiPNLU8SfEz93aInVDOxfhHmXfVqVXeZScI1X6F74NOSTI9RcvE6pEapevF6pm0DCV9hyc/
vD9keTcbCDfDFh6di8lg3Rue1K/eUAHm19Vlh95L272F/TBxAtz9DMhOrqJZJvpCpWZLMvrWNjtU
QpghvwAS1knhTjcd2UeXU8bhUOE8eoEVo6IMjP7f+OAEmOSv80kt/Q0eEgqx6sJKdY7UNq4kxhEA
zrnqS9WEGqpZ4yozWqZF341rFfhnvRkKWdyBOG+nI5Tr7pqCPUAx5JGGrGDJAlBqYUtOwbVxYtzj
m7BgKSq/o9xKtoF3TwLRb8NTrvDpOtqQoxk5I00013azKkTtMYBApz3FIDMj2lF61Eu5AQ5i7DVX
dc16KmDR1dyZ0Ry2+xgDsphPZzzxxSJmUABdJXvrpKcmc6OfsgquLVlIg9mfa4bTiD1mVtvNhito
KbwI9cdoW8UC3EFOrhAivkUMX0eq9IZ2L2u/8folrQ78q10jR6iUv582vdIZ6sVamA7iHcks8Ia4
F4L7QYyCVTlRqREiP0VVzY2r9U9ugepgFTq/M66oVTs9mXZo1jx2Mff1t2JLIvZaxP+xITAPfoDF
OMU2o0uTUt/ZjHOZXCJpEpVDDv90ZFx4C8n8acBm5ER8mWbw2ZqjJzoV9AWjpt5iLI8ZUYR4iVCr
Az4wvu/XeP2/Y5f6t6EjjPAT3c061wJx5ZaLTby4xrhffS1PYh81okwGc7YsFyxfa+PjPgJMCR2U
5kAldFaO2c9jPMKjomUjtjEgibd1dbM2017KrTSQ+jwyzqRIB5lRfiu6uZmftLkCD3sIm/OmDI88
gSdA+rJDCJ66MX+NT0qPkaX+FAUmLQ1+iMmkodSlKFUQ/5WvzKnlGxDGCsKDMjFTKX8T/JSb7uiZ
r+xvvZ9s5ul+liD0o48geScFk7NiYVvtcir5KDv7jn6CPqIb5HeUNnarrgncxJloq2EdoWoh0nCK
pFg+wRvhr4F1cKOABrZ3ckvyplxqzsSHbo69yAtQd+Q42OBFDvO0i84h8s9RgjmO5HJlcSmvj6bi
gNnO5jHcWYCf3RUfIxVELHX4xj2cUll7J0BWuIhGPSa0qjGOnwfkrRYOS3T2jf/bDwZO9hcsrXLV
wIigktBhBe3I7lWZNOb4O45lz/5CQPnIFCd8xbXbyt+pfMz/mmT0lc/11UIxXowVPaWQ+DzpdaNu
LISqE5KK41tv0TPaB+L4REeHigpFcTWNta3R6dO1Ajn4cFKoQKBZczEZOSQaBLpB6/ulCoVIo79q
Rn3RyfIwTa60mArZUG727VAOhOs0dAIsTR7VKF+5zPlLy2M8IC1EQVGQGeiDJl/EUJqaAazbDCtC
xSdPe8omzKjlOxvnVjIi8AT3uzu2oGf52RF5kVhxTj2ls2VIT0bfvem0tifqPlKXL+L22A/WaM7V
lXpMURkN7hzUs5nHs8wVusIwyMBeDW61oQue10lbGlBxaRRrEscRu1MgvHl+37MecK8CF0R+GjZu
KC6GmewPLV9r1ctRg+4EJYC8p+Sv9LrafojYRE23mPwsmKBLHwFaeltbf891A6BCnNEN6TYIjJb2
sO6J/g3AtavgXjopMp4DdagHhflCFhkTZm0aK/w1HUX8ypl7RL1dLs9x0BZiQdyKIzCcdnhesngd
mw8gubdqDxG7Ue+Uum+459a4jtcTXydJ5cWIcEQVg11gUTbRpxSn10Id19wMp5vy67cx5gwG3lHH
LJVyqka75C55aBE0iVuAl9bzfuJG6v9hitaugp/eWw9CJqitsv4Y/5hsuI/h/X+jRuXLuK6Hn87d
C719tw9fqZpPH+V0Ln9A8w6wqy/fpyfSCetyIparShM88V+XJQWgPHiA2X7FYH51zsF+VfOR27PG
XEYR4xTHycQ1WP/BOnvcC6HZZtthcr2IdG63GLeG2UeyWR3gdfDRi8yEb7YUOVra+YQ+eVydKyx5
4a6qe97h/2hRYGX2eTHkIgCcKUVhR2xCCRd1QJVUqza2uCmpfymnqtt/t7gVnzYVnNbnq4RtdFij
ZWY1ClYi9k7H+fahljxYLqMdhaDbiWo2fH+F04UTvw0VRHwjEBYZFiohmB4cjXyML+iz+T7ik3hJ
v+kBrmTdP0I849rnkfxZ08MqeYDXnpe84R1u80z00lk7pN70StrUq1nh0q2L4eViP7fMLhDv3LKd
MIlLxt7+00+LoJptOExfLKWcEpreFFKLqrPAaBGqwtnvQUZWEftbwGbzm1fc4kAr9bgLMRiCgaZ2
d7V/GJ3mn/XfKwUL5ra2lPNKgDxOzNidZGCVzl6oSd2r23+AMRtbTjdMZm0knWTvo2tXst7nI+bv
mSKHwSRgJuR1qgrpNSQL1JwN6hBC/fHNvINMWedDSTWvKVSPcH4cMIrBfswDX0vzqWW5ibqWH7Cc
rjmCG0nKQnIrxQX78n3aG2Qo5aK/YgH+BjsX26yysKhtmjFF/u2xsMph8+F9DNbdLMEPif3P8I/y
uuseUb9OLFyP5XPe5HBeRtl81ZSzIpqnS9PeCjYdl+NZT3yUa7V04MEZmtiBdkpPiD5lFeBkU7J7
bca9tksksOKJ2oWMPeyRV7IPREw9HQZJgS5rxtsb2JPYSHk6NxlCzJn1rt37kRzoETcHz/WZI2lj
zjDItEVenDYjbIHdWG9PqxZR+O1/NSgi7NiD/rn3OF+uYXb1UUy/VA2XVXgeX7dTAhIwjhFfdRgh
oRZRH+/GfBnPP+FCHZOM78lOCmco6rvXibJDbTElMJjj0PXmozh6FMD8ucR5kkscxP6VZ3p1F9k3
+LyR1HOZopFaGW7/uuDndfSiY584j/mnaksU+Otz6NE7Y4mBLUfAp2FtnYGVBFFvmCN5uqql41KF
2c0Dy8DQ1hKBWp89gK3YUIaD/6e7KVDhcd3qlOBNA0TQpR0zvytNsXC75pP9aOGUbVlam6JH1PHE
aN2vew/GEhq+ODFzmfVkrsoYhaeA1XHXRMV14qtN/k9299IIkjYHr+cC9HD4vOV/1DqpGVRdOt3j
GJFJfoF+glhzTFkiWZjV32NWZSr9wASs/HkHQpZjL5GWhv3DXFf2zOfUHMkWNTIgIBibXSQEu5tc
HorApzjEJA8XJKPB60xJg+L0wPa+tO6f5Przw+fX/yEw1UXPmxFngmlBGhUszt0UnSRCgaPGvBiC
VwTF+l0o0bSrTSlhl4O509DXcc/W1XDdmbopnaFv27CCPY+nqU/i3qugGvh35VXZhXbtWZrvgJuw
iJz5xBIc3Jp9zT90RzumnN93sIwHhYMFW2uwVTnWV4Oe95AGZtV2hubAVLCYjBjGHusTyeVHXEdz
R1lVuQ1+sm7ZZqlZSL2ibno00Uq6UT3XgohDQmE1qkpprmcKk+sP6T1K37sCgwRDGJYz3JIvCUMT
xqLSdgbyoVxIfMekIl9JW6REVj+ctbbRFBTce8OK/ICAr6Rz/klSsUtekgrr59zwGdV39NlmpElW
JL/g6EucL9AM7ebsNwD425CYFB6UiuKMdfWVwCw15WawsTWglFfRCeqkaJqSubaHsiYS4DaD0VNS
N+6W4PfdHJ8+uYjL9NCdWWdjNTyHh0ZCdc/hVxMcqUvKFCGdUig50hhOqqbPvbAGyqB+lDpKk14z
BWyG2oArscQR4xY0p64fx1oLMwbDhiU3oi3Q/nYu0UEy5NFewJ0yeIsnNRsqSFdfY0qOvbYuyK2S
SHJC8aRiGYysYjUcbSDSQuNTXve2O3bI+OcMImyhC68i/lpbWS634ELr5gethLuOanI8sidclN8O
B+k34KaEJKXpqZQMkrYnbtos4o3BOuzRfTqpRn1ekFoO7tduVcLcC6+tmbmIHhiRb9PoPIEpwixy
uz7bLw/BBPX50eJpXT96lZ3KtSQvBKMP3flmDlsh3MN3eTjqKG/Io6kMEf67JaHTMKsVRO+4f9yO
w2+GDgrafOp8qOAcBAYsVSu7Wi3jl/HuCjTWLMaNUNxK5AXgPsSEw3O3Hn8Ce023v6bWgrVT3SBX
w2Chxi/MnQJB5GOeiBGEpwRCcMG2clsUqiRgPKB6BtpTUO6E3h5hd7Z2UXv6m/TVdXveFtniXfSV
40H3dzljCiw5UO4Zh35npQioSnGd0Y38tn9zJhttZO54Z7WNH2awjo7Q1QuSdMDPAoWQDEhgSZ5M
cXEz9fXD8trjkgFKXgDqIUEgpAb4SKykXYzVUfOHgIgALYC6h5C/RaPdQELREXk9ZThqDps8niXT
HcyZ4PvOVms3MDVBP1ZuMwhsjYR21JuG0sR1ARWzDSiEcT5pSEmw3HATb4ACm7MH/v3VTkU2Tv+I
A9inOfEo5s5Y2IetXpbmVXNK2Eg5VKMhQq8JJJYL7tIsmbDcAoQVsyvGOMeu4uOXSnp9M+gX7w/f
mtv5SbWU8I1kBy+X/GNOfUiJ2cHMhy+XG9SpJj6hwzZnzjDW2qdmULgais6XyNUqnYGKx7veWe5S
8PGdVX004Drob3eDutOt0W2NtDy6FeFVNJMsLfv4iB9bsv5RF13tcY0NZs8GCtiPZ/AMTYLXxyZy
PHIsC2mpETY16XO43f+DMFvifVZyzka9nCMbrw4rbP+asm/B4EA66hdxTMLk3Tb0IzqDLSJ8hU+9
W0QYtuxwlvWfJqDDiNPl5J6qvprunFHruaTE9C3yQ16FW6y/9uQDQ5SpnH3ym3NlrJIgM0RVCOTw
A+q/K2sBn0viI/J1WWomhNtO7iNXwTDBHqq/KvmRONJ0l/pKfnYnibH3DAzU7TRN2xrlquSC9kqq
mTmIFcnAvneGsXkSE7fu5ufdEG3JQutjmBi7/3VGqsRPREY0RO0SyAk63++Ikh3PRf3wI2zk7y+z
0XmfXYGDeZKSISaR4DlJq0oIAnjcNLyRrZoSH19KMwV2+jz/Jh/T2eM40NspyUikNJ8rFa2fhpN4
S0oaARs1w7JZQ3mvQOYGDNOJCG9Xy7urr1Lyxmjud0k7K7LD2vGpHK8tC3XDZB0J2Rqf1LuHpUYr
T1yLCJ7o9c3Sldl774uCEgJa6MedrXK9UY6EFxmVXuwgdNXXgJvTWun87//SwzdOu45uV8gPZv/H
1ts7saKl+cFCjwDts3XEuarZc2XdwO0NLFrYguXrK3Z9v8DyeAtwgcOX3DSZCDW9uahSuVXwlicd
KBh418eFROjEWMUlv3dyY270U9PpOHH5XZV6rHY78KX/s8EYu7YrowhMzlT4dhwXh2g2Cbqx/PON
rV8YfjZ8tG47CzgJYsOSTzJXbVvVxlozv8lbby5so9GqnKddeK0MgPRszee9TVHO8r2LF6GVMJ5T
etEt3FHyI9LmVJGULMB23m3bc2VgRZc+DbOyKgX74w0q9qJr9cp423VyQ6TO34bceR+Q+PUchcLq
Zkb2En4lxM0b4ECpzdsJwtngHSG+tiFx9p1fF2hgtD+1Wc0KQTiTnWRoxyMLD0kkcmQQW70TM96e
DOMNF5areKdV4IKIIcs++gdGbbfubhCpRVhswIc6A/HxzyEv7ubaUmKy9MOsS2CPHcrPCsz+Ze0s
D2UD9854wRS7/53lm6CRxdDG3cp5Wi84oedEZJVHNPvLxtIzxzC6C2uW3mbOybmHnVp5JCp6r9dv
Pnx4rPYSwL/yrbR63UOIq0vLPBCUn04SHY+fVbizr3ZGY95fnXSKLBhXOqLqsw+K1fJ9uLsvgiuB
HBnoFsQQhyexXCwOpMTz6OD7RoDNz4L/S9geCQ50UWQ5K510w+LjhYJISjo0ZADu760bKvfY9DOv
PXUviBO+4cJvqCA5yQI/HgRlGRKsbIqsGPg4qulEeaHa2WOzS+MFWG7jxhDBF57X+zBb+h+T3EGY
dzQtMQSqWxlG8O3a/aUW2ptBCF2ZB9O7Vykz0w9opvP2bQKmsh8O9nzr5jWJAWXhyCzEWKIdLng2
Eb8oNznP6o7SRyYzvrGb6YHq4GlYyRWlhfpY4yecGPUJF9YTfv36JlIN8PVh0RI8D+TgzcN3A9/4
RYopFhg3PHgkz3B5CtfLC3FMdCt392o4Xl/q8ZOSx4c/fDvFj5csvIgLkUZnLApaA6Y4TbTRWxXs
lMCm6wT7PVxcGKnWF8hFR/Yj2Xr8lWAcJV1XlkxocUwMd0+ZtXAFoQNGfrcz20vzhYt5xm38jhAA
2m461YhrZB9Gb22foL4rk+wzfw5augE4CIpBiazPKrvIMYvhz+41pX9YZg7AEHg5MLt5PsF/GeB0
sZfHVkPG8a1jMaC9zYfa2fowQibdwmlIpxsr2+b3ZsuErk7DAc9/aps/rwJWw5R3VC4/1/iC2Ejy
NJYHa/UwAvjscxuY9CS0nofApN05RC79Oots5z7QEgNKW2vkRVKOpQZhqRvqgWbI9seRMS7xJmtV
rmcJdHwg2AXElTi6qMIEOKW5/1vljVonqfk+mj7F7F8G5uUj2o2KrJKGV5SzzpQ7Cy0OKVT/oKKI
qrh5Cb2SepHr5SqI41/9cps2qtYziuPO13GBPGEKWUbuQL0kqDj5xe9aSiTWhqQICNN+NBu1z6Ix
grWiojvqr/1hu3crKfAfObUTqKi1ZGtZ0hNUj7vjv3V+J5otCXql5UsmvYna3owF7SJPVTzgPJ3q
bOWSx2VSuUsZVpW+isPqVjwFmPZs6S67Lmwhxowxj8u+7KGKXjxIl00avfBK+Y5xfRZfXXPKF5H5
pl0nN0qxMi2PaARamNcnV324v8Ksi7xPtWo64+Qkm/r4ZaPJw8sjfZXSq1aImwuk6dpw6QRj7NhJ
b/U6x8wGCGFSKuMxKC0Ou9dOYP6AodhcjcTazMweQNhyTv7CpEM3D/kVe1Egw2Zu6Bv2+fjl0R4o
c16oPHeRHpKowL87BhN4P46fjUMgdB01MTktM0uKTaywxDRDmlebawXQKEm0KlbcqYvlNweD3+nK
pToAKVfqjNjEVm6gEm6pFk8//nxOxamQ4nkOQPMFe9lrMjA65hRmjlrpYHEqhNESirj0iwUs6ZeF
S7mEuwEcMFYyuKm9OWSpvNs5GBaCSTpMQ/sCJs3RCIhlLEb+x+e4TL2RBBIcRf7VKCNauz5NZ5Po
hwYE+G8YehGwaSjDnzztBPygyDcRDevediY1vn9jzAnQFZagKKWVjYQH+cyowq/APk0oDI7ZIsey
UnspwAsBY1i062Qh7EmItFR920hvLCZb+1IiewY8RRBhHGWB4agORY/qOsg6wwnoOlcyVMBQo5z+
pCCYntL51bPUjFOb5zf7P9NbjEhxsOnJBrTTAifzamwqFc0W/o7rRCI+9uxqJSuaPsl9WPlOhGMU
Aai4PxBTCt5IvwRed/5aDsmdHjP6NHVdkpYDIy2YHXfYktk4x7G+Gog1+o4E+PICQo21gzENe9ka
EmulFdCQsilYnjNyuDl4L0KJTxcPfp9uyPbEHwH9xLHGMQRshyML7UOxShPdd7FLTWkefF0vRaPg
VDm4el/P3FuJIsI24w2CeByGZKlh5Ps24qIdP9AtBUW0LzigQW58OgaZOEiIY9U4dX3rJyC5trnC
vtI3jT+UJDycDHO+uV8FGl79uSzRbz9vEO8hXpjBw9T6aZGXt1RcvyELX3ovchasj8rxpzG3wwbu
g79ZiOuzw8Yg6/wRSGvuDji67NosGZ2ecNQ7ScEpM3BNkfPtaM6epffwVxSUANoT+AL+dcsMuFKX
27YxyfROnkTgM2ZacAxMIvhl/PrIBelIN5hPgIvEEWpzOfLK07bu3a4iV7ySiWoCMa+515XHQsJ6
SG35kk3rCaVVCbi8+5Nz9sJNdLYkgqmzs6u8h+ihrhX2JQW1a9waBvXYW6ZH7IiZfJ4qm72UcaT4
s2YirZ1BrkMWu4U9F9EqYMH4a2IngDP3ZnQeEKYUYS+JtJigQIUn/PfuwrCcCdW2vXaJzUC0HgY6
vzVIXaDTeuy5hvU+UpHyLxAGHNuQHOoCDMbQHMSJTRqC1oqg28ieGHkWlZbXVVPuagfIJxx91xY8
2WH99Qd3ZnzKVR8+/WbgFxvxIcTVKKUgcYZ1PNydzD8ZNPcLRzD2C4igUb6pW+NlkUJRtOWUA7OZ
lxNRIvdR2IanvHuaRiTGHA8ZlVewZdBiy8Vb/JeQ8SR7ZuPHfMx5jdXt+EAKnpSx4Ke4E8EYV4gB
3Erugz0JcpAkG21x+4B1cuDrLr87xMJSGuB8oTiBf/3e5sFGVa9vxANrhqN5fnILa61yc8uzkJSz
CV1JtPt3lFBzwcXx6mkgtn53MzbIE9vP/6i0yfELIQxGIj428/GHKXuU9tahrr+t7RHL9Vk+X7k2
+TfSS/r2nm3BuC1NmmmzOG7348sDf7tc4MX6g8Gkmbfd3jN/P0BJ+7+iTpsaJVW6w+CNPeeNW3h5
OhoYGlmctXe7bqbnkFjmqjSXnYDF5awwx5gTG86U6g3G9mI98LHuEgHNvS6OpveoND356TQ1aBoQ
JfiSKtaYJPbWudkf3U0dX2dDg7YPFUSej0xi54g4TkSMPh5SnsNhGbtK85IhFgzelWuTbuytshQR
H921Z/+x6vYBTbdfSjCNiHOdAimh6UbmozMMhtZKgjwSOCjXmKnH4yAGZJHSM2vC4bJ1lh1AfeOr
1uPMel/IBCKpE/fSsFREbM51HQz9t2YkQVP1CRr7N+Q/gHYxzTTl+/B9MBWuxSfawlN34SyJEkQ7
vjkLGKP+RTBRAhs10ux+C4Eh7++QkLtEO2WedVKiCvcEW8ReoBeTiHmSZO8SbjrSNEiF9JQXaHCh
y+bvugOyv21jCWrFlQfd0Pl0mwsR2O5JWFs565yjO+Z75O+0rSdYFILmvVsCEPHZRHsUZ6Jn+DYx
OIfo5KTPzp6dLL7lHTFT0TndM3+wy5Q8VdvV6zFpu5sx/14QBtrIif2Ev9knO1gmnUydZrdyc2mX
x7QUflh0MW/YsPGhKfF56CD9Y3dAApLn9n0VnoZ5xVoKAjWCpC2JUlRYDhgxJVHCyhZs1RqNEs9K
6hEuNgH3bEzfZDj2pUjHJA627LM6AahaPgszfS5kTr9k2kYaFWvvtMtAG1i85KhiErs9Afq+Pt8Z
I+tueajZXnLKIpHXa4T0rLAuLNeKp3AySI4r+yxaSWUr3QWis5qFhZVmHbCip3swCLp8T9sTdAmv
tav4g+EEcOJHgG6lO3EQevqDLpJWZUxJ3UCrq2M2sKXUbf1KP8u2TYE76pg/QvnxyBXpwfDbVY1g
H7MEuDv8SstLe3pcZ/zxafmxlZOC6fai7KtLb0BuxdBlMTX8EYaEK1vY6yguq9eLNMktCmxxRYCZ
anhVzkY/QntpRK1M+sl7cpGT54DvJfvdV4u0Q7jIpa+4/JLXqW/b4YhH0N9+ZFHOIKBE1ox/KWCA
2NaoTbwB5BD9PIVsCRHv82uqIOq7fTkwbVinL2ZQcq74nohhzrlagjRXGpMFNACvpTwC10MD61M/
8L+mGaXNS5X03kWV+tNjQ8EWZtnDnskZNc8KFm4x4upOT4/xtbsenvjdoel8JwfxeFmoNmn2bjW/
3v2ICMK4MaDBHNPVo3r53/+I2g8cbyjJdx9pz7nCPcyqgPGR4mlS9Xgyj6fjuupf0zlaR6JDVNYU
YvnNt9eH5NI/i1T4N64OOnOVOSzOSnd2IY6OHuXtBP5J/ls4GnKjP7jyvfJsCNAB4+g1+BITZi+J
0HFwJm9vkyM3vYP/ir9TWAJiqlkI2tUijIllxelZi0/tQCGGexFv1UrS1jenBnus+RXFc9toItXV
w7KYQ2ETPKeVBX2uNe0/1CUGBMlEDrn1iSLaWg4sm1CmhVnkcFKlg1wmFSsX8B8CO+8eJVMhAgWL
G5gbwk8nfIH/RT0qBvxa0MQeoCw4nRSg3CtpolsXJ5RLW1cdimSWwbIjCkS8qPmpFGcVBZCoHjAI
qLGJlwufWothMaYesUv1k33XDQIVQB4ZMQ2r8vMN9ud2uP0CXiycvE9If6m+mSlzIHW9EOYU+42m
RuQ067zgboQq74zGE0XPWhGW9Yn/1cxeadsWRhDy0iDz4zgwkFg/zIht+RQeXe/qe4dTLZ+9YJER
HWXggjbZrfTdbs9FO6SRg4Te0FGARTz7Ah7TPvby+SqiAZacw0uNu//8pPFiX8VdJMDr0SulVm7Z
f2svVUSLnIzSHANS2F+3poZFQfJJ7PVp34kJJFWp73MsCGmqHGFQy6wD02eUA0qwMVgCSlAMnXkF
goSNX5smOg4Cj5Iv7yPdqL5Jcvz1nfTTgB+oOn3n4ufNbjtuJZxSdPwAFFvl1FxAOgOsnd9tdApm
N6FfMn/JfWgVNSb4T03LiS23J73Vs83iaRYhPOR0wLvsL3SDmnCYVWdVYW1V4LlPICkpzw8tCAB1
y97Jnwh8/RL3LBNBwK28KJkIeOwtfH4GwrHT2Gbw5liWuAZEV5yeJFGWskyl9UWuVSJqmE/lf3i3
3+G4lGo+hm5Ace+RAy26+XxHjvYo4zWZbAJqmZp6oBJ02ntR/eTTWEXWPXuoXsKSQ7m7jr11Z0CG
X1HWD4bn5fTniBdnc5gp2+ta9Q9Yh0BEjm7+ZZuQz1VlAIQluPte+TEKADgNIVNoEArjj74icxCM
ZfN/4aL8C/qkRj1dxD3ZvzB6mjp1dB0t+I/pnaBqMuyKlvt08MBjVbM0srCk4bNBvCeTRdtmTC4l
+vYnXjpyjx8786JD+OIe5dOXz/UBXDIc+SOXvfIVPn+tLWDSh9iU7xHif65BijQJPtQKOlI67hKj
7mdPLz74c26xxKi9WjagyEChHbEG8GEyE80spCqbYUtg7TZ1b6g8nsdjoY6RZSFynZ9d4tzBukrx
7y6tldahihLXOyAQOhvlK/QfTIiKotRjOv/+XRRZxZDB0MnCCJhKVe/hq+8S59bR6oobeGyVwFTY
XQIRPE5q/5DfrwRvSXrhs+yp4xEfe+7m/QRwKqNkz/r56HN2+DVq5aUZ/dVt/zoQqfgb72Trrwya
+I6cxTBN0y2zwZ9JAA1cO0n8MrfjtnWMLFU2pNa5Q1zhuECLMNiKIK6kweyJLYAgQlXNDdzHT1jA
G/mXaC+D7AOX9Qx/ngX6xB8g13ORXIpVu0ekTG35IOuzGtkWxmLmlcjglx7x2Y2rcjDRhVTlYOQT
xKNC34YvYq6EyII2QOBe9aSJz1wf5YGBqYRD3AyIMX5NoOOTaPMeqdoAoiNybVqj0JqkJOqRu60b
nrW4Rk2F5HZMztdu05Xa92XZRSQrYn93HWd2TMqLsvYA4/pVjjaSGsEBEq2irkwkTpw7qTd8YAXR
9B7G53bIlcWbIj5xG8lmTdBC9sw2VntMvT+TpGvR/bX3AG/uw5i+IAHpEWYMoYY4BU47mFI8OO/P
ytKAl1Ope/Ndzv8wtIVD1DpBRxOjB8LoonOLgkL6J8EFhNix/PVwvSfdStrdj3rCXHOhpEd+aeVV
Y825uDrcf8huutp8Ys33RbCAqfyNbO/C6hwJK921PFw4x/u542lrdlZPiusYhqBHcIfT3QiHvuBX
KUF5owz7N4TEtyLLJCqjWVPJZ5F0T94h3DPtn9QGDUDA+re5FDBo6Wxyp6rrxDnawtGAIrED4pwJ
6keCFjapr3XXE4+I2d9MZW+1Ci3mDBz+LN04nlngcwWb7NIrQvO5riYuNJQgEZJt+l05z8cBuLfI
cyHcRLwCU/MbVppXF73C08g0LWBvzjcGolHzybCLvPjI12TCKHYEXUiscdaGJxGfe0hMMuDGjgy1
95Ij7EdzMJ89g/gjr+cZi8izfQXSS5fTnAvVZnn+bUUvrdx1j3oVqAQYgGr01cf9RfEdBRkDWS2w
YokauQaxjevaXxJWP6s//J8HenXwqiQiVHvogGv8sv7wMIXBbIXkqxezVYTRNd6g21GsxhtXeC4m
VZmZoGZnV39hYAjlxurMrOh5/KC6zD0qCC7WNEnsKaYcc/d4xBrIW9ljMLtdNXMK6Z8xnMtFj5dD
tXoDJ3jigUYUem3JU6OPZdsptH6mujWE9OybbiHDi64K/QN+8PXrX/gHj4Kcl7EcE/isak3FFDJ+
onbZ4zDPlDORy3OcPqOYMtGbv2CAyUSFcyByxlttR7bZrfPSu0SHufwiQ/7RfeHUw22yxV8KEleE
4yVOP8v/7h11gVoP1DIVed5QrlM1x6lqenBOZLUr9JHx4I9W9A27X/UDp++Lf5VMCVYFjM7GXd/Q
afBNt4aP8fF3/3eD/wnNN2fAtDpsR2koLyQT+/jsLh9IBufr6eraQGQG3FBhMllKxfbER+zK5ir4
hLxlrPx8u2XuEU8LPELMyUHmpn0Pz6Ha5B2L1kxZI3fG/OzJxs5g5I+AABiojILaHlwQNc9kYKrz
NhZ7LLoh2UNqAKziDJzwnCNy/bV2W+SkrCPfvE9i2rRa3lZAdw3HS7BJu36ger4NS1o2ZYoP8YuC
iq2M93oOPAe2mLGjM/ziRTeXnN7UIH2MetoZShMsi80QC3tyiIWNRQo13hQ2Bby06D2qoZZnsTf4
V0Vz1wSvvwUi9Fw8+x4V277/0rfx3DziXr0tM2G3tq019N1M4+99e6ECeL6mIB6+FIYYIHH4Xl5f
JwTum3/XKnP62rM07OyArwXzSLuEbB9VFAnxrW2/zgKe5XoTn0ViPv2Eb2sdJh7RlrIp+jcknpRT
Ibv8gnyErMqlC0TvrrbnwFo9kfcPBBO5OXnG3jYGYgk69HDImI33+kmYiBGSzhEXoKgvcOvlQt5j
fKjFp2llTkFOuzYGX5qcDwZyLQo44gCOJK1kytGHGRZmGmUIIdN6VCGlqz4qaOZ98ISjwM1QS7MD
/CB29zTeaFDS5FBGOennuMowuL3YhERXM79APDqpl6M/7JvIfquH0OgnWvuoakoMfNcaMbrw5B2c
OJWYCK4anLR9YYB1B80QNZE5uABP9tvnoVhQlHZPj+GuQGNrvZRPsXPuch33mb4vVFMuGbo3NQQZ
VkhUT3J8CPwf8SFmI7RJdTCTwbCBxNQFgJvjQNrliGrIius7WaWIAA40x9NRUndxmimkf5WKS8HQ
cMYA8U5MLSvcQAd/rz8ce5tm7IEnRtgKhLquUycokGrQ469jqaw6d7hGFONNYBP8CYevjxDT1rA1
pyxw1q5rrPduTjjMs8nQpN4hhgKz55a8+JxLk6R9LglAW3qwchK4AvZHL/JCxkUIeJzMLuOx14nc
edyrG1r0dJPIY2XMrAZ3L7ysi1MglooEtvopTsHxyJBR2P901lHj0DJtZ+PkefYmrwsNVFin76NL
l7U/5ne0E/WLq9ff1nD3WQ1GSTakHCoL30dqTfwvZSqY3E2K66iC08ytzhUxPKBmtG8ezu09EOFs
5BcjPgnWTx0FcL+q6UqWyuMZpOrrpiIlWFUkSqK4csqQVXInBZflSjrV6BTJgxkUMRQ94kZ0BlEU
+LoGkIqFDzL0vKMpyaBm9geeaWGCQUGTgoh1n5GOGSv8pONd/BMB4n91bY0IkokPlU0BpXbikdbr
8wfy/lsVCSBs8+FIPUatHAXYbUe1we6GhvTNlNxWnn61zd9/rGVNB9SfcokF0lHmcKmlM0jHmwUt
3A7YarwGCJ0l2xUc7u+OaRPyH/uSdptsyD1X9tFx/sgRbEMDY8wKYAWrfTC8xw7aE7l88WhjyyiK
HnIsYTVm+uY+tx4dXG+EG3dIRuN1zQUAqBrvTNVA1pfoo8YEfYvzHAvWp+qpWcpl1+6Z4XvbLqc9
0GUCyTY44np8tgyezxfV5Av0RlQ3y8ZVMuucMupIe7qsUXEpR+5cNeWHCxzkecNRTelXreLly2kK
t+PwrmPAS6O1Hve2swrncxMI8MO4IxbtHn7GJD9pT3mw2BukjyE+wf9vXgPsAQq+BIdGs27hOcip
YMX2+CXsyDPUpfYty526efR+cka8AGyxNL0Fu+HdLlIMdmfasOytDne0TbIpCm5TaifhSjZJh26w
m8vPAEvSc8+U4VYh8qAxp/D5Iv2t/65ABEr4MoN8DCTDujC8kNlBlhIqsFOR5k+WIJAR+137BMbG
jkGaw91DsZPMIV98xE8lkw6hfrKwDGxZb13wSj6Melb8iI87wqF9JS7GVgCYz3HhfJI4fOcKZAvK
XDderg5ref1srSh8yiLC1/O7Lq+XdS1QeAqH5PEqECKq2oN91InWauv5vQKNJwPgEn71BSihI/Km
2AwFRYtReSAzMouu/TeoyUoTEK/dV01Ee+PSsYSG7Ko8aWWXM3ubbzi704gIDiuTWBaX+6/JjKfA
VfrZbbGOWtQ3vb5WCPJuFDXAcCMstDBSKOjNulsmwKYGHKFzEwuk6/amhD/t0oADOBVcKKXqF4R+
aTUCbgrutFyJ3pjr+vzNyMXhj2J7AawoJqgRUxDSoE23enJNwVND7JHec2UzuIzw/BRxB/pY/1Os
CCZ1bbnOFehRbPI23gCS1oQHT8eVqKYmTnffAahnbNJTJY05UsoUhZRL9QfPATJf6X9tyEFl8pkr
VFz0I+UXSktMZ9PBh4VqsO3tQ2QqPYcpygBsZR3sPavLCvsKVdApxmc6COkHqDryX4MJOnilIhGh
UMJJgLfPjWrntmsE0cgH9MLL6pOY3x/fi/o9XPwg0IJdfgacLxwaNKM3TRAFQaY2GykVmf+qjDUS
Gr2XlkELOz7DcwPdlqC8ySpYv336oZWa6FG+twAR4PQUDJLlroU1QV1EM49vbWpDbVWKNbMlwlRe
Pwze+L+JqpwhkKxdJC21mW5VKpl4lXWFSxj0W+fQs99sX270mmb+YeeU8GKgYvWB4e+MxxszeEeb
un2qGUCGaPGlwmQFTBnD2YKr1Wk4wjMT3TbCFrdDjnkuisuilSTGSdki+kPnkxn3bvHsbZjQCBd5
2+kU+6laxAScRwVxtOwinH+fLAHdyOJJVkGwoxv78eT2HaosG1gwfqRqm6WMORJ6ZRIXWzxWt6kB
1SaE1A9BczOJtZi/qG/0T77bw/yXeCaRSWYoWRsGK+4LffU1FRL0/x5RS//lFYlc6UTHoQFqgvSM
d5yHzwzWyZhth1KSKL9j51ukCBpWtzoAAHGYV0WZnUCuqvy0UF1JDjLv4+tzzB4XeOvG59eu2lZi
bfl7Whfk32Bk1pVThoLjPgd6fQhUjaSHhqKGUGRLhT5XAat6jVgtmVga9tBTYjNP8ZcgMGkeJ2jg
+SJ8u9+8BrfncrJ4Sc3nRChnnUyBTZczP/o6KSNO8q0MVdXX5bV+mvepZpWrzebl5A3PV0wTHLh8
elk5TC3JdqgyLJXr/HtrSnNtjgOeZWspb3NND5p7xgzgUZSpmteN+04yw3KqWv/S/BeCwOEz9wOp
80W5xpFaKX4IYuJQM9q8hYTuQA5nG+yKvIzEjZcyC0YZ8X9kJubNpAGqIResguRUAGpgUEqDm6vF
U3gWqECHp/pxMUbzoz0gb1njOuGJM2T8/mM/Hlhb2uIvx2+ZeTCL2+2/9Q3iAIsXvT1y2HGSvHkP
vmauX2xmcRn/5l2rcDb798bIq1uQ40s5hflFY/GAdj8CvJqQVC9bC7sfsMvCQ5sdCXSzZcYGp9hv
QPPoAdX1eHlfxbvRtzEBD7tIRcYMbbpqiJG+D7losgLdabcuugAhBDZ1mEGcAhe4gW7DL6m3lpGv
SASO9Eev3WLd9RR76TncpVTboBzKziIM1hcf97R1UXOTguq96m49M8TQDi5wvlwlO/vWREErwFMX
1BoshVJwO9lJFp0dBp4UsmCy236XXoO2p4uoApU+sr7hbSVyDa8FGbbVtJELoC6vM9kJjYe0Fbs5
wsFp5TS/b5gcU+CYuTHmtmVlSjpcH1q4kbFxodQ+jtrncsm2syZnh0zMEoS3YNgPwHOVmzowVRYZ
8znjH5n8fOsgYEBFPUS+uzN3U/S/Kaplwhom8XE5OmGf5iRyK2c+vGqhICzMUiWWSw2oy13XhH/q
J76PSud/Hbet73SRBl2uQyo9TDSdKV7oaaLeZtaCoYt7uGTCstRtSCSDcCSCrn9ak30IAPlYEtTY
xuSufTn9+JLUGtagDmuuN/J5Y44OAsHvSZu1OJd96KpCgZUBuMR5/O6eRg0b0QAxeanthUOAsKg5
Zr+MBBFhDMo1mtpfIsin/22Ia3lYvomvX08u0fFvTz5aCkFr+HXG2D1OHWIUuVj4Gee0Cfa48K1e
hKM37PC80ROx3eqTbpeT7AKrbdM+NesNNIOoeGq9/OOEUAorMLW/Xv7zQt7foQZKTH3Z3tTils5h
/+DqVzkikt13q4Iyor2cva1KEAly7krxPMx0STvgl/O14JO2c/t5ahf7x4uiFn2WxuYmHOnLGnfb
zcaK21p+EcDhK4E4/Jyrs6O7JqHR7i34hKegmt0KGhboqdXEtQgzO9rbn/QIEapMyEHltL87cZh4
s1JtrFdIte/SYJxsdkLur5GZQkip4LbNoMbaOQ2ciFteh8J+NUEP8fYFWSYxOgtFU9oRqXrdcLtb
IxzOf/mtQWYIiPFAEsSZgl9w+vtY1PmsUltKRtebpdCf2mZoxmu8qfRVW1vN0/N62CAKsGjmIGzn
QMEwVqlLb9BiG1HxMDhGIx6nRMNl2y0lz26UoxZhHSelMe2jX1EqJdeaLSvQkp6znrwWcJpWJxxP
jU7lLjROxboAELQyqMc5q3OQxXA92eDiMKYG9HGXFglNTIsrCuJtTx7WhO+177pNOkIdQlnDsgFQ
kMui9aCKq8X/kevkZGLSxMIYc9hjMth2dL7yPOvzAKhGyFJ4zSdjLkFRQ0ZHL/S70rmE02mNPPBK
jrglA1YSafSRuAbu+7hzl9zLhxNAzXRmrOJjwVVFBdLUKOUhmJvHOQmvPOIIEwXqgj6xkGrwqtfl
4Iet9qoKiIEFYBPmlhQdpMHm88txM8nObtqIy7Zxy0QWnpK0/aXgCu/hPGWLJkT/N7ZTiODl2Fkh
4YeocjertUZCk9GwIqERsT9p2YT8mQb3nlogv0C5eoHMBkKfKyXwPDVi5Ns93RWgnB3LEaG5FR/3
R4QrceXwNDRoQSVSdnneHeBIpcXV8/Z7+mEvIJVkjJ1reRvt3Kam8MCcFJb0z+ihWmtR48QKFxZ+
PbC8cy6tqaCopBlRopA25J71mkmiemr1VY2gW14C5ntyk2JTRmD4zNLXHzDY0C7U52ipE2pvDTym
I85zKXZg0bCR++MBU9gsbcr6koYsX/O97QoNTp8smRz1w0EqHvyHZ9U3wwmfyYBredmEXG4xW/HY
X00jTmpKqVsjRpaqXu4p8tl/75cvPe799L++Pr8X7hCLtR2dlpdlOSkchwZ7NfCyfgeuV+Abz5pL
ArQ1iyQy4prWzWVz/6K5McQeP9+2ypby/Jx1y6JJy7oRzwNCm1odscjy5kO5WWEJfJb+4Tc4feAL
v6VMXJiVhm44F6lRVKG8cbxRvhvtWod1YssNhcrxF6LxMmnyHHYoCFZ2UveF8pR02+mVtzz7DXE+
bNXm2WNSmV4tZciWjF7UnqYhncuV0vA/GAT9NohLO1gW+vft9XN+tv2hWBj/d2goXVDd2IjsuCyj
Ed7Yx1mM2vCm4dfvyXv+25SwAIBLeQX1KBufkdA7YCJ3p1WOLlPBh5nTnvbQJkQCbExYlyK0Vx2f
slC3tyZOsK34LacweMTQ7ERMCCszZFYn4vh3HVOMC9h713FStk7HKnnrrtrbrKAdzeyL8N7iD/N5
DgbL78IffXaYuWX1ODj556sOFyIwScMa0rxa7UwRSqjgRBkcI/7hvSbRaV7U/JnUfRxkH9powRYu
6mhSr+sXPsGAPiCb9f3MfMRp4qZoo6pQ61Ers/kONsyrFU5HSFwqdgUifqlO/scyWZMo37OByhq6
8LYD7g8ib92esLe1Ffkna/D/eLALJGhOzLbLh919eeYlKUpLB3ZCO3MNS7WdB5YFVZLAjjMhz/0M
uFcdBrq7yD22+fjSANfSZFWK0HG2eNRlE/ZAjsQOCCbbHbSFWngcFqHPp9Hx3eL+TiHpshwt9MxA
ZU1Uz+aWglEHzjda7tAswKLGDTe9ABt0npmP7yzhHizWR2XOmVH5GHChVEihAbpKM+F/eY7Rb5j3
XhXAZ3ajZY30gVnURaDxEnG4ai6ZhMDCNJ1nvjvIIah01TB8Ua0Sd9mNwORPPAt8ABE03dw06C4F
wz+3pH4fl0wgNNzTBU0ovNadj3NzxNwUQuwVuIjS7L0+OyJg5UM30yGY3uuY52b2P/ZvtG6tX6UR
gtw4WrOQGEmmuPlrM02edlBim2BgbKebpc0IeNfp6sTeY03ocgEv++I+fspFgwCAWfWo851Ifc8/
rBznhI9cGUTkG2ONORY9gHEqwNrSue/zVvtgzM/XdaFt/feqmhmVKvprz4sMnrSmYQMvtDAtDz5i
7ajEzts7ad8rM9d/PSn6rBZTjKm6ZKz+7BveRLLEdHNG3jn7sPhNsztl8TbRLhhgBA2WPhQ4nhNu
kq8A3cBT7knGvf2jvB7qDw9ribQ32DxG/buK9UI1dbKvmG0NFLGlBwPqti0+GbezJZmTI8wD5wxd
dxuHCk8v9Dkez+DFV8WsR7iICE3CVHAW+VRn2EZhNS6GXRK4HjMduPsoy0HU6a9XMcF3mTjZIxM9
JbAcy4kFCfyDWMYm4ZVHUyEPekKmr7IHVxQgM6/arKuwKfFdY0J+pK7Z1WC8ba5lL4iyglifzEkO
vU5EFK7Jam46/vWfxIhp0FtaPJahAbIbLj+Ui/O/s6hp1UxYF5ZsQRcjAyFVS+Zm+SLzgwwJ9p1S
PXC6zvUDl7N3wbqEaL2qyo11pkgMphWR7NRQH/JfAr54GsdbPvr8hFfnI5atES1ay0O8s62s7CQq
8RjTdcCail9wbtE/WYDlJ2gZ/mgR+GQ6dUp7FoUnY4Y01pc3JqQlAkxpa8oeTLFAPFeDorwGs0Mz
C4oLUYbiZZ5gBeLUkuMB2BVUG+fee7WMz1naBzfPr4EKz+PUlrZvKDkm0E1nJYQLs5hRjVaTMOrD
wqT2oMKvg8WGwS8EN8+tKk+DBejKdCu88A1kBRnlTcdharvCsAaMJoIRZ+0M+3uSHBTtf2lJ04cQ
N5ev4ViFtwXeVfMCfqDIS9GdAjJXIe5TMVipUAd8xxCoqRb+TCQD2X3jH/d52GCi+8LdlAEQpoAD
+CXTpBMT2QlQIMF78ptPCwqYWFeSSfb5xGAaX+56kc5TKCa4XdoApt+N4DLKzFjx9wvybpMC97mQ
4/YbdjfAnSvtMSkgWNvjebt5dS6ReV+isjBSDaUnjLZwlDhsBgPB60pl9P6w5uRK4TSx/iLD8aZM
uuHHZzVvqS/bixCutjh/f1syWciiczP9AhKH2UxkgCQh8UMZGZlLEfx2q/1QKHXNrLKBJeT2rrDc
M4N3wCGkMrkOHCah/xKlCQ3dDr4a9sfV/c2tjZlswMqQGxhBbxJ14HYE6xCrHzjvMWTH95RGyc41
KGEom0/4xepRevhePfQsnNedceWXuFVvX5JpK3Mr6wH2jccpoAs9OIUtUhnt06THE9itNiyMMM5d
eYE4tPoEeoHM4loKlrt1Jk4PzGkBSMC34yUJLWMnPiPHsod0uIuKx9TASOl6gONZ96RiNILIG5Kd
175puzsHCNYX2sYT98T3MDAXKNY5VPMDvmrTgCuFowtZe+GkleNtgEp4OnxLgfLFxTIaJeuGQz3P
X9p6IvDNB94eVD8fqbO3ajb3niWB0V9sEMTK5izktXo6QHVv83g1PGvcGJBwSiVirI5vlEr7cKgb
HJO4bZ1484EVddFzMExgKJrbvkTjFY8r5AHwdpr7ZHHzPyCUL3yApLoGzvsmxvwZn+m6z2ubc3Ab
EIiLAJGvIfK5hw76Tp6nefM5LSpGLK0JJfKxMv0W4F+h7OOO44Yjei8DFENaasoZFKIxYUjLb7t5
c5CoqxiLwKSRO0sbfLdmn59MhVKk8K7osihMr5OrTyb7XNFxSVApUKzy3rOMPLbSh6tC21C3hzzV
kFVLEGHpUfd7EmefmbbR2EqhxgEkDXQB33Bb8IcnGocnc4zzUGbnXxO9erSCPjI+vAXK/cG2cr0b
+6K++a1UC8gOa0XbPpiv3xBXlTSC7iGue3XL9i5GucB3/Q4Rw8eo7TuHBzLrm2Gmg4rixfhwQyjA
ZO+eGz4XXEXYquxWqOHDFW9Nc9WdUn8Ekzjw0+Es252ncDZRaiKVor4mJM4xgbdi+Wx8cRtu7EEL
Jyis6D0wN/MYDxUUK5zYSOsMXo/9RkVqgu32jm8dBJKrHVFTk6eZpLR/PbDJnovoUrYNXQpXWaN+
lLdq3s4Uyy7Fh6KaOdRMgmUs60a3ZLJyW6pbZH4Fus/WEOPB5y3y34kvHbhSx931pMVNrRPRrjOP
8Kl7j/8WhGwApEgNPfhphCr1ynq3Rx9U/AKtJPx2XLUvbiMotP/lx3MJfJAzrp3LdzyBscywPGhK
oboYe4/iS/zA45vB3R0/2QiaUZ2pIPqmUtRe4N3q5ioPD7HjRR/VPmsS1qDeKeusbW6x2w8N+PbK
DVH3YvInEtfruad1p46kWPHRweTGJBfihW73wZNpKsWvvG2plv6mYAA952Tc4aJ6aAlBkjKdJTcY
OuxeJI+SyTQJaY6xQc4daXspLDKWDv0W/cLoXkEPTUtNNBSWn1veWfe0p4ldmL36aGAVqz3jPppN
AvcP1rOIHGMS4NLKN+DEzv2nL/ZYSXl2qhL6GCaxz7v2J80LhXuKAI1XLmMBqAJVOz0uKGfx3jP5
AHbPtY8JqGhq/e052FUdqNSX8D/aHKm5AtmOpkiw/MCCBLrkAGc4jT55AKi6/mtptglZg5mrcFLX
7hXoyJDHjD06joig2Bws6xkixfv3dXW4G9XZ5hV/RA1MNVWfH5KSt3ZJaSt9EOtuXRKN2XVlqNX+
TPsfovuYyay3Sx0qY0bcLAsxSxFVJ2SYRbEK3XbAVLE7A34wXkdgyWBu1s+RzYS7oP7ky6xtvqNy
EfoelpzGSFTMfK0qGdyZEwxybDLAdkx+hZIToqM2Lv+0D+kSMaOxo0/85uGVbEB9OOUEJw9fAjzE
Zpn5us8FmkBG+yERnFu5f2b+g/T/uCCMNRKjyVVmmImT0IA5Hunz+44bfRzoL2+MPdAyC8WBjTgi
iKObfqKX1SluyCoNyDuVbU0TM4PhmZkgnlnW1zomD19x+Fg4hveFluyug/9hgsv5gc9f7EdHoVtr
hb4Qub8ytx79gBV2af8ciaZ4MnUQltYdVQybaagpUM95zaETjqVFfW5OT7uCUzeAHCdmX5vC2/ZI
caIHu57eqbg8A4u1fP5njU5w74JP526zdS0QEvrweCP6BJI7qpC8keZ1jjQa/Z1TIfQc1EC7MEme
65tfwWEcZ5KlrrtzCEKZJW0JN8c3lG3CSOFtU9WS8jcmk0jpaWfb/JshVFMOt1h4nhgxQa1i+Y+U
wteAstbkiqekmkYErVSPJ2dV/QKTSRLhbNLt3d/kJzFiCtLkpCEUgn0OtG6NFRGed7y4SH/jPu2O
svQqL45WnbxZfNbXeJp0PHT9F1dx2GOLVQ3Yy+Jb1lgx4ZK6SYGN46dFhXwxFtiFqExqwqTwOQMh
U3rpIDDx0+4oZDMqkoaprs2a07GSN/7B/McLQ3j0a9u++4mfn71Gb8VGUz1V0j5P2NcpiSAriMRh
9SEn5JbCddHLqM398jqwBTBcIx2q5DupXvoIiuQ9x8VQrxAygvN3l4csXMoX2gF2zEHEmHEFK2GD
/iBd8x0AvVh1aiPm6Gf451Rsuv+Edbpqf/vwe4jeRF9iRpIjFwIfACCl3eHqZ1YfEeHcHeyurb4V
fUb+ONFGKj1n8eoJ4opQQgxpjarWB+9BHp0l0qqPvPacredktjt8ZGtb4TsATLSEPW3w9HdG3CJ5
KCm8sIK60D7uyRW+fwOgU+wbzuW4AGWwvKBw7+eNfyd8ZeKGZOyUOf/WVWcPQq1jdidokgI40pLx
WoxMlPAkT5ehXc8rmw417AlT8ziu8ULAXUO08jw+M+6dotzhiD+arKDu6hEQOGF5t6fBQ1+Sj1Hl
arrT+6KF5UkLpyFthumxUrhnDcgDuMSW93S+gv8n2l/mbBJfZfmdvKSS3v9hLa9mI+iZ0pETSyEM
i6KOAlgniDYLJSJrPllYQuPDQ59tB11Zv3GKrtD1Es5q0ms9VsP7SknBwT+yBsNb2m9ra48oOEIc
d7ngfWuc6IRWNzlm7fVBWvVshXUBo0uex0ud+vNBB43/HWgB7lU6tKFw4Bm7jN5pz0RAHxiKMjBV
ZpqDN2OgPSoj7SzEjnmaRvfxJFIu7KXLrcTOfm7HDFRO4dOcKmPkm3nFg4NaQO4McllPVJygS0Tc
HtU8420ZtLz2+N5CYQ9RO+X4evaQ0fd6gIR+2q89VtlRnbjJBez6DT2WIhiyz1gMGDy4rcwM7c/O
kHO6Ptu+Z6ApV5PTaQi83MqNEN4ZwWDRrMPcsjpJnLxaczTlOUjOz4aC1WpSP+fOCMJ439fUiLmO
o9ZkxP0Vo1Pw54C3J2+BFpW5euoJUREfrU6hpFnP83LIMXqjEgw8NSzKvKAJleft8/ncA7m3RdBS
TxAtEfjhLO58KOX14Y23Nw1eXvUMLd24p2HUGubs9xzlaNT+cM+NCTUvA87D7Tfn8sUZGxun2Ftl
+U/J86RIAU/Sl9TIEY0FmxA3ZPWml/dZ5+X1DlAvYs+69twj2SLAp/1RdHXEGk9dSOw1vxf+zqxS
HCkiRrsAL/gb4HbZvCCntVb2N9lh3w4d1of2ppBn9nu+V6wMOFwbMvU9nCcatsbrCNqse20b5UD3
kOP8VPibdpXGo1vBI6Nn0JmiH24z658vuzzNINbsjqpMeh9tt6qbkKByMXggDs726Z7R4dm5BOJt
MbT5ONoNuy6v6OqxpW5Y4fP9ycDolCjj+2NEZNh6GraCej43WVnqmM1RzoTQ7rHv3CwyWQnq6lD4
nxoeZ7NJuUMTNGHZ5+FoZWPv9eypSHI1N7/dAJBcP+tm4lUgUG4UcnId1q5UjFKKz0VZ2k88m/xA
Kk4jij/DIbHFLX9CvDoG93a166qqBiqvN5WPmRHd0sRazWGnfyOrx+1vAUnpPjziio5DDGhDOmcE
f9BN7KC0PglYOgmUY+UrGw8EnG2LqMGP5Ijm8BsCBjYy26Q3mPTJ0hDqWN60ETrr3RMmRXroIIb4
V6617kre/sMb9Txi2D3jf4JrKX3ZLVQX+6B9BcLOpy+cszbqhCIuBSpMAsH9aKsxrisq9dOeGSr5
qGxBKIv23UxDQN6GzFYrRZxZIs8i9zSB3WDN7oVJyWQ8opdQ832XgxoNKJgnW6y+LVrUyw9pFXqF
9Kj534nxtReIegWQ7KGlcdMI2HHphiLcwhD7enppCzSQBeky0bsI2bTuCPmtOsHdml2mUpHaTZlz
vm5DWyehuG+0NuBrYFBL+hovaYz9UfMGUOCIHJSBcCu4bk1t2edo2fI52IAslb8dJrbF4uaER8s0
Q1G/7YmLjt1QuzRcjX8dt0Rc29SrT+VmIICaibu+LbESe2v4ZbQP9I7lyjmZu0XM7HWRbAkpsLOj
hmCOM/NcGUn9N0XZ34OpDz9JRXlWyJFpKZuxtxE38fVWaLbbgzFcZbpwCiQ0g1+lmVEAp8Hr30w0
tqjCMRjcjph+JzDFAUDmjuY1r4ba7y7KKLaibcxNTgw8IG4csp9eaiVcLsdYi6GebxTPHvG+qyd4
SzTIMEitvyaiBidDFDRrbdtKwnFuWJIFjjRdS+yP9ggMoWrMCtIvaSbjKEKxTW61DICzDY36SHy+
5TYMOmF/5PAaRVBUY9aX8k87AjHKWgOMzS5NgisQCMYvRddnbBimGnoWvfeApXhjeG2cN/75eTSE
Uf5KujcqthqUVgji+xwJpAI07dJVgn9F3MTZMgwFNgLYHNVV8gFCzM0RBb02Ofd01q935qkPwjbV
l0lvvT5GbNk+0T1WLO4vgKjuvWPCt8HvkH7ljUHV7tOYQwlIVtroQucDgeF+o2MjkWg6lIE5j4+Z
gXp0wBgvH+TVHm3TVv0UrkYKG/fro+RaLW8LIBlMsJE3OkQUAqHvs5mIGM7dpK9Zs+FjlAUYZ7G7
nY9PDERghLJEgimmr2o8cJQ3DMwVNXTxnPEKz05u3e9tAN8VY9FVDlqB/+PKcTqXhEc00Tz2/BKB
h8LTm1QVYehBETkSoYfDLo+OKrVM1z9Xd4+474jmP4T68zKyRHhniFC0gxqo2P7BMSXF16SRLzUa
oLaOcIBa19b6Uz6yjGfla7wTpkfdmAOypzmWPZaZ65qIBMyJeJC1FV+HOH6hjqUkeHlOS+cxnOOQ
3U1XzFquid8YIWdIZbrCAWiBSrX7CgAzI1HRqzGeFXUlFGzdJezzsjqrr4Wn35zszErc4apThiIN
CBXg9i25jfGE1oPT7VmuGwGdDiSRGlnuA85Yw4ZQw7S6pIKu+oqlM0OfN3mxOT2l1AqnswzCDhtT
4kdVM89GSR7xBVGn0U4HTQSts6gT36Q2sYncMtFJeVJDsAxqcZllgf0odmOurJjsWLM/GIGyGm1L
Yn0LczuV2LjomaG6hvK/yu9lBIc9znpdTQpJya7g++J+9M7ygGJU1KwXwhes6CXhKiqYvHQ2KFhB
deKFECMId53cPWO9xdUPpBlp68l8TaT2Yq3by+88c6ltRMk7AhaZmd7nbDZUxePekuPSE3uotTGC
iZiY6wDHBLfdi59UJ5XG7YPi9nu+pyPIL/BvCbam2NEXCvvP55iBFmzy4uryetl5lJ09ID27kEI9
acJYthVdK/xJbuWrapWFCGsa4iXbaQHL2jVGgaGrHC3opkbqLvXNGXaYYAKl/DIowJEAXBcKjc8D
CX3zTnfBgUVPt1AaVQTSa/Isu5M9FvuT2CIeMaKbkzF9DATJgD0d2XTk9A8bZdNJBLU+daIAoyuH
d/NRRJkcRBPji6goRFs48SAJiAqgHK3yePicxk1Tkq2TicEKguOCyajMju/GyXXiRfNPOYbNZHQs
UaIfd+txEcty+PXJvDrEyW69xUEOE0bIRMD6Rb3pyaJQvGvWqSdaxIuYbReSNrOfkIPjDHgN/B6f
zsGgdhVhgqW7Gy00RupcVfF4uNziyIqP/DBLALo+ZxLYOnEApxkNhJDd0YUGmo1hp/B8etHxnBEV
+pezcmz4aEnM1lL9obc73aOx5RqEjlh95MREpTlpFR+Liaa2/lvJCDoVSLf3ikwXuVFmV39LtYVb
nkZElDKjwsChCNEw/NYyRJdwD9iTAsaSvqLwZWSMX5zik09pmKyqWeghif2PauifK/DtxdFaUP4l
nQT/WnrLq3Iq+5TyR8RqMm3VoW5pBAt3Ac3eXlyBsMpJqRl+0aw1Txj1FDxNECvu1KAnG18skZFj
lAeJTkkpTOxoMIBnrnKx3h2b5kXyAb6HQOtFgNLLfrZNHYa9sxrIyphK0hEWpw+/DDORhg5iAdJZ
uwR3F1alcpdIu1j37+Mx3bIeVRYzZ1PrwRVZ8xZi0oE2RPxC6CUw27q4dxhEVsD+omzDxQSH5/nd
PfjzWHZt/q3GIJyPXCG67n62oqdwt1rDaZBVmQ9j4lUtg0fyC6DGAFPtUDlXswXPdzXBhnuX4LQr
iDrm3Wh4vOXvWB30Q2ABAMB+faqON8aEU0/SwqhS8ru+2dLWjDpGP5OVDBOYbl1T58LbveZRZ9kt
HMTbqZsKEDmErul5eYufCkPddMhgZOhNc9x1xXNP1ecxi+DkqwTX7OCLFPfpeDeLrhmdNk5ZYA3k
heBTALKZ0+mpxMpQnBlkKXP1SocvheDao9TdiSz1UclD9R820vOE9m8jpZHnnytZa3lslHwt22RI
Zw1g3ER8cPLzEgMWl511xWRpGJmhYVgJSrZvmwBmIHDAUdkopv0Q5BV6DaGgsF04PpXUREYDYCLD
soqg+AQh+mrtMsKX3MzVEgBKsKu2DW9EPLSJwdXD2JnPLK1OepR++8J6QUfwYX2wrpVnNtCYDhke
QyYULuU2o+vQ15tRFeTulj4x9BPcqYRBWIUUZXIfY2L2SMxNc7shHxsdba/iCKcR03RY83bVEP/r
TXg2l/p2gDda7HVpcgdF1QSRRvpL1n0C26akgxh5Bccb364glNaTgAB6Q6ScgszmZz+/jKt7FEsp
J2qhv+fLSApmAqO4NdB54VWBZ9uebRc6bmpkEJskc4RkJI4NKNyHHqDn2pFy2c0uSYjkA2G7GUM9
IkIURt/BhCcIosrQ77C4HuSqb50I6nsQFbCDVGoZe8GcBce9Jk51I+iYEMIvaT3eqqEIRHKkIl2o
KJcf9LuWzvHwUjTUeb6NzeGmcTTJf8NDI2jBt5iW4538wJrCgzKKhvf9cNtvjBL8iskWc4NZ7icA
FsKxyIEQsGDqTJUHBb3XvdmO9Hnd9WmxpZVFl1LFr5NRVwYBS/iUFTh6X7GM4DWNPRCThNP4GhO/
O1TTczLHCpEAAK/QO63DryeHIHAiU664Kw4olq6siYyfz8B2ArLHiYjh6iRGLPu9kr69DBQYt8xy
XzrC0DrZtOPFHkMPDZ0rHWXn9O3H2c0vNBRd+SLh7mqXRiYPjTBskXfgsgCDexpk3jEGqCkEjrx/
r5rcT36YEaqZLdpqaRAl1wGIwnLA502yQ+xe9gjeXMgZeLvJox+puo2Y1LsgxC36ouI5ZnAAz0C1
qKz2+ygpdSSxwaWsKvAEJMetXoI3iyTvTe7VVqnulrIEbdWtY9ksF0fAylIuojMCJ2vF6zDKPjQq
+aXPVCmY6xb1m5hrLyh/lb7aqNmApu2AQSt/BHSDa+EoNxELqZ4ObLF/Y/+H56+TTnewuUxWC3Lj
WxZHoMCPTaNjzgXwRu7kxnhnFFbXr7eBipn/noo4K5+wo88agYluVs8avKSpQUNfmVsgAk40++h8
5ysdyaGXhs84MeOtKW4p9Ig6MEXthz/m2eQWiGESsF57AhBpjoX+vpMfkHLgIbuYuHxEUh2y0BvO
8aeBkuSVmR3vKUE/vNKeFnGVTb8hTl10m5f9dILBqpOI3QWFf2HtcEUsgJ/MtwbyxbWXEW19sMkU
xEoZgeqtx4j3xBSpOz33oKzVKmbPVKYdkx0aFgzyBVl46sIw65ENvvH65mHVSzofn5zQb+ZNnPXJ
e6omDT/pW9w45BgH5mN5PZa0QZuDhoplsc+io78aBFuZElLfnALmY2i0obC7oyMldmcKJavEQLFK
I5LHKaCixFuHKmDLGFTIdJjC7S3Dc56QvP3sBjyWOkeG43m2ZkHCnwHJ3dKTbabgGGMNX3xusWcP
sg+n5BElnJ7FoXMAUVTZw6GsvvKcpI7ueQm9NLmEjb8fzbdvs41JTZqWiatIXbjQg8fGsGCqv48L
UFB9AGl8ZkzDLFXTBFPTL4eJZjdkb1C5gAEX5Pi3+OJmjygC+XHW2KKS/93EbGvN9Ui/MPFSMwPm
W51AxkLBt9x25HPbV940LFZqzc3mHVb7iuGY6xSy2aDyZoQVrmnkq5c2/VDTp4Bac/+cdXsP8GaF
ZCciwQa5Mw7RdvwD2KmbgpfzucyeI1Dpqv1w/2jgFmKwG8cPe3pJaqwFfgmcnBgFquLD18OhdxIs
mnrNXX1px5dVDGIjZNG21G4d2uwcL24Xn3aWHpm/xiTSgILDvc4EcnrRi9pqj5rDd2gnKQhXakT2
ku06s1lEZ7eKiei9iRKCCPAf67s1jhppluEyiql22cZG40kcnn4Eu1aVh90c2CXKdOyLhDRWGdIY
+BT6tGm+p8y3i6aqdi64mHA6q2DKdPFi3bp/UmgS2oImxVuZ/J0TZQM9gK6nawG5jMacHOh1tn2H
phDxfWiuj9iXfrVC51u2YBm/WX2r1axSfk0VSMj2E2hAjApxmdyWV86JxH9Bt7EFt3BDwXsX0yxJ
P4buQhcTog1dzKq4Dnre3QgRyY4RDNDV63Ju35OqQkY+N7Yb0Czw3ZrdIFyASdvFV65iNcytrAio
9NSAwL5LuDQWxh3vmdrbxMrgC34kDh5/WI41lw++pqlni75MvLHU1RsL8helXJtZZU4Co/FPrh1v
EsEdp1U/PpW1pJxhk8KVxetJA/59SRRt4PGNUA8DTh7J9cEclNa/E4QuvMm/66cDWxCKjONJ6HLq
GYa1Ao8uNbKkT1jElOTJDk68l23dtWyjcVW1zFnIKkfikcAlutf6D5FbJ6/h+ERz4D1Wq4lClnpl
AbDCOw48l5HRi0K8ZovRsEYxawn7HuDLpdjXREgJIz37mut7VrXhABuEdMoRElKrAFG/Fwbglu+Y
bpQM7Vr1GrPYAhhTQ+57aBzKdYE7Hn3TKdm6GLTxdE9nTrXBgtupqBAq9zwS/NSS0KhZFh1CKtnw
wYVqWvN+PfmRVaVQPPts2sdn7ieldG0IJPOvj+qiRRp5qiUnVbarBspLSjqixgpRA9B8d5i1dl8g
gND2nLSX1cthdAfwUCOdWNutiWVWsprEDaBUgs/VWXX6OQKGFstx8cbeGjgyiq/jEsnRl852MmFa
o0cpTAMRYawoVK8zf5G82+derwYTIqppAuEsi+ZkruS51ZOYjANVkQsgc09KHaIFRyg1YUImnCXQ
VvYaStvCEJfWa4DjUpael9xrsOSPL0iVwC7h5SvVg0C1gCDKxi4SpV3TXPk6NQ4931VZ8+mwNHjo
IQbG5fNVYXmxwXIHd7d8fBX4FDffYVyx345oHYuqwulWjqykS7/gEZO4GwyGPkrGUjG93eboMISc
ZyQ7ZzAZerJBuZjTUc3KGkWNiLagrD1HP4zboSH4fhuyfPAH06I0OA2Qt/l36MMIx2R7Dd6gnhHg
PcN/1WjOXEZxdzoDuTSj9XA/X0YsbRncALyRoYDIrk0gqFveIRGcl8TYrOBmbRv+cTakCQtqCMJb
BJn9ogkUCcAN7ixgvkpQOp0SP2HZynCc+aAwTu3KsFaI8W95ItWmym4mrCmXELSpTi712pQ3tARF
fq1K0PqTmypSXqITtawyf5/srSlsfCuY6JQg7bSoZbmX/kmhZd3D2XIAoHOUZ5McT46JH6AbDPxX
7CPs3bIf78gWJ8lRGzdlLBu1H4C5YtA9zRHOSvRKTvZxiwBERArBn6eHlQzL2iH+7ZomqyELiLtc
An6HdMxINMet+4qL24Ql9EQ9k85PV04M9RbzRTousbozKw7lKAdVvnirS3Tb/Oi0uHP4FKzQtTlM
R54IyNuk5tBOo6ULs3tksMk8tqz3bHhYVZnx8lsJHQDxwDKvVW0JyNIqhc2nwnmywzMb2qEDfhP7
d0p4L5nRgjpCyl1PDX9CbikjgzmqGxY+X4n4UwaICRsSs99BDgs/4W26sbGEJ0eXXdIFE+Lhk7Lo
kex35mD3O3ZEXXXTbXwqQdZs8jsJBCldbbJH8MRrWc8KUJPrhjRQbtE8+XAz5vvwdeqanVa6mZOj
cFpVU0o5L9I6tw/RkB4R3BU/5EfUL1Y46h1Dh6e51lSb7LaBochLTde9ukSlAg02i2xemg/+2goA
pw2sEOEU8cABYM+a0Mnpw1BLtEEAip5/r1eJfawwO9t1vN7hiuxvSrC6VdFj3dktoKLorrExhIrJ
FrSF9u8TQmC6QgV4eoQEBIZ9fhMJluLcMjZSoAHe9L3JfWDpKP77dm0fiBSv6PA9DDq8x1mLq1FI
nLUsyzUggzmca8PJscJV7gE2jiJ0iY7v6uxqK9ZYrmoZzETjo0ccIpovhkJmf2hH65Sy9jxMZsi+
p2GoyDFHWlBXnjH/Ix3G625boEZOfi+hQ6EN7hBfLgSt0ljDWEfzpDtvFNOvxVans0617OUAnmiM
gAo0fvpTE/yF5UzjcqJxYxgWNBlFP1a7O0ETRh6BquzePss617Rr6BYoZxngnz+fGfXZHCcoCcpf
7gfk3sY9aCgo9TzACKgJ1VhK+ylgy610ZUWGPVVZkUeOWR/abCnHYD7fcOZi4PSnl/cTbfmbWnI8
7rO5r4nqYBdpC8104xojAHSENdoaoG/0sd64ULiXSutuJC5x1GcnWYUS+AVWMJFEn+iFQ9h40Tnk
6AqoSNJOzMw4ZWWPCUBSRM12ZXkVXqNAKTZfCYWt4YY/hCnO5pmgkF0IwCcKJe9bBCQAq4gm3lQ8
gg1It0eKjut4LfS7UnaiO4zGHn7hCaj0PYUkJJx7xTXgGdFXNJYrBa902xwuRgPjBPchiTamtG/p
ZRAD4Y/J0jz0QlvEJhtbVb8C5GMIJEzOWHOeOz/TLghC5BjvNX2RL/IpubKeoFAhdlbUg28KLz6W
DWQU+796BTI4q7TF9jRrJ7tD3VW56t2HxzsW9ljMzGfRnZVDe2H2FFd1h1zOGJ6QKGyEBEEfkvak
8CN74p31JtbyUPFdN5HbonZy0ZvrX1yyEnNRVJnMT+czZdj362eSwV8GoFd2MkCwvFk+qDNtFXA4
tplApzsQIyELJIYRJR0LL1L2lDiDsPRro/Iy/zEuN88u12otLWnE7V39Q45laBtuYKXp+TfEjNPM
KSSAdTgcVPnBQ/PGZrMfOarzriSrpDTVn9XqJbc90dbYqpaDtvSWXOMlyCoGX2tuYzDDVcB4CH/e
65d5iyhluCdYpraRXWpSL2oUe2WpOc/XwLkG52rN58iya4KYFT4ZkVrZakyM9cizJcvRZ0EFicGU
LLy0wKkihulRWVaPnn/MS6ZEyWGPhxvnluDhnaXzqIVybW1shzUs2f7IC7hvSy/UQ6LnqbOKBC/G
Pv97kv79giaxFE/acZn69rB1aDvZH998z4+QQ2ftSCeJ6RkDJeCT7PL++oINpGg53K2K6vupMFv1
KllnwhR8aG/ZK06j790Zc+GQsgG+ZCzQf3xdJZdBHV1krW01QvToqk8MMuWh1JEfI2VaQKGs763N
ocEOJgVqrlHGJjrYwf9DwTOsQckxWGhGGzkclQqtIapLx/BQC+XUlhmWG+LAJIaEBpp39y9EbEuo
7o03GmexWy4O/BaIqfCKhPwXVKH2FBRc1jZSTdXVy2x0FGgjScxEyv7mfQFJe3cWrDdfCPD5Vv7P
78PUNCshWIAr+GJa12f74qgSRcwwwF3goiq5+fi1NQUFJcWSxDksB4WBDawP/yEJEjTrbHhEDQi2
vp0c+3hFPySz0WRWU+ylwLe2gm2f2bzzqEVzju7R9R5a4PKN3XxbOCR20Qo30r3yP24onHBat/RM
Mcu+bMzqVCCzRoTm0FTAkZMUHFMhIm5jqJ7DyJwsO8jVZ6s9v1k+GfhkPTRk7SVNDO+vhpZozXE3
5682viqRqNv1qnb1uxgfPTOkIqe1vuVF8MA9EYq/gnRpLWxyMBLx7jPUsBlp8Hws/wWhCyyZcv2m
nwcuyNZdzalkzXs7ZZ0Qm3gNig5yQ6b22pBU9cbLp1f4yYmWyMht2NEkaSCCD4yMz6pkGe6irRSj
HyifMsEWurQ7eHpqR62v1HSweBaXeYrNlS5PNhs11cRXdvxd2+8WUHABrSJoemGJANoANRJIL7V4
VyvPcQiBnwMPrkNf2A3RSpRlrLfoiJK6r5smi0WGevoB9CfvZm22wf6eqfcC28Ir35z/e83DrKiY
O/nudVRT0YCYYJYyV8OkqPz/b+6d+Gi3NWn/5uIyTY105vzBCZ8ZegzKiFxolu+NRPTAME5X7tNt
TpRJxQKZPabvWfc8WwqEEfW8L0q4ftXWR4wff0luskys7WQNRLKaSCNDuk0Nl6wcQ0LOGc4wcWQw
uLeUgL/kIs8EG2FD7X3N0cFP3CTkD19JQDDdk6GI55BausW+bIBBxeVBckYF23cTqDzVavqfZ8tN
p/3yCtAgmK/LxjlYTgjLGCUX1r29Mn+DeFFi4w54PxUwGySpmcfjxxwirEahzA01w0pMFFUxRGYl
C1sNiRLMGSYYuKl1bnO27Fj1HnuI9liDfhEj6mdDTyk3qi0rU4k2FMJisL+1YFXgP6ePM4xV069O
tMCNCp1QyJQpTBfB6X+20MRbfvm1Xr7x3aKFvlkGNzxe+VZbvVleWqnCfWwqu2yTpctrGaNBXcJ/
Hoa0nF83XMy+UK7ZHpaiqltq4z/qa3DjHoct3DJL5qw3+1Hl+VlUn5La4MHjSWUljNqFEbQlJiBb
Spc6Sba9NwLFVXiURNjujskf2Z5PPC3O8i0VCd63RCnNBVZl8pyX4CYvziF3cfyRkyWx2DGXJL+I
xwUQn+QPrZ/NvVAGHkknRVj5/yd1fWeWaUWdKxQWobfeushVBQ/JJK9M70daPn9DgkvFNaccV8Qj
BppXl/n9mZIvx5FWxUU6V1Jl9l/0C/clT1C9cVeOgcmdR/0A/DUaqdffLyGstm52sOZF4frZGbtu
xIWtOM0fiKY+nD/fDUkx/IMgv/KSyEEX5zyQsgnOWMjqo1vm2PobE2j8VBVPh+3p/NSqZWiO+GDz
wfgcPdJpkAXoehzv8F/ZdFtRERZmSd+b8CrRgNNTrUgJqLjq3+3+gNZVMXA7jAMwkSWqY5+aYP8p
Wl/Y7SlJYCTZle3ndGP+eagq0aAgoKyiuIEa62ILYJ6J7I+EANJbkW4jtFObpMdU1kJA2YwJUzEG
WoekMexun9NU3KT/VJIue28AJbWbolmqLkRLCK8BCv0gnuexPhrn38DGuyfGcrutyBjlY/dTjW9e
miVOgDVfninGT8ltH1774O+mxx+DQ8JHr0jEtH3irDYbpvBoc0M1xdKBDCQx2FFWwsi6L0bXRTLH
kqqjIto1IA0U4itcr5VhRRpYMjpOTjWaQgurWU5frkkUA/QZ7TUFT6me4zRkI2oXIv6F93sh+EFn
Y1E3nxn+Xff27R5LgBe2zNqDOO+fa11aOHmN8w24zDdH4L9bm/Xl8oCuND8Zs9mBqrdRhQg6OTrE
IidKFfgw+WGGYNb8l+k7Pcx4jus9hb+Ih+03xaHFSbPrdWUNrOvJiZB3cUCIhGPy5bKob/Zsbi5g
JetYSpw5AzmZmAxLRhyIfe4fsETL4TW3I9vcgazDYxfp6JiMKFxrvX1degXTKQYv2JAWNKe/6p9b
0v2nYuXzYcE4qYy3jAXQZn/Sid0pHl1Ws3EMAOMqrcgtWxRPH6Jt0HxOGNsISkiAFNvYLDEFsSj4
zY9ZK9PtVYSliIBTDPhA+n2U/+/Tt2gGSTeiERz68PEHYKFPGUxzCI9heVlP1MSD9lkITYeBZDA8
VO2bToWYNjnuoEUQPrngaaP1GtQPEWU2ixHUvVfH5GTlhWeV4GrbrEnxJUogcbgTSnxBVzbQT2PR
kd/cjKk30rbhIobwhtN6+G+e4pw5nB+tUuTpGh+yuxAbpeQXCY+U655J20Hv67nBICyLSdNjhJb6
aOJdNzJ+t7BnRGYbuizXRFqlSJRTAoFysih5EGjRwF5w/Jmo1LQ1WMggNV2R2XDeYlf0e603txWM
M/Rn3vXoUIbPMpS6esvVzC9wTkLsDmSTBhGAbe64Fnii/FQ7ScXCQndFDhbeMa0gN0Wmw0hTU8l7
MdK5CX8mGd+0bcVs2w4zbAQMMR7t6rRHB1qPzc143Es3wHArfkRb+lM3rV1TyJAVCZ3PZoWsXT5w
4qOpRGEbyrNppAzAojg7wCreSVe+2V/gRv1kHqZs40nmoQCr2q0aH8iowxQ/Sxw2XyEOx3qzCM8n
Y06d2QI5xMDQ1Kt9zdCVVpP0Zk/+fmI9RsWNblPg6FfhGmLC5toSYel0p1BCKBDAJHjKsOrABG4+
eqU14zG9NkTA8wu1EO695WagwiqV0EqLfZsSqk2zgQnG4B3qmp+SI5cPLCiexqSevI9BKKuOLvtf
ouaZTwjm4gm3CxWXRqhHgRl6FGGpYqFpJIunEYBAgd2m1Cx8y6/7/6rr5Am0c3rkqyM3Zod9aSB3
SZUjSKcD3WmxPa4jk3RAWf3bik8eJrDUmxGJyC7sCg10uOKubXAeu86BEkJS8oPtlc7Z+drmO2zs
soxFLoFRBeAsbmnLiHRIp+E+CrLv3VC3qMvQo37CcIjZzPmJEP2FZnHlecjMLuaJxLcu3fO95iPX
7xh9JXLHDunq1D0zeBb5iC8rQAVSjx0C/OPVJhodNS65PvnfprI8JZyGGg1ZCn+Gir6h0tbaURjw
fL7uxfPZD8llXxZqYFeuZUmFaCZ03xnjjsKYFQMH0zwPZWxWovZ+nj7/Ri31niEx3bnCnoFJJ5qC
MlLF3xLKW6LBnq6M1M5tiiaABEhzM8LFlKX1rFYcifMEEOexbfnTBEtDmc0n+ZGIxOgRUWANuEtk
4HTzXVkW1ikf/rGjX84plr9f3ll5VAfmglmjL0nlkZPWq4xpt3/tgkb/WEhsUInfEXbYgYqSCVZF
Vgv2/nmfe6XzK/4YImIU88cQoZQlOV7hy36ffWenXBB+KqvEjnPPuQM1iYk0UjtLeNo9W9FFFoOr
z/H96sKLSEagt4YezdTireqnH+h+oNFKvjSEXn5711qnULZXH99I6PWp3bNhCvVL5tXsA8BWGUwn
xRYOx9Qnrr744GH9mhtRnpLosyBO53rRVvb8CfwxUf3uOSqcWTl1YErt1PE+wGcieYUqXVC2ELOz
Ymc8JuVgGHRyGWAWlYC9VwIh2PE9wwvhtJpAUExa+mAByDQWJvLvH5FjSWE37U1CT8HlayKUnN2G
cx+iNrxFGN7rKjpGbtfc85lhfme8/uxbmK5cOSyjJi7wolQn8M7KGt5sif0nos+6N1TVSp8PyxsR
X8n+AeN9E4KMjwpk5UNEHKN7Cd/cf0tI3/HSTR22WO1FOubGv+2vG9ClTrrYMV9SVOcZgYElRQ2W
0BpHxRiNn8vgxpec6RB1KZov0Cq6lhFX6Ppzz/ycnzuFrMJXA8RYVEpEi2Ai+1nrGkI/TRAq7zRZ
5ibg63H9diwOMBqnvxkl+N746oEcalkzF1RXAnLcGStsvW9MxKF0m2t5EmfFAP4PuZt9h1Tbp/mx
/C+nBfIlog9ERuXmnHvJ04eshTu0anaVFJYh8XZaisWgpdytfiq50HmBig03ez+trABZunz4JZ1L
snRkUwrK4TDzMJsUQaQNl89HHeX1KZATdD6cy6HF1tx/N658gR/7rOa9Y/cB+AQch6f+vb015T/+
ghLUfeVB3p/3rfZo6mu7TCJC1aO8QVAAkflSySSTM1S2atQDQbcaZMLqDnmz3pO76rCKA8BFymZb
LrkMpfr4jhvVMInuCPowBBiiqq7qr9WgBKJvXnRjQbnRSm6QqCHPRSUDleQduze0W0hruY8axguD
acINtZt8gKIrud3Va6rwNOxkxzwxIOnM3PviwPnl/pFfFfEdH7N2h9FMrQp85EB9JqX9spbo0s6a
VfVeWuFHHKoon8BN1ztK3DqH/lTHbPTUEpmeXIBC38yQ4ucqvBaaACHxSRTNKJb+zcAJUByhggRD
dmq2PmAGOa1yoznva9wN9wxw0X8qDnI3S/H9Op8ansbe87RLse0W7DYGKYFqD+dO7a/FOAlau9HI
elvbNQxwKeAOb2iqUotqYGPwqeqvpo3mvOSyYYdKSGBf5nI+Z9vObz39x68oLqUFp9a62vZXUlKt
iKZtFMSKCqH7bWiLmafpGKywZj84SDa5Ka60rrOmoMw5WMtAr+hEhBnLwkqtO8B48964owzgcckh
bfM0izRwi5OPBC6T32f80R68saAtqW17TkWnoWu2JTEx4Ir3GTFcXKqJ7sk++USfpHBlhNcj1wmi
l9fp/FtC6TPCSZyScIMWrqp6Y1wvH07E2ig/QTLX+tRQK901zE9gyVzfkpqtvKciK5c/LvQTi0JW
ML0HWPi2K7JYr64robX5Db5xqkXyJfkDijB92eVjrGOwgClWJD9QR6EesWH8vSONytEvW0lItMPb
mygohi+s5uJ4V7C7TQyeDZHagjpMTjoVueZ8jwgyTSZYuTNhr17YnBar4MBRiJMBADsrbLCGSIWB
XSX6jrpQocq3wiKP0VfjGUAijjH/sVoCDmd7v6E45w9E52dVfQ8/8TUNKMsTg5r8/RlfUUPZeUGs
7GhkqDj6FbFNuSMQ29yGKozucZW47CmV8OWKcO8elnKkSklEYsN4gHCTGEfLSufy8S5eCLX6TsyT
i/Uf8eVva+fB8REPZ4qzhBVQcEhGfZN8e61YGCJUXQAmmsYKoeiPnn70BZqY+4bN+eiLVP0EBAwg
62ZM4ZxVMavrykSjo2teV+LG0GegPgCxEFGj2R5fzaju6EmFFKPAKpLtmqTgMOwox6e3v474aZ56
V5ruKT5l4IbKLJBHu1Ocote4/gHcn65xdXi+dVDUlHGRPR/VDooqRCQagvL26devutxmfFsP4FHO
AV3N9M/LdxNhtoFlZDily+Cm608OWfYvuy4tDeX8sDVP24gJZaFV6FKwWXEnlkvgzSHAxOO91jGZ
ZenZXTiKWmPD3Ckpnx15VLGbhCipNrbzM1iKaNNLDdMYH25OUQnjPrV8Lj74KpQkmB35guwfGkIr
SIRL41ewmYQUE9/c63/Vz+g+TMXMvyWUB+Lzj01pE5snLTEpxoomLwf9JAbu5qbpybxanFtuf/ww
2tDAvOP8Ly5eUMAs6Dd8nPTexwVi6d0u7heXenP9pHL6nbbEj22udIUOgl1vknFNrW8eGaZAdB+D
p8n7HJ295ratTvP40D5aumDpwF9lwbogHhlrhARHK120cPzLmVIG4ukNgfCRPyvHA/BQVwyMX8XM
r6IKnoW6URDDPeYThD8OjX3MpX64/TtWllWZ0Q9ssVSEPQu7cXZOgfdMYrFjmuci8md0OlHqhnU8
2CnZMB6ubh2SNgkfJYuj6YpBu6ooEfTko11AND22/r5fUID3eQzo1GjYDfMHb28gFkDhFg6Lhqdp
hfRi1JTBBtFscIEjenN6mmxwvuxb9fN9MtDYxw+9zUX6u2Q2ytyLxwy8ODEJ6O3B4SAsIQmXehDj
FzCtfJbGqT8OiZlIKSUsmkvSQd6YKMOTuyyllEMBP5tg0qnIpv+HWBIj1bXdc0VZp8e/pN4mwkd4
J1IqIOutgdYwZ2xUe8yW3zSHB5Y1gNhIfT1YcP6dEaAUqORajGTX1BQAiKycAU+fvhZyZnJqmPcZ
8qXyyMXS+5jShxz8iTDMWz58QZQ4pcOdLQCKFE/znNdkxxEPQ0c6RY+RvY+RM4rKHn9czu8HEfLI
GBXITTV5XfDTi7uikig3WyTq1k2Rhb7wo3PNTvMkECtKVwiQYKBlnT9H8gLwGHVr1xl793XFcn/w
6BlhmpRfqY+D3YPgQ4u0jcaQASU2cvE16eSV8BpQBQ10jqtsihtszutQdpWHT6tlySaeM9540Xq8
nYAfuMLdaU8NWytaKc8fxIsQSsIJFHRcatV0coR22Jlfyi4NDs4x4jTfYR+ODM8/puDHnCu4Tq+Y
oB9xk8M4Cww8/rGS4nNiGu8YzyVkhDVC2yozuc5bfC7s1ki9SGNWg5kUyoExcfcVLHXUrKQ8ACOw
BiPqvWEPwvz0+t1zT0SlFcOg0ZZ3RpIwQO9Yb+HAKd2x/fY+AI+qGU+ftMfb5NnROX4HNgxi3+XW
nK9iaisAIMJawRMMnJE+Ldu8JH5HWmWIPrsEEFmQqp6/N1c8lElyJgVxKJmHWZSJ4dMI6qZ+53oy
rPaTPD65W4LmnQSNWAv5oOBA6OiRnaVdSqhzzf9OeGcp+On7xpJTI8IADzfYuf46KmmguKpa3sCO
7qoG2EFaljr5RQLO+Gzo0caH7QhDUrPvMLpRpjDAIDcCjTTGO+dCb/L2z3QG0GtoQcdBpRYFm9LQ
17lq01zyJp13KvvFC2A22xJ5K2rLQT3sNW5vOdX9ss6WmUtHtMYjf4NhRgeSE1aa1gBWMhH0QQYT
ccBpEuLCwMdxHV2jq0ZFglYwxpWXBbl5U3C9+Iw1PoZ/jCvtJpVdIBAjozKKjOZ5t02wACTowFJU
AfpWeWHXBTK28E6n35kl+snlsQWLBrw/HHb5EzZ0anN+I15Y6r2/Up6nYjFgPNCp4jhMbDghK8jZ
Kedb5Za4OVv6aaji//6QwlKbb3T7KVa1ra7YaJTewV/t6w7alVBYNS2qM7ZFwruGctGz0TTHSFnP
u6CmwEgxdyN6bAS5GjhVoB3lG2EBy2adC6YzY04Jtbcbym187oV99xWsz/l+tVP0PUZAkR+D4LdW
984KYNRt6UQGccXeJRtmboieRz40QPRjuZsRmmh6sYwUiJ9J/oD8eCvSnizlv1dkEt56fpX9/RUv
kIU2a5nAmbEOmYS1yu0FjE4jdAlfoMs3w5nwJFh4IleZu/5HP9vbZZlrj3oWQfU31UfhbReGGT+w
f7ADzmtkzzR9l4MGq5Z6UPseiSqRGNPRgiS4yvIuBbP3MlNSU8uQ8cHLF6rUm4Xm+tk4riwlmI62
hQjjE7l7oNGsnqwXQh5CUNdXllcLjf6cFO6ZT/YgcVCKtcRMDxDw9HB1PEz5Mhl94v+FLx74r+O4
O5TITpVlWbizxQ9MS6tsRbYNJInkDPWXDCYf5a7sfW3Pd4KfMGa7Ys1fAkFG78EtQJC5anSqS5M1
eAt9zt+l0o2Bmd576LkL66y5IQkaYvyp8Gg3fcxqafL33+6zglcwvEIYSDD/vMj3y7ywu4/zYByt
C1IXldpLOubaBoOHtyJXbPw4bs1WxVloz9YssZBeryogyf8iqXbQLdq8GtXcnvSwl2XLnVFbY2WJ
vnY8y1ueWHelBYdQ/6o04sbti9hGiCeWS8iTDUqQ3bab7G+9g0WHxGmPY6yiGXgsEx5afo5ilpmr
kXgy7sMnze1yu0bfF5Z8F6WCkLNylmjFFN1Wg2YO6BDCEeGxXj6AfdZJiFcmIpYEm4JCKf8Qai9f
t/vi2f8L+moCwtO9j70IIzlaRLn08PsK5ZgnOhzs0cIXU3dIOKvTsQ70nwAPqtLrZm5MGHQWiip2
LFgchD73317MPnThJ0IqJ4DlB31TyKRrBnFtVKVbithgVO+rs0I/FvfYAcgKhJOkGhF+5tctjZfu
CRsTRZNNhaYHwRNR1TyguxDnKtJy5TPNwTay++6a6jMjUcbveOiivgxDv7nXR+8NyTpma0F8kaYr
zzwSv8d3i+RfFTYqUYtAtvD8zoeFk/5yZB8H3MuMTNitnryemy8BUwrazmndHIrjrJSc2djwHh5T
3xkzYRk9CvFvlTFphnlUFNeZeU/2xgOlheOY/5PeaS4erVtlHCzk/5o5OcK16vfBQFHq5Bla9dZj
04KnenfQ44A1/br7azCH/Qh1fmjgIvvtiCDdMZcihDkQ0p1uv06X9G7Pjko3TygR1jU28gwJfqBz
LVm2oh0b8Oqsoixlt+DpHECrDCxx6ZudIBuoddBsbR+oi45x/e7ACNIPNUiXgap6UysDx1NdssfU
s5jw50ARdQa0SyYXD4KUcqNTGzfpze+BH3Qk6CHvIrZkpl4f5Ujle40FnHTw0OHNz+4Ou4aV6b2S
8HX3BCOyhJDEHgpiZb6IQzITnKUmqPfseIF/CankZra3Asju+FVYEy15K1Uk883hdNVkfNb7R8IT
D56Ns+BNWITXx0I77G/onPjTe/QBuK3knGWX17cN/DA/7dZMxwvZNrZb7mhuh5uFRC+EMdY+y4/b
JiM4jLc80/Qn9dJ1ZOR9FiW25e3+uAQMoFb4RTE6CQ363oeNt5VRisJF0MUcWpZtMiguUwTpdJ9l
Be1mttHC8JubhrLS7rCCFDb4sZntvA3QVw8H3/3P3tFUMtwkLRO5WajC4nB39QcRTch7vUPL/1RX
pA/c5EtOEsmdldcBQezvGzzBgs3xm74jLIOeDfYJxCEZHEXA4D5y3d9JkT6ItY0ObIs5389G8qlH
3OtzG4aMCaJKXgZufyytlIqxz647+Dw0T0iMxcGDS1NUcILxlkd3Ek6LP8LIZUREQvW8gaK4TZ4v
pC+I21U8XaoZubaOpB7Sq0pHH+j7m88BOeDdOMkWOwhl96maAkpzZ4g9kjbqY7YPf5uMO+0BtW4o
wVzuGicSINvG1mEbWejFeVrsf+oWUoJMZyxv5yY/EX7aQjo2Jm7kfuaZFkd1H19Nqe/dEJnKCOvZ
TnIbD6qKav1r9IqII2XiOAIlzmq6CmY5pszCXy72f/E6D2AR0dyxb9YdCuAZ4FHF88hiqiKSA+F3
/uf1fkpISGTLRTpL/4LGu/R6N082KqnB/2vhUKSXahOjWOKkILdZOKjNQBuJk0AqOZ8PuzRRZxH9
CHBTQWhvQZ3NVruI3Tk8zFgJYp/EhVztRupC+6/SZz+bUW3Sc3jbqLv4wWyeogD6oGg0C/GOuAxF
jAXOQB42pqpqvNlXYkK75x1PfgLF+He5PhY2j7SZtMSP4zcA1rJwrejWCcqWKAuXYtRs2n4LsMM2
Yxkg0GP+8XwZ6r6kvcqPm7vc07HCWkTL6/vZjUIrVkB6S78UwOaES9xvruJkmyaWJgbYEx2rAKyt
TiI3eKsWatyxUosLArUuMiEcE8QhnT5l0At2uFqzxs/5IdY+QQfzZ6Pq4MF4pE96aXMgzbkA4YJl
bs+ZlaiYmdTb8+yAJK/1b/KdAi7BJaPZbpWO7WrzE3bNJL5c4/ZLJZ+/dqI5Trixlw1J9xXbsZZG
Vt77hTR0FrV8l8kEEyFYL8PLPTKMAWPF6O3oGlEVX7ZIdLApaNtg2XgDS6va9Ks/VANja1dCi4C6
QvJMzKyGaheWjqeVZWwyuS5x7UU8HwhdUFpZctdruD/gLtNgpjD5CjY46iSZDlqLKw8U7d8Z2wUN
2aQDN0bdLc5T6xNlo124o6FgauC5dDq0gSgycs2jClCZvM3CMwjKZb7hokZYbI5JGZ4YHkPJnAxJ
mtL35aYm0/qlAhAh2tgeE+W3Tiqc7mQ8j0OHhkQKYecdgxZDp55XNP3KTddqxLtKxeu3LYH+uJUW
TugG3EBVlJvtn0pnI+7lLt/ozxOLdzgVBAmoHpHKd3EuZNrLMCcEnn0/ZC8g8A9S0H31Sa6P3AB8
ByUwWSkspcJ7dMpwyA8kExJ5CGgUaV4GhDIG6yEHztbsshgKEQkfKVPMGyCXvRmCE95PqzxLCRpK
cFCqQ7Lb27zAeIlHV1N4o2cqCcDrlypuBlOKogXO8ftJ47HcJeinG57ofkmraV/KSIGi+OJYnNqJ
GiwCYoJGeFi7KdKPUe2/nryHikrftxUFf4M/z5sPmTyrXpuG81sRjWQPNWg+BUPTfSbLyXzGmQa+
fe1pZuqexMANDkfzVnxoLWn1F/120WvwdGq+BwM29J1iD+YN+sCAbHLKyTrlQWKdikPLqUpFuIoC
keFpU3ZtFF2IPsEjNRuqB73S2U8EOGNg5wlln2EDY+EcKIQyK2tKmfNIcNakR+/eFQesvGGzFYNG
irSipjbd166114lHpirY/snbhxpCnXaARsiwFfTFphiUYQxcIjXkmRbcLxUZqa+2soxLh7DENXQw
4b/E9DZqG1HzCd3o+3GffktcDIaHICifACXrmYmTKd1e3TgcaM4kNjCVue5nH7DbPtcYRCicYn1d
w8RjtBOl6Y3hhCBdW6/SDRlaPVJCt3fPqOty7fTjomMTn/hDGmp47+L9OTGN3o2FB5x6Ca+xmwfs
c2q0Qes9tmPPNRQWl+SD6d+sKHhDEj+TCLHoxfXIcd3LYz2cmazhAqlJ8oyGoKxfNp8n3t+kblmR
J0KvKeFaoOGMQP76F75qhZoSyiNUGVSu1gKqXKsMHT2SQ5fljfmyg051dWueMfsTNlHWSFQAnF3o
4f0iIMxuYTl9gIfAiPOA+G+z1rR+5DBu1ssGg6wiyoOzZqhqF6B2700XkIsQj/6YF3CQOJlQcOuk
7VgcojSx5QpSmk8TJd6q+rh40SkapEpwk1P2WZRrLIP3pdDsnVRQApbT2+9kwIA8FXa1vw1VAXfD
7WkC38kCxaai490E8QSFMHdl/NPSSajQZYxD3ibv4t2M+v9KE3ePYOqCzguhTOMyIIEQtzPLh/iZ
vh8ErW39Gd1m8joCvnRk8Jczy2p5DuFq0lcZ2GzWOqgmnku/Cl6KirEwJ+L1Am6GyT8LZmdhffEw
S1RLcUIZuHLKT/2gFslmAytAYqmOMEFqlQV+g5+htce7TyP9Xew/BY5uMqZeX2/EZcz3MCAKhXtB
+Fq0EuJvb1Wg1+Z6LzwCatPhpSTbA4Suj60nVbtzf1VXBJ7wH+Qzn48zYFT6OcEv62wUQHB3bwOV
ajMS/BJOWIFp4aetDw/mVKJK4NLCIpJ7a5NRBPmO0B2WSo/yTXQNEtkSotHLPnkFg0J8fJ0Krxkr
ORifGppJMBvRz5n5x/6W7T0BqjPsmAMZFdPTuVjpvdMEeGxoxa9SwX0ka94JCSngvar7sDC8rDng
+YxBKmM6oxhT8iYGHUObG66LsUVbXipoCCl5ZbMpn8hFt64GexeMha4MIx2GD+/l15H6Y8t6Zzry
dNfGbmFg0xb4WTKHLyaHanpCjly4L+tZtXrLCH7mwAK2Y+X7mzmGJ/yoYMfDN0slLPzUEZXm4kaK
SLnZ/xmcd7kJcb1vHhZfcBW/XRu041+VB0WKrptrdHKZ8EJdF6BYx19KWDAmB7npb12MtNafA2Ml
izWpNXy0SXXXOXs5j9ocFsUhmQBGM8xbNwZGmRGx8kNrfQqv8Ud/fWaYrrKoYJb+IBW88Jc+ivwF
k8ZL/iSkN+/TM5gtBKiz4JUXuthTIVsCvWvJP8zm9H7sdR/qlvJUmsSQZIeEZYPNCgwNayDkxVD3
QU19orgUiiKh6T5ry1yI9FnJU6L2bw1Y647LrCADLYybfsGIIhJY8hy+t+rYL1MJaSWi2YQQb3nJ
Bmpek2A9jMfkGh4kcIyg9so2Xz0Q0eepUQQxZzfYjk3bZH48/U1QKKxfZ73ev1I0KGTFKCJeCKNS
cWw1x7Eoi+GrSPncHqFfDzg2OMjyMv2XQuuQg+yuR0WGfL53wgFqjFWZLBuZMjm+v2TzXjXvTDD4
o34sepP6vPdDkgd3a7G9lnVUKvJLdyu10BvULC5eA/GfmZPQdQaZpndoYRCkDjRHJ4PPBwEYcTYT
5kI9EEB9iUNvc92nZAntGhaD4CUu5534TnZ3LI/F/y0k+wUYTATov4+jY+bmIYNyA6waoLYeMJhP
uB/nhN6p3ueE2AQXkARJymUN9C2u4+cFTBMhcc0dFkiqXWxG8A4GyglK+HmVx1YB88kW830vijmG
9D8qBF04KpoDgjp+dr4CML4l4DPPJpbq+EpqX8v2gZztN8ppIncKhkJasALK+DiXEVs1498hZYXq
fdV+CFckWVed4ptFWhFVJkHtnd8wqvU+y7QZZVQ4DQ5yyQvGfOr2JhpHEgjOaMeBJ9ldPKfXsRKU
byrzhWmiYOtrIk4bGwCTHmCyA3+jgV19Vr2lJLiWfyxnY9pUXsJyJSMX+edI40DRWCBkIbEYmPiv
elMTz9gG5AMA3mm929jdAPnAh5ztqGLALbOc2s+ilCq7MFsvunLBujxOVMfAkpKyMfnRf6dmoo9a
WQ7Z86ML2yI73GOMGREfLjhMdOaiaR8gxCfIFwZRqOQnicGWyPcga6kdoPBlA7fo2VFp/N4tr8xm
FYlOA5Ijeol327Oto7v5b17dwpL4f8ijAYSMCh7cC6tc2c8gH1Zjs2THDKOBIya6fm7ch1CWaBl+
IbQNVcdcrvfzkzQQK3nWsNPyx64wuaKl8EOHyw57DTlpCWWgGT64gzAF3tdw9wcaCgvfj5J95Whs
ZHSlZSbQNWRCioRQQehIweDo4X9j9+atC62AgyZVxbz8QlL4dUzOe42UIyFOopvyLoPdib7AMHaj
rsDC854pYuRvE6/9mw5AcJkvpsB0lTO0ICDhQdW0v1o4x7C7J+6at2e0Pv5C2vh43lYOGbixuZKB
d01kezoB0jfSgqt1XrmIrDVsNQEb/aLeoxF0SJph9yaS9SSkRTFDZdvnNa0o/aqudwjLB9umRX12
EexQ2gfTVQ6xsg++mfQ1pSpCWIgQcZIsCqgnxwGSTV9Nbmxh4FLLs0JUFW/wGXW7cF7nnAwH4cm2
BKZQCYHPZWd/zUBxQW/qxl2ocOdSNjoT++M+98O6Y6zQI0F5uwhxs0rm0p+xVyEecv4lxIYwoFv0
/GR2f/EsD63tZ6uclG823+UMdfGOLGX9THhtzOxxzORjnIm35M44AP9ob3/ZwoUlQsJoSWRNuY1E
E4hpyU5IpTh4Un6yIU2wGFSl8dOjxzqBRjy/U/yHQyQ6ekZmtcb1VyDAyumTS/qjUKV763J4aKG9
vbzvR0B7sDUhNBukZtnofyrqEU1GLQoH7UlwYGHBUQXJQCV/gEfMRKZNyPR1Jx5qhOIrY+bV34Fk
3l+V2PkScN1wk+/LXjcuacsWoBpjkVsQ56YaCjjQrfU6ILw7wppYrXuzSRVr1VuLK0fcxBRYtDVz
Rs0h8cDRa7/z+AA9hw+HGmxWnPi14auxy9WivjjyneIboEtCEjUNVWba4KFfquGeuEPKYmlIWz3n
hUurIdd4L88uf4RmxgNh2VMk9tMyUtBcN3aipCnpJ24okVNKERutvRHrtu35h2DRVC0z2XQjxVB4
P+T/JSHO63yOisbAWA9Or0eV/bZAfEfZmUfDHff7SRdlfn/gRmcpYvNnzdbz3oEdVMOO2lg7ki9o
Ik/SVhmP32+Cn39bivOAQ5becACzNW+m2EVjLBckamV8hPXHyta9pSMl5v9oaRtkSMXgHqbNAKP9
pNUdovrcyqkRzt3S+dE+ASujJ+fv7l00UBoF3DZWteEWrgS7LEY6WBnMGjCfhMvrzKzBbd/CnnjA
5pQvgze5NNbYdvSC6CfZ9n2YrRjpgMMxTH+5Z4fzRJ8GUdAYcCsBSmQaPFrmyYUx+Qo0nrmx4gGO
jep8ccRgFv/UD/3u5l06PPv7r0n2j6hellzSwU3qt7V6Ze1MEJ5NZVAuzxvPJCtTfbV2Dlnp5xGS
OAn4OxKkyYLZAu5EumMM79HFGS3NYBFgzc9aRC+nEZwnyP5E3t9dRf5EROErYxXVmUu9Nv/Bh2PJ
iJSO8Pf0mto9fyIfY511RWYqIWWLqX5213HSZJrTj9WuwwirxFvI4x7/xRGZqfZptc6Swt9a6yTJ
hnkuH3ANGOrliGumEkVJ6Olb1gKoVlGE9TPnzL31PGAVBmBvsxt/2lIfKWU+VCq5CdGuL2DvP5Gm
oj9xLMw02E0oNzS0n17izyjmMt4r/+W9tV+inxqU1yKK20CKwMdsxQmI+0xDWoKjuxPGmnAZoFKP
ZRPiXLtsomYJIMXHYsAYym5m0IEPUlLJtw15EImdgppgvfBC2CwuSfLk8D5U74K+ecx8PeeLjTIn
MZlOL0gDXxPvFTL5HwZVfQoDi6NjzJiLHWRlbNV5ajCqpaZvcGb3lTXElAaoAA8dWlK/x7knnld1
OqCi0l55GIF01N2hUe+A86oHwhx3QKrkqfGFpkm3f5ZPr2YgiUXY1g1gM5viPfdoARSCinKS8qeJ
cv9V0nc739HLMJ1KSTCvFzxmapgcGWlDQQ5HpVA923AJbdHtHMSAyyIU6V+WKC3NXRwXIvyk+IQD
5aiJpGUyTenAPdL+IMFBw432tft8Nte0t0SY14bfNAiJXpE0wXGYeK/SHPVlMUQUwUqXK9tpSZHF
7ypN3ScTHgOvBSBanuhMByqRjWs2myyNC3PoQzK3ZXX0+P/HuspV9pL9JFkKfQUnd7hmekok7yhZ
Enmri3+vgKvdDmYfHmDxRQf67V/I82yHH5jlqU5wfbDYofcLdnFnz6q8i4VBY/K5YA6OONUGephg
uZ8yRTyLpd8lkC6/Ugn3dVrQpcGWbbkm+bPeftqep84FsIh+enMRoQBvlqFCLZgljvvXDObJ2jbj
LkHYih8wTfY7xSMe0jzjAmoRhmCMG/+OZVByHn0lswV9hnh1zeSgdjgf2fvUfm6/n3P5TjRJkNb/
kDJ9pywbwXVC04CWXtBfeopP5uLdF7UNGj2/ZpKXDkZnQAXgYPmndMpEt89mRDxKmpB91rKKl1HF
KphkC9025Lofhi7/JFMyMil+4CU74ubjFy/QvLJBDZVXdLPCgonXMaO6eb0X7aEu5RybRXmKyE0p
A+BmKTuIqBT6iJDx6P9NSNK4TpTIFgkPztMpDmAgT/H650fL+OW1UnROkpy5wWsgFIvsJw23j8MC
qugjTicF+7qVKkGLQOqZ9GUFG3sPat+FxToMrjqyAwB9k8p1+Nw5HouQVr3USKZV7QTjVNeWLidQ
ERlbKYFEOATVU7juqKRkmwE1Nd2HjVvjlFOUmvCSBFQR2CZcAAUREhAMhNqCzEC4nWiUwpQmDV0p
q+PwmzncSZdHgHWAwkwjlxol5wG2o7cwkyMUlR2F5h2TBazHnUFW12TJezijAfRPo5jvzLOoJjMO
tja8RmApWgruIDU2gw3o2pgqVEM4Huq/HchwWubxDZX4XeRxZNEaMJwKgZ3cO1o61SOLHvCpRt9c
G4xa4VrYRUNxqQv43/Zf5hwIPZH5BOMCyFoewVHCeuCeUdzLrEHThY8wpaQHowi9EYkcXhX4VSj5
y9obzI5bbtPObzqShYAVto2lR/wdPplkFgjZru+zykxVu8dGwxuS0znRVx7dcJT4tUHcwhAp1xov
6b0wvr7DkNKZ82KlBGmgv0Jq7bqxNzormLZ1uGUK8NLhBaOLtdUNhBjz8gzdRz9TC6WeBJyZx2Mj
TTkVVlmU0hoKs4Wf3Uffg1nLuxlKHK/R/oert/3bfhEa/8NVsuf9lmHMU/t4F+0lBUjoYjjYjCgt
aoH91PskP9JVvn/FV8s4PfxiIPrn7pQmVzq3jDr1AvodaVaxliywSQwDhfUdW3Z48Tpt3UOg7IHM
z+odESgdMZZpkPsZ6qSGpgn6xhUL0B10q/Mb7v4PfBH+kp0bFJROEgEB29XGcK1faurblB+plcKF
6KttLsQEkZ6kMvlgoCIWY2TtBcHcXNQWJUdCt+5pk+FMw/69uDIVZmYxpu0xdJ7Cxqav+rEmGqtr
cuYNUk+2gathf6VEwBz0jc+p+35kMHR/NYwC/Yn7pUKjIELBDoQ3JpF1a6A4MS+bIalaSXNqXCDf
5TrfUKsT1hSFuKO42vMdIsu9Nye5egwYVAVbQ0q+cnNLEohtxhUslekLwYPPwAhxvVvEicPD0Xb5
643uR20lr6AAKYhxZyg4tcokf8uwZ8cHFcYLrKrKmSn02mjTcE79UgxnYRzBWGEsuAdDR9mHAGUx
vmsy05yb25Jqp09lX5vTKyDyjGAJXt0J24HgKyzipLoZ5JI5bJqZvhmuPrfWWDnnNl7wUGnyH+Va
J3T/7RosqahJytT8KiBMnRyCRd8R6qLdaOmZf5YitkAq0lHRBAlBbn0tPn6sStFS7ogP6lxksG8/
wU/L+Yp54cUh34GwDx9zn0xQDOSZzIus2dd33xhDr+Pk97VCzXkVjHk6gF3hkVP26n63DpcYzc/R
xtoadb9++tZVf/WviN3UZfXf0RgUZ2PUFG9ATse81g46mbL0jlUyWA4giwj0s+LlTplo/VzrBRNv
OUMharYbzIF2OGsfvQPen04f7ZWW/mhPptoNjZ3b0WTh8g2fweXP0IiPAhNjjUekaqbTYeF8eqsi
df1cXAxHRK9iXBFRPTQ8gS6qUFQP3nXwbPxumojGkykyYv88nXS7O7kmPCMi45J95D+jyNqT1ubP
pm0l+S3IKVOVal62gR1/tqjrG+IkQoLXHlHeh3F0qYwrlfroc4vQVUng4WfSjIzs8J0nHxp1IuW3
YQncBKjMD7BH1SiJJGudL7laCAvqbs/cAd+PtVXE6Lt34qQmmLlRCyrsdrvs9VTw4XOlUkVFtDst
2cUPMET6uq/L41kH8qLshVfGLseN15/NPpFRhXWq1k1MHuHy94E6g0RJBwGMLztNCDL3i05ok51K
ngZhND0PzEodv/5oEVN3ZrWArF2Ja7vkab91a3oIzdSr5pA3XqOE/kghZfWs+wybLX6jp3jlQnAJ
BibXXjz7VvEPq5X9GV2owX9cZa8LSNG+CVAKs2zIO1eYe9KBoXJBZtgDe0CByEcIUKO/8Zcg5Q62
DP+ZODOtIz6QWn5e1ykifm+Kq0prv7DNvqKYtygDNGcOyCA41u8bsdfgDLIm73v5BUYfQwKBriJf
Rr/FJA+w5CvbMcsEq5EDDMmeFdEsEAQz0AEUAuG4k/z6kSjlVyd3BgVAoR/8Jh9YkOm8WfX+l2jU
L/zr/RaywzVNFeyXoCdId3/9bnQ77/mBCKKyqygHS8pNDRY+FuD8GiPp70iSil35HOsAsIcXjvRN
+uFYdaBJ98sOC7AipwZi6evB72mlY0G55wji1uiva7gHdBE994ANiRHmmxYxsB6Pq3apPCgC3w4d
xCP1xHchb9HKBRg5Dx5ffOrJ1zEN66VHkDROVxrCJqZURSpJWjxrISI5cxUWiGSwHQvdgX8c4QCZ
noMjnstC8S3H0N0lQOpB+M0DT3IJ3Xd2YLaz8y3Lfcpf1f1C7I3ycgqrbToTknAAp8qYd+/DmOcV
6oO8zvzVldZDgyRHM/INGlwdQs9WRKiWSD9n7qAvgZheOlS4/B3+b99PnPcHYRqiGFnepgSVnOvG
4OTAnRNLAdR6x6CDFEjG0TVXmar5rEBl3bEEEqNFsKepYR7UsYvZsuFiU6HgXdkyxnxV71AuTBEz
11kPkOMAuPWvsH2m4mIpjcomXWcWVzO0vafclV6oXaF/Fe1l5oPnCPhDfda0/qn8DVKqDVvxnnC5
sxjMUasL4E2HhlRquZCBfTtfQAeDQVblKIHiEdNURcb/tEyqx2foPogYslbCcZQ/9A6nzm2eAd4h
B9IMNXfzXxdRVRBeffM0MXPg7PUNLW763ZkXTGFFQj2f94LwGnYMy8bTC+0xy16WR7iCsh2yUTzE
GxqziCvyXd+VON1Psy/nAeGxXAzysnlh52s9sEr7/M/WplKkSgqgdbimybwcSg2eawqH8I7uu8VI
08KEiwSVIr1HnUhd7JvhD1LbDjA0GDtgAo8vUHYzNLcxU9sYIZgLe+Qh9KNttQKY4/kiPscGAzCG
AIBsDQ5jOO4k5buxQSwt41pbd/2T1JAFQaYO+aOLIvcPFUEMVEXa9WKmN2ZqCNkjNXqw2oxBQpWO
Ofn8GagKHzxwphqqm77Z/1cAksvLlIh35mYPA/4pZ1v3a4ULR8Ube/cUj3RBZiKOFtzq4wn2m09f
1Kwo5/PxiE3iLvufyw7lFt1e6d7op70+qXjZEqccoaCm+JK+251jxNwlz5cnzD1np7i6sAVBYNVt
LePYvC2a1MJ93eozEurO5j0PD/Jvrd3qmmuIoevbAwW+FSIwcu+PeXzYtKHGwZosvgjkmVEVGoKo
gI3/zkVWSJDXSjyiFrnLqu0/m1bDY4ftkkz96YVB6VOYnqtNqncXLEHS0XArHR9aU4SggEIRrRJQ
bihHMqQkjyorhXT5movs9HEO+qVQPpwwIWm3irZnOYsdDm1WXzz3Z8uGLANwaquwIQO8HuKERDUY
8oyOM/tDe7vhJJeYq70neqkCQ+zFoBSVoEmRezxEvPlupcNEC4C89vQyrbpgVcRvxhpjNibspea9
uOdH/2BtVbPb1+5u7IWsKIK72bWfYa/MNJxKzcRJwihzhj0YYO75SVIHpcu9OMGOaH4BfzEC0tvG
NavUVdGQTWczzlGlLMTW5jWvg1QiPjCnytI69mPEVEXjAecfSqTn823IfRZdlhcq7MdaAACnMroK
pKh9w7gDhKfBtYIaPQ/Fy27pHniaH6KoUJqCAMlgO6jz2rWa+7D6tFN2DpETQlyEaunjr04V+rEO
99FiWjeYAPMRDcOUvVKC/JO6q5gSb9ubLD722blR3cJNUC8rIXE4bpwwpzV0mtlXDDuPiRJDSDDd
2LEn5t2HjkLq+yol3iD0K/3RjOxQ75sjjR5tBzw8WlKyRR8r1CunZmTuvZ+pM0XnH6CmdnTCWDn+
n7vf7gu0sYjvpti9lYficbRkwKTQhHTO8NaBLcGnvEKozQe0H6wmVZ+EoB8922UD7xLbASynJZ5i
b1tuSx0zgnmOtMut26tfMBRNb/Ul4kKAE/yBeb7ehURjPyGjmU0raxV71zWLAXEViQka2G3wGkbO
5qoybiYNWDP5yhTozBJhzzRMy2xyOSkminj8Pd8ylzx5TSETj3d72MTPO4Vk8jzjRIN/lSdqK1PD
BJOp7qSYeB1UFZG4PzgcDPz+xNap4OV48BjDYHXOhqkqjYa9vo0VuIWYTz+rLoC+WjKNmEaOB1KN
C2LqKYpIS14nTdfHSGGB17UdMj/c95jVAzt7VcUQTufNz7ct8gakODi8nFYp4OR75BLhEF+WcVwp
Bji4iOzSTUC8jtlrL7FYJMRC921Ao5chJTa/pwFfwbUxJOHLpoxUe0Nanh4WYE+9NxATY9IzCYgv
2UMwI/AikNio3pWAyDtgJ7/5nhZfUVWRltWeLA5NnBZF/9FUf0KSf+ZfZp+mPfXVQadpxLvxodMm
xRTjpFI62ss4VpYvfHxh5A08/C8izD1kn4hOtLxCOHLpHCPbjPhxp8eyAlRdYtdXRZNcwIQBPk+8
63AA98GlNnZg8CZIuAFuUOl03kbOh0hr5HBACSI3caS03eOHlrF5oASaPmslSHvJ9GNVEwflvjyM
rdBrXJPl/OMD61gLNhr52D1anTJsbNtLvNTIGgqLV/w/zG4iM28NxvZkXH6UI+grxA3BTQDS7hh1
HKLsXQhNogEmgPtRhQ/78PL7D4HfbtRviroxDZf7tuywcO8vVItHQhxgs7A+C41jOgPBNQWsgUeh
Gq7DK2XTMsvVrqIhmPGYOBDKpxWvXpml5Mvl0P46EKiYhruIt+Nrw9hvZhz86RW23JjWvBbCh6dH
AyuOji4kSqOZXQp/renfIj54c5OfKbNkVQbB8pov45ZAQYwxibcPwFlQuU5cv4CXScpAmY767ala
ZWnGE7i17jVUMRafklozEZ8yqElX+twxR3xEaWOWnM5WmCfpTtt/tdktVokjnM+3zAltswoUbRDP
NpfB5Kdw+8oH6CdBc6GWhipS0EgBpP90iYYamt5vX8ah3mcC+fVzJ4MFYIa17xl+AmoH4A0PxLk9
B8XXmzVmuUhT5YoSpL016YOC+Bs9/WqeksXa8mtFUF+68S+kYvrX7cNizWyKA+K4+fMlgYaOLuJ0
pLPp7Wpwuez5OHlIjLrXgRIbwnt0jwUqXtqe9gMU7Xvf+q/h5tE9y4+8Ro8R1+weDg1eyx2s6xYm
2V2GjOIqFJydNwQ3QknA5A4EJ3eGEXkq5wQ6ddU27RtXrtSIE1xrkJysAAlAFF00XAEw6jzzQBmi
R0dV7J47SFAmRtTdy8sS+1WNcOG5Q2k3j5gJAYokM6sIol3O4N2yUewCRdv0Ojeer1qkTcfUIXtk
8mlXZ0n2+QITuSXWRLHQ+qcGpS0imZy0tmrcG9+4cR+WI/dAe/gvQha1HrHVKSSRae2o18napjse
KZkkGpHG7ZTd7/nGi8LP9R0Ox3v0sH/I0kzcBdoz3E5Sp4Jup3yLEpcP7O8yVSwTqNzAmozSp76h
TzBXcHsne0iFenueV22QOFzLfa24BZT/LAy+kWR8j5QWHiyLgpOhcS5bhQr+b26kVCZJdtkk7A88
dLlEcO9O1lq/yuI76PiJokBhlhDF1pKU3b5jdDkrbTBU9uJVqDSySruf3EhMvi42oY3PKIgKFg6V
7hH9OD8w+q3P1jh3UksF0U5TByJmWEUWfiFa+yuo3Rv0xu+0+YZPcaBdMcqmjcB/3b155swncRcJ
FUW0nrpow8usnAfYmbLHnL73QToQCnsBK5ZH098CjTmGSSHzFU6qgDbPU7AR+75RiSOIUSZl/2yk
zqgkhRzTGJE2Ie0tHizB4OrTLVquXOT2bAuklph0W7VjNu3VjMTheTsKI7Uf04kgc22LLMyE4cBt
jLUYi5XhxHkdyEJFeFIdh2gSOC6t7j8+JwKseWbi/IHQzk8iLOUK19TW+pkD8x8MSbLQ2DgyB630
E/+EVytkz2aSV1zWOivYFXug1zUjMh4LfFCvkietZnBnZtH63E18j/yRTxaBGW0K1jm4wJVXRdKx
yYw6fQBnQSSV5eLBDAjN1LJWGHzl/qZq9hWetbChY3cnDNz8oIbf6ykSbDSF0uVlZLrj33Nh805S
M9jVy0/AZ65eclZpzwqVWJbkiAPNvoCpiCzBWX57wsJ7BaXPkmH1aftMdXqJ7AhsYmAh2fedfDof
Oc9zkg2VVjcRij5mrdmf35s9p1SgqZ4MFLawwEUgR6h5b9+O7tsxJbEF4Yn+48Yu6TEMdx5VhzpG
iV16vT31p/fuH5sOpNqSX3GdAKKQAttzoVII168LXHJu75qGWLg6FxMJRRdRqjnSc/cwcWaILxx9
H3xyehUWeqD3/LCT1vsSqFgT/LeuPoQNsaPP6ug5MITdqhzKE+3UyD6443zyI+4Frc7ud+Wl8f6G
3SaICvy9CVBa2Z444jx5LhGXgGGOIru7SChY8XnUi47enb19eWFKKcik3D14V72fB3Z5S3NQhciH
QjMhwQYw+liQK4A3ieKbTP3F+oqw2y0+SMi1iqw7BprCVKW+SF+BSQMML+KBPLfJOup8cbj0lyS/
MG+R+SQRpdrU+a5HORrjro5l4SeVJXOPEHpZdpoXZKbS0sw9glHc8aUNNbisAZBXY+si6afncqFZ
ox8edijAGO0ENcfITZuaB56CWSJndsUbvU/1wO9Xg8yN2kAhNSZydp2zJqQnMqWN2UsylE5gp8ib
Sdkf0IpuEZ9avLBTdkUq1cXukLGtqBRIznkhGUDJffMOTP3PFs1m2+YH6X6IzIGwKv6jl1GJ4Aeh
HO8/5m+TAlPWwFiFeWXvAfxXrZqaraqDeH3lefJxBXocF0SmF2OsS1LCvWiD+wAoN/LjOcLjBrwm
PjR4E/TjH/zUPMaUdVjunoF2CycrppqJW29ZdmyWtaqHpRe1bh21x5QuqZf2xgVDIVUFEW4UgBc8
lM2knVNVMCGujguA0afxFo7RFF8SUqErH1lvjbgqJpqOW/QHovu7DZR/dKhDrDX5xD6msMdWFxZy
N1YOMIJdDhdFn2XjXc2vaVzzF8Z5u1boCeMbQcI0idxYU5e8LJJurAXAyo0iRXaHXR4iavuC9GqU
61o2E3BS/yhydVpSyXbF//+ZrSBHna/ekOELlylZhBJ/eAssznLhElLDIfD6gpOcUe6vqTW5FxNp
nOg5ag3Ua+ZcnXymLeyRCh/LMRkbh6hH4p6CPJzCZgYCguTwgSx2hHRn21A8LJJfRvdwO6KzPjh9
FVoN8zzki4oI8VXrZEBDAiTUtp8APkUGDB/9qivCUoYnGAR/2C71GhMzEbu/u1rWn+aU7GBa7zeo
aopQHhMqFCkgppk03lLwU6BE77Kgluc9IrWPibaCJRYggawtcCSSnGfO1XJ9drWwPbfuLPtDOQnO
NEU+qalKKgxy0tbpf5nFYJQqxPUsQVGx3YLGZjoEy46oDGzC66ZaU5L82xg9UVZgkgvzi2DxAxAt
zrOQCraGNmvbMF1NCtjLlwBjO4i/Jopws4fqI5YD/8DphqFN/5OksZ2xlNBC6rqwIjfKReahEblj
pGUPgqnZwrikymt9oPp5pWZQzciZbZPGiK6ODBTtMv8nqVBvUbqb5HftB07Ymfvq9VGOelr8accU
jU7ZSjZMQ+/1tbfxHyp9Dw1JgUeJHdEQfPF1M6dSG7l6psJjmAQCxXWKLFQKg+2j8bYXG862wbxm
PCxInLmqgGQUaiUZEBJVh+SCxksaiS9KEYutkOu2xwwj/aw6zpg/eLkeD5zXXXZonEd6iZiv7IKt
LOIxM88uXiaQcbSuEM9Ai+pp4S2hYtLO9sZ1LxUrcSINd/SQqSRq5dmekXNbCYl16igjBpw5UwGi
8QWiAP0ZUfvxpoBWIjWZ07fzQAfdTjEXDvVloj62JJeVz67oIXnRcP8oJqM3+Yl+AD9yH/gkJ5NK
8lHfhStIglMU9Zp32N4fKo5DatpNQkrkT9fQOunTv+aQKlaFxfU9yMwO5wHBPHaRjHV5AJkbOWc6
SvvlDTt2Is6i9z7HgkJReHP4Q4VVWLVtz2CKNVP1fH4piFopI+o6AazFWyI9gefcyrzLmrb9gSSO
qevNil8iQJiuxMbsMgtyO3AtEeNlbjv96j4wndeD+jUCw13GJcNw5eMaR8J+Iww8SQetz3pnNU3J
NuwI0ZUP0t05Zz8n1fEQTm17+RtTHXwd6StrKc5jtlFJ9z8H65iwLXLLMarAsV6+szu5N3W+S5Mv
ZQQTfh8nh/nPCg/7xOLI3DtaCwV/GajUS0C7gH3sGKgXgxuhskyLzJxhrIgDC78l2b5x0ZrIVp8v
0T0d3+GIeN0D3v14SqT2PH8Ic1lwWoUM3+EtoPkMLoanUIXlCW9BYkFP2QQd0h+HMnb1W3u2ySvk
3lEcCZnTx9QOEHLeRUMFuYGv0YxFV6IGKand9Nh7+1oSUfzEMdbSb1CWb2Yb2i+PV1HPg9jdwHHc
B2qKb2njg61EtBTYXDDHsAPD6acAUqcRb95P6IxPOYijTqzKOCLqPAA0AW0DQ9bdI/AI8QCDUecM
r8KpY2Mg5FlwcA274/EzihQ0ro/86R359t31zo6qALO4g/58dfYdUEVtqGOiRHOSDykzbL0u7nAp
gmxeWce4OCTJmHBfOYm97HuI2voIUJDiBiiv4egMNTRbOG1M4t3HSj4UuWNagXnnkqAfEPGSC9m+
SVmKP+6XU4juWXmxnbczG47wnP1jgx5/wVVxoxr/sCycul+JrAjm+scplv1OAQoWvigpackb2nuw
V7VgH1bF1vtZDntW9gKBrGaRt0myO+aW194/WgZKGvm3qiq7e80nDugSy7lqBzFrvkVvgWtGxlkI
LH4dBzsQYX17Abbsg35vje/mp7Uo5cA5MWO+z/JpbkF1/bC+AqoPmWa9muoYUgjbA6v8vLZweXtA
MfN/OMFFAs/2UtEd/ZdqPLnoIg/hKT0PrrGizfBbTGI9HxMQuj6E5SLJ9fU+gluDhXUkO/+9wOU/
VBrokhzJRLlRbShQx8wV9YX8U7otys5A1LPySqwe/b+ABzrs0+i1x1leK1keDMGcy62V5QNDQ4KR
RwvdcgmUM7AKSlrLrrNlMAQHwPiaCR0m8+m/yApnSvqJCdhMUqLA9AhrZOOsCuUHCwZkfN/mq+BF
3UoSDAQPpGjtb3cvHx+Lw9/zg//PQE80TTgsz4w3/1Ipaztu4CQNFtDVa0I1w2AofeIqk62aG1WA
wMsdFrRcVMD474EsYEcudXIU5k/EjrdG9S/TzpSltnVc8OlnB7EXpkQLb7m2nyrD5+CynmkW2nQt
CZJuHr04drghClL5xBxGV/TdOMbGrtmh/6raAmn248el+6GMKTGn9BWJUwWPm/aIGFIMEEHJBTaa
l8FaW+XURRhYb8Ayu6ma6naRthVrzBtUAJRv/SNAXss/eGQXuJEmXwnZCUgw0f6sFWLO7CWjZ4m2
uUY5xJLJrU42SzLfm6iOYlhHRL3IZTfEvwouNTTQ8RLjEgKucSzyW1VNUWJFtqvwSb50GJKUdGxg
3clCatpUarUe8AAiq3k5bhPpITrqGQZ/ix2i0d1GTmlCWPvBc76QtggNdX/QHkXDCKdBqdHX3eaE
qzkA7svqZlNDOVAfNCJys5PDmrB0f/pWDgZqt98GB5X53VjsglxgT0bCn4AwwLBWqE7TsNsoSJY0
K7gxr7Zh6bWj1N/ZG7I9U6ab/zxeqid141AMD9OPhJADaN3W4yYA6Nt+cI1euoMkLvgtcmJVdG0s
yWUPg30++hdUVHJjUPmFxESpQalgKJKvNGi+fvZesGYw0PIhC+FlLI3gVuqzKKWvcUkVpcayi4bU
2j7BGZGVaSNAVGlgXFoHm4joKFM5kHJ0oIPIk6DF06CowKl4jE1Xc9lQxRSr1VfEfGPIO/6Q6X0y
TVTRleoAhbLOaKF4VRiEdsF+2BR+OHWMamNJk+GHW8wlw5xL+v8n01AWmxMv7zp9hjhDJR5sWybA
kp9SkmbIZfZctu6nJcXZnDRP/HJ/yTYgMdLJS4L8aAv9iyt3JuVxAq0ivy6mgeTK5nfNvV6Zayv/
/5r/kSw9VVFiCvFWk2oRb7hkJbk0pT3NK+Am8qJHz1qv5u8Run5iMyPoltZsrxTWRjELWvs/0yYV
UqJ4HQDKgG5V60LTj1ztoqVJEWFePC8tTMx5BlI00ravUzRYaZJYH7nCCPhp+jqfdKE/3QmSZx/e
oYu/whIm70Kz85+ea3Cd81ya6KJwWeF0wDm3Io9zGpvhshJDQKf1metiND/mRn+9iTDQmZiPLOw8
LyWFUyyON01jZBkTAfZbJKGGZl3YDZy02Ie1ZlQzDUUjWgB75Ka40Pv4ZMUFFbnEQHTxH9Fob62H
cAVjroC2wj/hztF+/x3cS8sPTjUjuCNjCTjTnFR+Lw4AoE96YrXLxzjo6jRCXazefaw3afUq3SdJ
58NnvIm6Ec3cBMCF8pORXt1oGMLb05/QUr/7uVpoyLb/DFwL+h//nv5G1aAJrhua97AnVDPO7TWL
K7i8cjTGFzwHutWDrUo8vzkhgkw3nTeAQHj9Wg62mtOYDydpCXAI6eQfYr2zVFULDBNewVOURyGQ
zpzNIvi0SgeIaFNDrZcNQ6WgyZAdy3OIFx69G6f4LPrlqEZoM2nZxVBigT3R6yeKwja+9yX+evfh
cFH3ArHo+15EwDxTc7MssIyMcYJcoukZ7M4FVJBKBhvEesoWPON5rHVNo0ZOgHD3HFb9tKxzjPKV
+eroAlm3p79fLMxFQSbkvzSNe10sYj6O5OZMycTIyYtce7vzjjBPwcjIegu1u8vui2U2sIy9sBUp
DAa13BCAknIUjK2DWGH40qPVyP0zjrCmoseE+KSUfzj136H30d4NNVOoU5tgSnyWqXYdRpOGguZO
KTDvnofSVO0FAlkqGmRpmJ7LEGTckB7bA2hfHyf1gLfeTN2RCb5fBao7J2AoQpa2wT4H7nFvT0Iz
LYw3rMTrRT2M5R009jipES+yL5D3dEkNs7/mbD9s4/xwpqFhFPymVY9x0TmdoDpK+s5a7rvG7ls9
KQStIEn8DqF7RG1n3bZd2hKxOhK3HBKcZwkLNiiiZrznRzk+UwdLVeRyN5Ek0BoPwJfYH3iSOyh1
qyDuOy//yYpgoFQz91nbwhqGeiwwBEf81iIFnNLSRW92xx5BT0z7JKQAf9l58bD+vv6JI82wSGsY
2nxAfeQkOnHRNzRmXfc0TPg6RDLUWmPXKXkO5+X0E9dwtgc0keja/KLBQFUnHBUZ1kUkAE1tJKTb
mV+bfjsCxubaXKv228vu+zxX0tK6vvLQtQgfi6pVK0PNpZgBJrusp1AJEwN6vcRQcrjTKrxhnsuA
ewkhk74s0d/tLSSOA7itWFPgmqjc0ZZnupgp9Qhyjf3ZkeYmOQxhXx54bJ+sMsfFPEcW3JMHzCnH
Xb8ld/dQKZlISt1jI5bbcv0zvdM6jJKLvYyvxbrdvZTMYQelHlnyOxaza+/5u79stCEUtj53T3QA
l/gDIo42EOUnZEATFOf1wdbAb/5gV8qNKY3p4B2KbBGFYXpNEIO3PY3YAg4JvDhWsMDU5po9Yivd
ahahBPoW2Y1zmXwks4bxXiwvqbsHLA34IgU4BXy9pN5WDzVDvJrOpUwbv732W74NE40lxiQKeIGH
jTaxe87wPmGa5XuYLvRqFfMaLFlvk6iPQSfECoI1O7cy9D2Jic8P4YKFjWTaCIkVVF6iBmgNK7+z
yrJFDMmKkt49wzM9SIrBGaaSU/OrZ0B7s7EpST3+fpREwsIwG71HXgLhX/udYcmjduJzTzybdvur
1prbcNzqvDVoZo9vD/BfkQYx5hjSNhJlgOKkqF+CoR10X8Mt+r4IXM/ijDkuBg4zx/D3rqI2WZ8d
XMzt8mwSOSVl5CQsvx1Zusiwl+MJwNPRlK+8w8WZd543Hu3hD0bYAdLCG/BeZewJC5GMbenAhEu/
5mZXlEdV0dw9AQ5NE1GH4H5Z6977vX5lj9QiIj7m4upjHVOPqBXE5ODdyFTo7X98luuKXyjFWMJ4
5Qew/77obouH5/5IPin4p2MaxrWP8OyTyJE4Q2fR7Ht0enfj2eUxvSHFX1hw47L7ORTHPahxYpFz
eJPfjPWY9tYHdZHBxDop9bjgj+WxbBMPetBTstYkZ6oHuQXBG8GhJw5lze7qOIEai2odlYJPUANJ
UCjRBQ7IaqfNxQdt39QwirIz7I3eYx9HtPAfwkPOEuLwnbMQz5wACZvPHWQqdtqxgoVsp0ecy3hI
u9NVBjS7+Scd6C+y7PeUvTrUpCX3+g6dnn9imL6kaB+pi+IJsB+fXqfDptvQx5W5vEKDmT7LIJ7W
Xyj+93MprchNnwU8O7E8a2va/I+zUMmy5zq46by1Kg91cL9+A5UJM8preAeQizVPe1oTeKL3AUxv
SJ2nqwd6x52WQGODgdF3X/f7uCxMK7Pt1Au3SUJc8RPA/9iylGUApkfjxTjbn7tvrHI3xSnkWYG8
jaT6jDhHTA2qPpOjJeDABK+CwTY5VhTu3vSUeD/+CNBrqbivMdJuLcMllD9xgCOitxKR42SQQCYV
2TuSo27/rtihBFIaN2BhmgfIfbjiPVFjLxJMuU27WKoRiRTnGJOGyrqiebRnTbscHHIGbWH9CEPj
LeMv/sJdj00taHCRRqCVCJ6q550qqsNL2W8Tn3JRHGwPJnmfdg18U+IA0yMDNZRJXBk2dSc7VcGV
nMNR2FY3qpX6EsJkCnSeJyhsMtMMnzFOCU4ebfBJ0IqxnlHbpHxCKlpc4/YhOLRIMCkW949kSEXK
mMEJUY/M7h5LLCLrfQh+Z44K1nY9BQJw4b/eXIi4WKJAl2qhcJ8YIm49sCWO256WDnICHYZOHCxc
C0wPrZbmLqSxooLhBW8riImjrmCcgbHRFOhCbPHROFoDnhU8Lp+SGGdgz3oiLOtJlyBamP3HZSQi
yLtN8uSBGJRi4Fjpcs9p4YFgRrsSDxQam8y4LdXXL34z0IO1Ei3scD4YyPMLpJat1el9srDnR1T1
idGIqTvj4LHugrCoDHTWa/mU7iNInLtU5I6X9mzO1s9FUnz9U1UKnf+NlQODOdvIRsLLsEAU/mGx
8EzpkWZKuU3UUnnWPkHetNWF1uXjQjKRKqu1CJJ7SIk3WcqDnO/3GLyc2PGrs1nQ7wqpkdRZ3CSY
0PzZJwFAoLJmmToik8tP3cNGvjnL7024ZS3OobP0qYmbjvnf5PUMZYXolWRR7wXUA3hLJGTEiNL4
Dm/Z5KIk5LxSXrtlgBjzWxsHTBB6m+dvAJxN2aIHD422YkViTminevjrn+faJTu6crgTcUYkxlVv
e6hh7J5meF6fiQD/QWIAzGIYndyehrEqcuELd7B5quCexGnaRUlSgIOJjnUNW0deUfmy2NpWMlaz
qPXoP16Z6Y8XDou4xUs61Ms3qjpI417V9zeYMzhXYL55pQyCOSwC4cF0XBMqYFu9BaL04VrTxNK+
FVG2TYVrZFSIVg5MXX1tQjtuf7nVUyJE+jXoB+O4n9X8fspJ4s9Hz2kpJplxh6ByiiyjNiKIwRy4
LFx94Ybtbs2MENy0HPM7MGcOvgchd3ibkk2pmjmF7b0VkrS7gPXGA9SaPr1IE1zcb4Cb3zFumU+w
ez7paChM7ZjhP4H41viAXDqFCDDI8/4Wc9vNKgUJCIsJ/CdvGgYzU2NPC14VPof8OkASToyw02ni
7u1PxLxGIIcbk7XA03NPRewWol4ghmAtfNpvSgU7UMI12OGaDDZqrOHaLemWqfCt8H/KBh0Io5hA
apjOtaZYCSAM7l0r/wGJJCCdV8PjAKG1ooF1SRzue/Dl1Jl+WXz/8esgkHdGW1duHp3t9rwhW5Fw
46Q+41GB6yqvs91XBKiT71TR82T6hjGYPJ0qBENSgecT42W7W+mRH42vfiRKtSg8P2NEao7Kj6RA
qz+iMnliaX8LgKRm8/++umYrupMpJ3Q5lPfRRZ07OjoLKVaycWILpCfD8Pj0U1R7L+wckW9bqMoN
DlkHH0SwtfttIJ13W21e2CppidYi4U99FwNQvxzNBFzuIotBO2PkO4O1T2k9vU4wDrKbGZEreZFf
NlA0WooWy5++FjEe+jtcKNwAnMaTWJmD8LAYJZwRoKlI5EJ9n4jGlhV2avWAZM79A00imCO78AEX
HBDVYf2hBxwEQQqdPZ8QhU7MNIdZqb9im7puSmvcpEZ7PBA/jC3jyepBULm0BSLQT20ycDYaEg5q
SMj/FVnFL34xTrin7XbBZ3mB9Lv9xbqbABRLGjpml2hhV0apJHG4XXPe/KVijxbuA2uj08xJ3Q/N
xVOLVECoMDCxSeq5pSRIvD8Kr1rFA/tOMmNP1beHrRXvKjURnr0lZAjSIlMRPqnOmQWSC4JhyJcl
hiflPkJ4+nrsL6ja5HHbXDg5A61zO37mxY/+Wws+yl86qGuKOXxF5EUTIz/pFF4rSMOKLUfNh1tS
MEathFIpIkqaMGlet6ktpjgFqW1Nuy1xg1wc+PxZ8zHTnEdr3ETm6ih1gyQPVBF3hdRLym/F/ufF
eWVe81OFTP88N18hdHqh7eXFuH+u4EwxH9VHrEcIMsu7vY0vClSvTk9nh6uXPAJghZwpIpvRVQIA
CDDfBkkpvEf6w1fEUWgASNirHLDWwiOEWx7pUWshDA7hUvMl1QKyQX9Z8YweXO3RK2z4lfzQgpvk
66q1WIHTTALDcpT/3uyAgNOt6Ll77ApM6SMWcRo0YyNmYBbClg8FyJREMo54GmKyDnGphDTYg0hn
byPdZzDcZD8cPyUZI0ovSemdL6OToypitnjyieAw7i/A9Cxt+E08ylCI89TNmwMZjJEGxoBvB9+N
CjvNiLLu4JGgUaxmrGrRVTDdSVLWiDLb7Sc4C5Pt38LRDNb/xa8+GQemYw6fCgatQAL2dfkb2QP6
Zp73iy3XkT1OtTObWYSm6vMsNkHAGNaeu65FXdcD3mVo4djNWuM1MbtEA1YgkP6IgLleQPeGQlEE
VU/r9puat5FV7H5eobwcYCFmJmWlGD55lh9v2vcEk4mM558Nh36/Rv+igvbdbR9JNLG8sPCWG+r5
D1P8dKFuEdQyodOPjuoVXAhMBSEr4n+mlU88C9IHem5yflyVCnR2v+7gc7tpn5hk0QieRNg7oKrV
INaWwgX94WSrlGGAbvOm8o5cWUT6gLtfhRybpveOVhCv/DLielaqxrc2kiMuATiiE2SyKCxfFRbW
9v1aHWamfOPb+VCpLvnXuyN+eGMu20rS2dFeIsjSQIigXHkHD+dhq8H/x0DAtv6HD6CxIfkRC6eU
le69k8nXRbZMNbEGvyzlpTFfonGIkZvAITvQx26AJdX1UyCel2H9ewELNRMPKSETqZM+Z54hZdXh
E2cb5pPrRyXmrccqPppecbzueOihCEc6VfkIdPqGaYbv9eqqZ93/RRhpSQEsNb9nBjpoILwUCbUe
kqvCrsGgFHjJuc69M80B7oh9ArfeOEIpj+PRDlhu5U2SoFfPCV+sXecSwe67MK6iaJo6amobAbGt
HvarZW6VIUJAa9iVQpZgdvP8kefUWfe5ZWEhqTksFBo3I4jGXsaSrc5Arao7v5gZnjddc+SV0iS/
88/o3vMTiXG1bUdp0VjtT0yWKQeULYQczfFEfkCexUSdY7HqX6vqqxVjjC/UnyGSjzwb9GPBkBfE
f3y8y41FYmqc/WuAA+2Isnoj8b3jNBoOl6cluBo66PueqN5BD1+4+JEluYa/pCxb6ly6moZ+mPfN
57eL/0UFYuxDk52JYLMVUSYEUdhmP/DTKJAgLLksYwXSVBZGSTbszPjYrxMDkMM6dGawMMrwdPgj
9ct7b9RJAAQEQOZDWWWt1YhT2Paj5mxn0GoejGLzCya5pzBY9KwQubSsZ0zpyf2aYR6vIoHN8ZzV
fZQs7U51t3H4iixZTjP7lmf+Tk/ymSAzSc+3jp7hv6j9IhcT9IS+AZgOlfKNgMMG+z0kKnOWk4GO
51Hek7JRilkbCEtM2AWrgBaSj2nPTV8tizIPpnoFu4D14P84g47UgAN3z5ZkR21tX0/k/7Ydr2cc
USjFFAo6IBeZan/fAyGxniC95zQSp2Ntl7c+9VMLJi+e8ruVSY+u8JLDx+N5yemMU1Z3FU1s1658
zLe7yfh808lphhRxZq+5VsBfMLRl3S5R0eMUiQSWnKRmHD/h+1WxhsAC3nuC0bXyhf35gXPF9YXL
ylDJzx7JfI7ZNuk2nfrXjrnnzUI0HwFGlI7c9MCVKPjV48O+mzWKu17iACN4GSrm6o19qhwEu/Wd
1PWn3i+DqDSb/CYNNPQO7NqboV6tlLj8YWSVTQiA1jsnb9yn1cOpNy9m0iCx2WfIQeSomNSOBwgo
LZvx7pAYfVToqoSNwexHYCHi6eA7Le2XvEsLe5HMTnd0gXgw9EuzZ8YJaupwp+I2ftZQM5jlD9Uy
IgNoWFAiR4W1yygG5q9xR2FW9U2/ekPjA2pLO2xBbp2W2Jm+dwfCQSaiU/xOgvGsjichTvrDTQUq
FSQxSQDdZbJG6vyqsfPkheAAs/xvbjrD7Leih00FN3NMNFXI9mzsg9Cv+Il9EsM7O02tEd3Amx8o
BjeiyhJevqF+Boa1sYHpbkj1km0Pkm5aDvUoO8fl72d1b0M5+AJcEdZ/oaWQYp6fEEPQGZjrvxOx
6ZlIrQlYXvBKANK1O4fq5ijRS9TSf26agXXo9Aez2Or4GUhXQpFywAhuiq89elE2+NlkZGZAjYg+
rUArrfysSlio3q71DqrqQkD3H+VajsajBRRxiOpyLAmydkMXNI/5Hu/bJ4ptrIkSuyODeOAwg+RM
a0d4ruaaTcFJYMHdyAWnvmW+kiv9hJZWz2frpHRZV1U7Wzd+DLknG1vrY9ecgyW1GBoUiUgF4Et4
qzWrFUFoygLx8N5NADmeTR6MihwLm5ntHvDn2ofhaOAD3ByPlo8NoYWkhgOd9/8vnC4h7FR1OR0/
xIPgCHprYsxJzTp+E+i4lSZDTSQTmyYu/8NiTkVAWVM/stYKQq8KOYEz6PrYc9ikWKQufEHLy6OE
6jZ5pOgwNMLCw1R2hKxcnLBxlLWCufFVhm1X3WTai11tWPEcooOJhFWI9Z+/KS4tEf1+4pzXLe7m
1EzRWDWCTc7aQOw0NCvQA/IMDqqKGOUl6XvIyzDUY22yKI/HCxSgzCN3LWQQ6deMGjY2cSmOrdfD
cIM6d6GzQ9wOpKw2jD/iAtwMu1rJfpYIwRn4SD/CD3RvUYZC7XV52iCYoIM2C8wfwS+gGzf83B6q
o6IvggBtQufs5kE/J+etyr6+eGChCY95WMRXU65Lk5KLKHIbSlkkVEPDqooBFfTK/qmtXETcu3vd
s+lpf7AXzd4YgNWdnMwuvwM/HG92cbm2R8xjEEazz/BtBon7UWlDBNEZGVDqs5DISxYeovtnfGpC
EK2JYRW1cM/1WSNYVyO96/lGOVBNajSBU6Iw/U+5eJi5+ff67MvZj3l2QFEOTanBVlEyQzdWu0Qi
MZ9ujh1lEkuYjBCvHb0tLjTyiclkVzvNXkOCDRlFIyCVDA8YvrGuePh26chqSSHJMOhELLgq5kgk
fWNs+s2v2JWrf0k4eyMISYuZMaNR2QHf5+A1MlWE1tCIirNcij0Dckd+7898sghvEBW4k+iLndFj
Vwk+pjUiMnKtMTgMe7PGrDYroW7Lco3CCOFqiWIAqTm4pXPOlzkLnX31I46JuHMb9Jk6ptykAeWy
Vhh3gh0IfrcuGmZcBfLoyrvePfUW40hTU9M4kaVdeUNrWwVu5ujPPrxDPYLavgOQ2TCLFOQ7hTQ0
f7KArjb0Cq8Y8Rvkf87wMMk32EMgzHpeGvmOJdnKHkoeNVnU9Glc2RcJgtgF8q/8LQM5WAJ5PG6D
VkX3hv5j/7w1XLd7bn4Z/mQkZlRkoIYwF0TGRq1f9YJln/EDfMQH3i944OVLLFQ/8on7Ha5Ooz6i
7E0OwnjFpJsoOXSkJ/77pJkRZhWOpIZarP5qBvh+sdxlqeftfd4VpUB1KDkemr76pPGkoXQazy3h
FIYAPvl4s1nvjV4Mxn2DYYYpOBCxQrJ0XGAqIi02SwDIlpDOq5lhXMq2KQkjKa58cpsMMoy/T9um
0g/sPrdlykBnGJlLFwK1YcQ/n2J2gvtZ6lJ3Gsr8dUstDvJTEhWspImAVKwVs/SjVSqRmxkoPXBF
Nb8CJ+50h3bhCSk0N9H2rxdJo+QzEqwspuhJIpAR219NtHBtIhufg7bD7DOefLc7/hCeXk8EI9+l
rMki11rehtP0yRn4SbuE/Snosks48WYxnVFKjHNPY8Cx+rvcqfC6OwVNMmSueJfdj6/OZNarSwyH
BiGmSFj4oW4kC4lLOgwBpjhoU9oirkeMtkR/NYGt28/VBbVFZhX3Q+OOF/9Qw6lQvJGo2P3GTrl/
OWxZNP4bBRubeD46CgQsUDATe0AvSJWqpQThOHk74aNi9iAZZ7AunJQ/ZRYKTIqqFAezZkT9V+2U
kwsM0Ec0lEO5aPK8RvNZA1zrP88XCMyyg1NWdRTDYMAgAdBekvyhSe2/cHS4D1ButySWDKHLzRUk
KTMpyOfzIug7aW80Vq3oPTVykn0zVo6QAOO4YOk+/UMO0mOmsAcESeRsclfbn7VfFTJiDlxIpr8p
9/L1MrumwVxSsR9OGCVC6HPuMYDd4yvcenSypODakWn0+x06sf6S5qL4flCCU9gL1oPzvioVwXOh
JRrcPUiizdKFoevl3t89X+qre6+EBYTXUg3Fpyx98VPD0Q5sBjY09j72xl36jmRtLtvQ2GRdupl4
vcHsWk1CJStMns5ECU7WiMp2YygB8pZB3hY/hVV5pkXB8U73gJClJ8DEgC8+0W+A2GhedPDWlpbL
FD0BFv2d5l+C4XG6Z2dMlDvKo0qsCKjB8a3zaHpopF1WJ3V0ujske+fTLaQhSaUwVsRIxmoH+iOP
TgGqL0L1ksv1NXtutDqle/b5pq8xsJpm/P8/7vdOFbc9qoqeEZD8RbN4YRIYxSyhBMTqOv3dJjf2
sBOralBN+yw/vp0h7BZU3GKsdiRG15IcodWWRSEThKbf54XTnvv26xpOE13g/MDJAtVsbuapNRcm
Yg47ys67UVvSzTSdBmoNCifB8YUhwt2q8bWPfUf59zv7JEd2JjlH/R3qvzfx9iugf+5+c2jpSvJe
mC2QFdjm/xEm+lyqlLamjCu+hXyc+YccnYp5nl67t2NDkd5ZQ0rMVDnZvLAHchmhZ/tRh5zbc4aL
ImLrgNreiEKljO7cvTXEI968+P2bDqLinRadYkMcxdGWEBSqfxD4mjToCYO1S5rZpLnn861yxmKS
oo8w9qnOQx+vn2X+gnG7VbuCiJ1bMwdIqiJp/rqpmllaXNLAx3j66WDyPUEGJELrFk1NG2aV1EuV
xW0p86TdBxJKW7M3GDV3fghmpxjPD1vWgzs5epwaxH8ueYyAn37ztNji5q9RtN8j/pTQ96G3aQyJ
UQOLsxekX3cCx7/Xf3RukkTiJtQFgqtcv7Ofi3XCn0xvSIUMBq/uVcisiHviS3/jRitS98IMErW1
z6gBufElZVnZqpjg5lc9HG6ZiA6fzytFyBgycmsNnqGLKTx2L4zpeAUNFt0bYtafafX3RZ0YYpOp
iv3zLhDQ2dFNYEF/vdT3p5bL5gMy1hUuNdfCy1t1C1q/E26+QZyiByNxautxO53gyeo+h7k+bhVe
NVYhBuBoOs/GfDGddLBxzRK/jfzXg+wBO+p8mG3QqOmo2X+v991sKkN8Vs+jvMLLqXI7fjt87pOR
03hita4YrgDSchtsrOpMkbuXPDPu0M+vKTbV5DstUwYgmo3XO38qkTYIrZKpqHAZc2LPxeIVS7a0
B7ulb1igyAwK8xv6DxtqDrDfmAEvVBMaKPHZDI5hgt43G40FNLVE55WdYEMAs7PKj0CyB71VCVPb
niFHOkF8kXvkp4yT5BtwWtfIWw5xBSjPRuXqtbmy+Pjdst2VVCNipLEeQ8XEwAfyYqlkMIaETexu
0E3+R5WgqLZBvlba9mlywlc07wTNB1p/x8sjZge6WytOGa8UKn/fO9waSrXaP7Uq7vC9NG0augqy
WsrU6cxK2FcTVGOCjDw1TBUwxZBtDg0VW9taJ/KsWOwOxFd3tHYPuIe6by7AXk7UTE5jam5q6tMN
xJ5x1zqjJdxPyUuRd5+i2/FoS2T88THxknnt3gIi351gotOo05O6I3iClMbP4yZtK42loxRiTVHf
FksfzGBXVD5xdLJlwsigTJKy1+KDR+4LuPJitOq1dS1Cu3WBenxO+8jLKGbY2ICrrm6iAf0oeh7Q
myCSa7ewxagbY96j735FBhjUM3GrIiSnQqEvOixMYoNUktFJMsms1PutoPUIxJFTMyO9Iwz5oBND
dxFaf0tZpg3+kjXTjEBzB0FgsYHq103E1LXlCrFP3zp7hAUjCY22QS1KxUO32CkjhjOR2WvGx76t
DMZkiJj9v+NAsA3F82fTsGOCBm3qu7n8VYr8ryAqQIxJcOsa5hmnTM/gDP+G2nwoPOrFEdXv69/m
rSKA1K5Dsr92hKEDfv2grTN4bA6RiLK5ElyskXAfiSVHb4SXD46mZl0wqWQVPwuOyWhZrybbIWm5
Qcb1SlFBEJsZxA4BnXOG0HBiWnoV+KrUpTzKi47DOWN6xix2BVxWojDzz7QT4LWtpg4Qb7sRqO5R
/NdTjpZG8XS6Q3f0PaZvnTK4OwP/FWz+See+JKakYZvaSVUfnEvziweZLzaB6rY2dEX3WtazU07F
cjVxSd8X6C3m6VMV57WrxMDyftuHf9/nOK0shUYJWSb8pd4rjCOve5w18F+spTV2fIK6D5mTSb7k
x9d5fXPIL6savNS5GZ5oZt5mMo1guOpjkKT9d8L7WFHMkPkD82lX9j70xmP/pF+GpgFu6G4NHN1z
wLzc2Wqy7NKTWxbfmGBVSPy2dl3mkp+ElsSIVZpHDPG5OKBrrTxk58CdWKfiNJxQxaFix3u1Nbbf
FPK9rdWLfBbAiHhNJw6GZRlxcIo6MJs6gFdDuPZR1C6eVD6XQOgz4CDo0AgSRmM5mSBePumdY0PF
mKfO5rSdisVL0hwJm9JMHX0hAwkqzKDUx323HYuyeAu5TUnzwz3I9aqe/E+DeNE/bx5Zx7YK38QD
wDdVgXiZmdwhE0QnF851z9tF/O/NvF6a4ssUYlHAIHIjN6vLDiKjqNuAfafAJLMdgVB2uQ5z340N
qXWhnQzdWR2iop5ujxrMDBPbHicCRjwi35CRZnGKuf3vOueI7Cghlmn5WfjHoJYdiuJ4nWAYmxgY
ZDaiHb3Y/xr4RW7b1oVc0Uvk/wu79SZXPRk0l1KHWhMxJHwRhRLWV55b8ieCPt2e4+vQiegNYrYg
ld+OxPKMO1iLsEhhpts9BG9+YwkDLT2DcsM/S+FbcS7nYZhKmbBChdAd+2I5brGoGATWLgvyb9Wp
IWgPxSgfS8adB27IkDPGh7xYfMnDul97FSJUGFFXw2JdBXjKaGs6MDoTB9S9gqxFpKdNW1gdaskQ
NT2uynUc+Lj1twYth3PMklDa/oxDjjQaIqPj4+wq5FtHmELwrLaf5Ark8J5uFeYjKGhnfpp2cIGO
A6pMkxXZZro06ntjPKk7eK1QxQUimuJ+aUp44A7FQRStDVe2YLPbFqpDWUH+00JhXpJUvynCjIEy
LAXFJMoPpjh9U5a0XetXRDKcvDjYdkwOQYPWAuRPvoEGTgQzgFkC14JsidthG8FNgWhfZ/SFHuuD
atP18Ip9OSyhLL3EEYIAQyvOM37AX/VtrEKSlCpzi69Nj+9qf0WfOzJAXb2hB4SBItPNlu7Iq5Ho
uYsriRKum+1Hpxggnuc4Lvo23TCGtamDHbSqbwFsoJ6KRO+D9JYw8JSjAyTAqHilCBJ4osveIOCj
ufuaKx3m+rYGNetXlkZhJeqNdnW/xhh6tJy44k+G4mbY0baxKPNm1rs8f0w7t0XChzUC2/dIRJI/
/MvR2Jq+QIwFc16ltVP0B96l6q1ItAF+hiKvyxpNDMK5x8y5oK58QVg6L2ft1AgjEjvhkNIeu4kb
MYY+Uhc5di9l5K404D9ZH63T+iDnNfRZjUYw0hijQUcXeTutvTRZUUVYLCk4ffmUNNALWoNLLyTH
3AXatPqaESJMocb12Jqn7HiWULwuHkuS476vFzLPEJlX3qPjZlU19c3uTs+htIpZ79ZdBpp+WmNL
55C9Zt4AyPSeQf3ChkBnugB1ohckbSLhG8BescWpknSn8lREaFczhcT1vPFlzCDApgQBitAGFLnM
VT5ss04R0hWJZZPirj5tQJD5GYD8yfYT7wGCQiUy4OYqYorI0GicPFsZ8s6FjSn4nmveuCth0LKl
Yof5KIyKh4vJnh1sy1XVPxT3fBMvlt/Tzs4dZSkPaJ0Z8qkT2plunUhOfjnqsyqlruubeQ9YEVii
jUvGBq0I642RMjw2t5ZuY2mOFSZpJ+olQnhcL6osDRdfcEPRS4aVTglruSBPThp9EET99TRdRE5K
GVsJgPgrBSmRQFOFfgvGeyJbBFs87IhF7GFUvoA6lfzPcvkMdzmOphbkktCw7b0zHyC9M1qVeDat
uvL1296Ho4E+/FN2ZbMbm3b4XYv+vdZaAOA4Ef8kO/5zniVeMI6rNxTDLjVCTJd7s+ab/4ujH69C
QkGMdeVEFGpUVthLcgBgKt/Fr9LUWaHaWlHpmBV945UiFhQzvsGS9UOwlXGIO6XTrwE21HuUBcOJ
GhSrIURxbutoAybZvAzdP5Wj1wTFZ6cArf/I8bodwBOlm0oztDJgu46g8B7A00McWxdKUIhNMUX9
5qmE6sQRmHaHNewtzz4QWB+ZyMPD+mPrCS5IBV4gQHMJ6yQaf5TsKKIT2UJcy2VDpfHzaU3ufKrb
QKU1B6OUb5aMTwqp3naFWJCDqN8yrIeHiMMzferPvxIJ1JQh0sa78wjNzPVn4Jc3xHVOCp8RgHcJ
g41mHQ+C1HwXqTciMy6EqW/i30SwPMQNUv1mMnuDbTxcg5kgkRJp41yq8vh2qDpfyCj4RuNbTVb2
ze/L8dkV4BX5IijgRWSLQ6bFaJwz/4pgIMaizVJ+GCjShxl0/qN6PMosPRd0hEX8kx1BsEGiDnwF
MBpjNPR/4xNYc/v1RnbBjMLoqNw/uLcaeg4II5zqBRe0+WB0DIwL4WME7XVkvugaVaPUnI22ISgs
R2uJJgIr8EiyUkeeOtC273QlMUz9pgrb7uSpLfOSb0+EDgPZjnmr/LCZx5bjIZjNtKnqoULKerPR
WGLvn0+PM19quWxQeP5yUlKRWxVwhiGCkkWF0KzXF+W/sr2BDbIEKuIMalWoniemu9uauwN9n0KA
/Ggse8XDYdEImfuGSJbglcZke27Kp/5BHMt5E9fDbT62jHAJbyl3vJ1ZtTd9wsLAOLX+6et4sSSh
RuTBDDW6Xy1ynehpNvraONkcqyPQkSt6j7I7ajqc27Pnggw97ZQzSHEVqBdhGd8O6r0u8AJnj2D/
LfYSTVEQskVkOQSZ3IVsAuHfk0ZcONIZ/ejlnLRPdtADEZAccv1T/3O8se9HYSO9OII1nkdxIo98
p9Txl0JZHJ8EoRp9V6nXC6l/eeyDSjYsFkfa2gRhpRcww6gFz7mOe1WmabME+4bfBQYN6+fPkKbL
t1tOEhwIsVqIf9cFQY9M+0b9X/m5JrrACQK/vsoCJ8RwPOPLVbwzRvVXcvD/2E+tsx8FZt7/pqo2
PiLt3f1W9iM26yRDji+vxZIL54UM5HEiZhjybzhX4TTbIs9PS7YTehBctUiwTUk02nelONZ9wje1
Wm0UznBRuPXeYSrBXaxNgUVRzoPfTTVHKMaIVgr28iUjaE6Zk1rFPRij4k+Xla5Wfis5VMuAdxw0
GLbRXh7cVIJGhTyR/pTPMaLNJYaLMEkYxXvmo6rm6ccJ3BcMwR/nQJ1x+PX+u9W5cyPgRqwuKYC+
C+RcyKsz8LJJHs/eoNlLzGI8e/QMeBWmQaZCMPDPphfWezIPTnUbn51SQQQL/paEd6MM8I0UyDQv
x969ZsVOViJg3j51f6k4oSFlv76Ksxhcr8Ji0eG+HUwu/b+/DamqKy3ijDURmRcCDHo/Y6YOv9Xa
JX7TvE27BoJ+HE6r/dkuOLISSMEDwT924tQdf1KvQCeQIHW3xVgZ9BTVbXRQDJjo+EP7jUgJiRDP
3f1w+oV/tpNLKEZs+bb68/6xKVx4rpGQYLmX9GR84GZdQfafu2drYGZJtNQ7cKE6kVLzeZFxqK/p
MFHHgc0blw2pMGSAVhDDrrm5glmaRf9B1489VIL9UFKcq/C88ysoW4EhtPDI+SV0iBO6U2vpKCv3
NNYssoxD0dnh3ypF7Mj2ooLnaW8njRPlb50tROrgO0VvIddiXYhyXrayl/Xcs1kQkDrr9Xc1ln1H
MXkLH/sVTEguEBFq+CgFUSpW0d6CmjH4LhAL8rPoYW3gHNJMy032ei8sNmoQc12PqnreTZ0LFat4
ePRKIys6s4B5CMsmwwfREg+Ef1IvckRmWptADRWCYIeq0trBRjAH6tikWrAewpkGRCFSNezXCdJ6
U70RHyxjrNBDd9+NRsDQNA7vv6xspfUjx5wrKs76bjOtEEmAK1N6NT912Qem48HM/j3gtzWXt/0i
bD7fMaaeacDjXWEFDAHZ/3HDRoeOf+Bd4HmF0n9fO/jMVa3bRt7mZvzkVZ2CqGf+flFKSyhyF3lM
bz3+tnzQmQmUq9DHYHG+Jm7jJvboHp9q0o+LxdLF4mmKmwwMujNrhM2fqruQcIzfytVfwCDgI57l
MdCzUoIH85oS/Up4u5sjCyCY76Oyao7Kh0yOVZm8sTx4KNvUd8mQSCsZ3Ee9j8TeKONBVEwOHucC
phDqiskI5FAgIJ+joqO1HzRU664+avhdbMwAKTTqdnK7IzSAgIbNqfhFz9X1qPQGzjj4Fh2Mp0ep
JVdUYqoqanTTgwjymZ12gMIzepJQQ4mlzFZIAvvzG2vodVJ3UIxv4oYTzQ/SMXowmM4MuT9/C7my
ORPSY3uRaFwaUJ5X/LrvlICbezGZY21XgTALU1e+ZkHRDwKysZ47vftNun555OesaYtclIMteuZm
5ovzDcU7wdnKLwE+OrEvloCbCqSAgjqFNSeOR0TW0DBKRREHICDSDqoIMzM9SfRBCtUhHw/YhbWC
WGwL2Q4lIAnqVJBQceujvY4BpEdccqgVBGsj7SaRsqF+mfTMbKp7pFSW3CuTA7k73nIZGVSjZgtw
eF7uteL6kvZpgtItQTaR+NXm45fueHzynY/MFTakSmDtDpDKunjXvYhqlfIVcjXuJkeAL3FLwAth
pLiN3twrQbiYd3L4x7Cq0F24dPpYIbAQVIZzWAzmSB6pRztt3SDGjCKqmW4WeYvypeAQIj/zUrkh
MtDXsMF4+BS6XbcARihEpwxYUen01drOAanlwUbqw4befhmZdv8NRo6YP1Gdeqc98d0H7Kc7Hi4y
XCsO9EXOvBR4dmDfOOA87x1Tg9rOT/omCJ14pV68BYJR/JukYByqwgGXiT68FM3fTdse7y7Ni/ma
SqO7dfSg9lwH/C70J42EsZPPSkyn0fcI7Ow5AzIvZ3DnCqjkmwHgYBBwqGUrQhWJlE+l36ZTYQ5d
xIjnA9ZaUQZl6iSKRSKgEHpq6/w7oVhJcVfEUJOFhtGjNK0inQzvhEPw8OI6jeYqkSJYMLt9oQdP
ex44IOF9qlNdN3dNsoFCgXIpvx1D+zSjwLqwN4JKlFzqJKkZ0l6zpDmgnzj6l87JQTeRsJ5xK60J
eJEZ0mVLFHcYmnAJx2yJy9YojRc5OINjB0OvzIuZcpp77f/x0InHuNO0O1+aM0CoUZ5jfLwm9W1f
O7Yomoav/wDY/oEGxmLkoAVENrdfyhFFdArDxkxqrtuYE+ugsLL4yBHnObqTNZvjyGcREArKOGIT
Jwmh6s6ohgfVqbL2fXKLmujFjXmuyTmhzSgDrJC/aupmna0J6CsCHwkU59JIJxat70+WZwagW/NA
NbayBrJIIemvwgtsY84RgciGjDeaTp7P4DAJIKfnZH7n8IGx9E1Lk79ZytbIdwJhg9715x7yhwUA
21vGdEnh+NG2h3rOJNb54S0QVXsDFKXcdF4LT3tNDkOJz0iMkuo/yXyyfjd8wZ4f6zcL9skz6PzZ
w9dMGSlbywjFKj+xe5/DYfRUu+8rK/Fh9gj8O8B9oKqgE1uTD+iI3EAaZedspURM3GN0y3QRTI4u
PjqB8YoH3IAPCkkUIIxrpD80iRmIC8wczJlIV3AWdc2jB+Ad4sOTaJm5wzPYA+36OVsBy1dEILWN
2JrGLrKt1c4v45xsOtzfQOB/tsQhsFCBs/zn7ZPRvKIgXwMNAf5OrkXVWRkaClwDAfH8tEYz7nbe
EV6rhZ6F367ZTXmUkOlYUUIYE3xgQ7hAwchsAw4q2oYhPXtSmw220jhBMprjTnZR4e42oCQ1pu3a
BKoajcb+8y6uchgAsqBy39mawuNud8BEYlCybRInaUWHoU47b+mbCr+6ecKUjZgo1wg8mVNMDjUz
CiOnrpWdl31cFuMxt9agzssAJZWR9MrbyPxK2PaCD+wymp6bs2/ncuTVYBVowJlMSLe+0tQI+RaS
8/IyTpM0qzUGqoVvgfht3D2JP0Et1YFymT/rmMLQqMSlBAGVDvPM7XtObssemAO+nEVSK7OYyApQ
m1STNL4BLYuPwsG81fRgOeqjx1BwSPtJpEfix972Do+csf/dN8E6zd24n6Ee3pZ9fsa6CQt6Oder
1bT8/Q2f8xbK+gDIUVhvjXAN62cp2djlktaYCu4nSSS3D+7hY5ftHj2Gx0ui9uzS5kW/ACqgXhCi
OBseJR5+dbsbISZGswmyiC92SqY3c43lm0XX/fhFazIdWJ/gA694nc4eATyxWga0IarjQ3gqTmTw
kydQEPPlro8/mP7bJ66uTfHa2lyHoWQNhaRp/Mhc6ZPpCyJR+Nh4gCKz2qRBuMAFCSATbMfn4ewv
hDNJUw/zY51l4Sp1jIVgLWTJbhPEteSS2rlPEoNNdir5j/X+n9U8wBDuz3/rBFQs9fXO5ocyGTih
kMfFsLn+bKo++1KSpOq5BZsV0lbK0rLNbNwl3jgu7bHLvpXrWAMnMJBDpfSSELNSx7CAFbiYZC88
dA6+RK6MGCl37KSFHcwAh5HoWJRTw5rqry2dQcDcXmOvlGuZx1fSkhJrx3SPIWMXNHw94nZyYFkP
DrNILfFafFoRvKfTlSjh5vpFClH97RW4RJ7q3/YxWixn0frlvP2qLERHM6HlKH+2moJhCBQ20Gau
yrh9dwdQ1GugPLg0S4mngb16PWAad2Sf5/A0yL164JDXRpo1Z/dDgQnN/WACqliGTP0vMAqVI3X5
8UhgaZwPVxC4h5TNCKOjthAOhsW9yeii12ulVOD3ZSBPxjWNFojDlHuMMqpuXa2QfBxUoXONjjPL
cXwVulJtFFC3vZuI/ZvOdjbV1f5Vy3nNwUHBJHTSIrqKz0FJMziG04DGA1zMsm2+siu2v8gDkTsk
lcltA550RBkr2NUrrosYMkg99GA+FLtaymrDXG2wbW05xPjnfLfLKWpitX4bW5OqpX+f8x+DRLbk
872WPzuLXdyhGgVMCod2OL1K0DQJc1aKwWhRiAASv36djaNKtoWkUNoe9MiQLUU9VRK3ydGP4L4S
xA6UaTHJvsNg+w+h6wlyiUJEXx6PeHNug44HxJtidqjxWGsQwek0dJtcHL6kT6b2Cyxfbfrq4gtn
svLUlFkb+0t/B7CwQkUmGHTrNFr9nSYLRLZM74yIhdxhr94oZvpn5sDIzJ2dym2n7K5Pfhj5qdVq
C0gBmYu/5C6x1iLWYRI6sgbZmXIG0mpNwJ/4xSQmPAVXoySo8K3xaNJ7O5motNKiOU/p7h7OL6jY
ZwyxGpbRct9XlZ1ZGl1wX2T8NqeD9hIGmfbn2MdAefBIDji+oP/MKOdKHZqw9mR/G6WdjHjLWcZw
tT+dXvI7sky+CPLgXcDb8MuTyIyG9GtWBEVQp46e2bjrOj15yRjiB3cApVjdOXy+cQPp7FFMAlOP
O/a2iDhtOynbYYflRJM80lBiGM+MB2JKh2hcLAuRndDdkP08jim+Pwv710IkSqbyphN9NhYji6kI
PcRsgHGEB7f+BiVpkXfvrUXJECGGA2EbmprA3p0Y3oJ6H4Ks+msETxGDaIUgm7vgGA0mI6NcfzxD
Xk+Y44hpwkcBrdqGlgeRFMLT1iqrBS9ekPvA8uDRAOS+wYzJ57+DsdTbGvC7YOO8QXRd5ah/8mwx
8Qx0BodheWyvgg3u7XJQ94Xd+a+VUqVglcIUIgbsiqIMFHzSuSRe+/vJsFTxQ1PRN85ABMG2HsE9
MkKfjm7lKeQO+Y9D1CbFCIItawAbKPDGdcXkdccEbG13bVgGSzKmLbyZVStC+eRQNsM+kNG+bQy1
UnP2gCGPKtcAsLxLwOtOqG2uUlwQW1oNcgx+91wDMgg56oiv47Xn6Bb8WBSqUkxqPOJOcdYe5mfZ
jKbOCkY/SrxY/xBwn9bWL0QDyeeW22MNv9Ikq84BVtXoFH94ABOiL+WwjFIuMMeW/txejmO+1fmH
D5RUPfVxHAmVmniYJ0+fYrEu3yVee7LrVWiNVmlouZ+ve66/fUEKQHWRucSfvVlZiCosPk/lInfT
ajmeJ//zpHr9ejfRBDXt5f1ikLIlrgpQqqPYGnJP2x5ysy6hB176kO+RJXREZXOJ6F4FTzAMMvuC
e4I6Gks0sjGWPjOewyF29KjYEOFrNBbRqHSX+go2ucmy9h8g383diVSGgIzismI5yMythfIARHGf
Y/QV7ikm0U4OwsIayb/QqIY3YAyy2BSBy9PCnhHgblV2eaMKR4xM3m6iQh8kI1AIoI5OALUt94J4
5M4Jh3EzA33JYwizo+uZkjZShXcpxp8Yst++kH8Mo5g1w+TT4Hta9EhNi3YeE97NV1yxcH6UYsjj
rlBpcEWJgWswWPyU1kfwiRTjBo7D+VdqguD/5VlevzvzE/n6gyDym/CyMruKWDlWW1Njack4RoxQ
OeyOdJy56oJUcHFQznIBTRhsRBo7Sx6pS+76Pv5PXhGg+AN1kIMJs23pmrJhcKcwpznKOvgXFzFR
04MQnDTcj0CY4z5m/p9Sua6AZSLWUdeuHMg/FBqUDVlJXuBfqnVtAd4oPnBCJgvWgKrlphw0Ap7H
wuC2zALoX0ysRgJXR88SMtxXgTr36SRl8fSo5B5Gs8GWWXD9L5lQjFcq4v//zkgOHiIw+oEfdbm/
xar5QlUxDDWpKyoj2OO0REouz7I3PXckcbsGhZDRn2jcreTvXwLbMbxSrU/W7pOark2TEhl96/dE
EiGLPYeAg7y+BCxUeTZO5jZ1RDZBticA3e+z/6ydm4aj4ckOwqOSCNp1VKlFB9WrqpYJHZSnXXXy
7cBD5EZOV+/QVRAFtdzVF9IFoVMM69cSg7o7FkGxCYaWwKewV/Dt6p3qY0iVRB1s3Pjg9HKL+nCf
gbShkVaMaPYi/JDkAGoLeyYUDbaY+mNPKpfQvKnGPV962J01C3Gk9D3MqtCl0Q3uk9/MCTvrnECK
7hJIwS7goD0P9ubuJdZSxjEyl1kMG9hS4BW6J4XxNzGY/za7G3iQLlHz7v561ijl2q2o/73vKibz
cSgVnv4pHFyy3lIPiZ2CQM5VOyK0sn6u/O6RGnndGHjMj4m/rH5h/qQXGllCcBtyP3evAIwY73JJ
YIUmp3kA2+BVRZaPD+gY6ESUelrnl+M4LtLSDwcRKF4zQOOPhIJMyfKRHnO2OsadUytJp6eVkxAU
VWuvl9g5FJxjCTspA8cfga2XR3/AUSedMVWSnuL19I0GIKAm+aQS8v+ZdeemjAYIKU3mvywTZESv
G5vlQ/wtUB+rL04wzC/aKhmuB9Wy/Ei/dvGzTw+neQCrhyejFez0NU8SMd2kPOUJfYkoXyoD6fW1
KV+DpLihxAldwSDjyKW3hBoLgcpqPbCB41eX+MLl5FlvmllnmNqa/d4+tJdhi8pDNODz3h4ZwBst
A0oXB2Ny7i8Leh+NsJ1suKMSrOc0IUbBsfEyFpEX2wK9IIELbDUTBFRk3qJR9/gXP1KQ6YfNLT/E
hSfJCCgu1Jg4tR2o6/37uatObL940EGjOouxmyJ3MgpciEpvlp/sYWXcarMBrpAIUO7ZS9HbD+AO
+N9zKOiftubBd66unoE59QoUJcyXpFvzYw6cQpn/8EoGOb71Yeu35c+eMUsR0lF8oOkEq8no5ZYT
Ehiy8SX0kwoXUq3f/NdsESlSK5XZeP5EPRb4vI/Ok5HqpujmkOjNEJiXqqYMhPk5GnM8AN7CF5TL
V6iYMKqvDFlTA5l58+xtYm7GqCPKbOVpaH+eygzeyBVe4gP1Xluus4yUgIYZtHKGJUVpXG+NDSli
1oPt+r8leNa/3V1LCo9ZZSH9vNnj5SbAiuh46cJhrH+ub1BDBhCMQsmAH9+NW7WcCiHBRcaUUGYb
lN9qmR5AanwrAHdV3+3amc3nB2KXjgT9hBNDcRVJTh6/g+H2UifeAUJ7KEcagBES/vib5J9HM7ny
jYaEDbWzDXSRt+WeITPRhjM+bMpcv/zQAYAU0gPsM4hohIOnI0gjSmLbbDobiMy1yWwnJaXKw+eV
CqbG8eUrwARzDU4tdQ+uSV5ElU/NidjEN3Zzlp37MQxcEgvCEtCk2ZWfYU205YmZsz+m5y/qqzW8
2WiE/Z/3C2sucvrOQYUFaRzEBrr5L8P0+klx1sKf6feCdG4kcJCTD+W3z/uHR9+M7D5madOeNz1+
ORGhtreFcdWDxGFEhCcMxjrWJ4MFzZRSe9cCq0neuQlssdaW8kkHqnlfbQB8uiEJ/D6HNKM4Cdk4
IEPpi3WzK8/NqgIUqG+C5qNYYIOan5Vr7HdAkf/leRiBr+YiWEpEAbnC+oay/gVb+Zs0aeD49foL
k6B1wB16jezsusTgnuhw/k6gsNkzSHw4QBKobgDZgGKZa/QGPAc0PEBsvE/gfEy4tsiZPQaAqmRk
tXq6uhF1EErzMrOjbJvEtp4Cae+Uzux+1RK2nLdqzNrNiMdyQjKs3FpQdFgINslso0h6ruG8tyoI
KXRoYtiJfADp26S2T5RBGn7SoW/pTab7BcSTgza4VFf35Kb1tEx+pg1saALGt4xcn+1eb6HQNm5+
ZlRAiJdUflh2s62qtvEu9dmTtdKzuTB0cpcp+51KMpOib8JtHfcGjn0RYMhf/lnlX7ewoiHPensS
0G3LKHJBdqM2tU2frEDeLpF4mDo6+7jPzpw5Zwra/aEOFtkRZXBZ25pnvs2hfqpve2Dt1LNGI499
LEK8kKtAFLQdPNBsY9gLvK1CT9PPQQoGKp+sJrPpuzOwUkLBMv5Cop2VuGRNd0mDIPxcVXb9oEAm
yTfK7e9FkZsSlBHx0qZPHbGOeb8/trMLpNP4153XP77LFuEtwbU2/0MRCH+/fj7UcCP7mC+ndyNi
nKgdHQjjPkDH/7Wxix1JOH53jIO+4KxU7Dgt1inkWpHAHMCmFPEmV3zI1fNkJgl7Ut3RK7nClz01
Hgk9fMi5Gipias6jN9jPydKOSC4111ue3pDLRbkiZbAYx6RCtT3lHoWVQQl0aaZKw7G5WiK7FCsu
mQJ0DBLOqms5CBIyA7yO+ba1HeRDZLJQp8oW7L6fc/wqRAZ/wUG1/S2QYaN22I1YHVPkHSjKQuJy
VBLLa/DJ8JB9hCIT0wCm60P9PBhVepYe50L9HO/zclAI13STXzm00ENC/brpLdDzN2Lravb3wsSO
YXlxGR7yWV9N2GGpaPz4Gg15ZLTKoNHucG7e2ESH5jBZmQHPMSteZPSus6WhSt19VZXepLLcAJi6
4COjiAiE6geTdnQo4rQsPwr2iBT/LbFOuGcH+tRQQCyr6FfFcf3AXgHIBQLk5I2mQqNSwjq8XZoL
GqNTkyoRzuIMj3VwtOb2V/XFNCxV4TzlMj9m+4fd9XfKSc8N4PufqyeGqyk8tnNEfx1gZ70RQOi6
d0p11X6ai/VZea3+GKR9GqOPNzyI2lKV5Y2Komj8vTutpEBQl9vtGkGNwUWBmdi76Kuhuh13nTpq
R5NXZZb3chZjZShA2XLAGk2+4R50DBbSOy1Bfpz8tS7w3ZmUdxdKKqBX2xyTJ8uSBmNrwn/dE9u1
a9z9nkQjZjVTg8+4GXnDLRRPLZutpujQnenY+B8cpiKkE10mWEjxdkeuIT+hdQVvTrAgAtaEdp0y
Fv2q4KjrqPM4WgExI1YMg1GOLY0jiWTOEhMx2db8kwlTgNRBxn29P0b2HLgccb/NziWF5mhuwKy6
xSzj61kYUWiINbyrNd0d6x0R/ezAMpyAPgvQMAYLLecW1ThBxb0bowwhAWJHE0YpcoJ0xAvmzKL1
30tlAqQKir5pGhBxIaNDTUp3zFOiI5xwKBxeetrLU813IaBOOpZcNpS9zyizC0geeeqg52dToB3W
aEn7cbbdiUOOQ6A7FdtC+IDW9FaDy5pMNtUfFO+rtzfV4ED0TxKl7wXbBPCI01B/e5IdCzNjCnp6
MVbhbuT/s5Jd+a7Zr8mXGcb81/yGjOq3dAMDRGfLylP0FXzA4CLtGp/+OzBnu7xvLbfbR2eWyOh3
weaG57gc83qBCrLxJJHiQMegDzZc8QTs0jQpsBRee4SWBWX62GLt5qfX7HyNrwJnDhXPqJWYXmeQ
/jEXaKDcTz8EW9gR+xgDnGYAM7XAe8+DmPSVfZTTw6UjVKMuotnb9XLsIz8QmAzGaO8mF/BUB3b2
mEy0ewndvlhzikAYmTrsjb9hGmKKL73sRtNb3AzipDaIDyCUN103J1RCDWLzErdq1Tmt5tbuZdK/
xq61FfFcpbLbZsETGXFlbA1N8NogH/bmysQ4zLU3gcecpv0fTBuOWFZcbinvbXYw3yjNOU4rHgHp
rSx5Q5YajBR6vGjvjNLCiGwpUL9ZXCP11Q2QqcJApIbwqszUafjQ9FLz4nSp4M/s3INLtz/umMoD
mfj8xloFp+h9aGxR5jhq9rhQZGEWqSb+ZE/wtRtW0SmgBOuebuuamhLzHhTifBUKORpZMo75EYKv
2PIPgN9sqrMK3g7Kfz/IKnIUtelAoN2Wx63/HO/L5G2fCNenBbo3Pzp1MZcqEyvLttPToPk6/Adg
lHMmazk5an24L75wUNeh5keYOpq4JoX+0QCJxYUklz/KYyIEYePWEeoZnEAGDTG3156ddm4KnNsn
4v0FOl2XgkJof0W1S9V5ZP0SjQSyHhthGEKa4JianCe0b5/Jqfee5t5tF00x9uEWIWI+zlAlSOev
AKoDtHlvu1dbpBH8K14mfkUk0Rjtna/JAXzxajX3zuARrWafCn1imnRXlf+prgdLq7MT1g9UWEwx
PwwhmlUqW+NMA8zobQaA4rEow5TTGC3zzLiJh0VjZE2ay4nZCFisSQZ7goRSUjgJ5Lc0C5qnROxG
yam6KeXaPmGuBHPcm2X5l1P9fhn/RuoZ/OpAtOe1d/NCGEHaKoXO7+FEQFgheRszOh7YtROWGIGv
w45ZOz8/3GYVKomYy7xLGxGglPQkmIz5xT7JMy0MhALa/Jb/9TFkwiZDo8eYJxjgdy82ITrAWNSg
bYj89+8UmGRCLyX5kYlVeyYpDjlT3sv2fWK8iRUE72JKPbBlcEvi5hdZZnaZjci8n87avgE6Ghcv
2mC/iPL9hocKe6v64pGBPAr/FDs/1c0sGkyy1t0a3VvxFgUEcxu+khWeQogOFJDciyQpQ5WMSEwi
/6cQGOrdU9bpPvAyooHQw00UmedjsUQKKafKKwgn5ooK3KCSMrztYQ01HXOc/KU/qtZfneWCC6I3
6QDWXHS5ePqi/Q9LHC56YCAoWsw83UsYIMwFrwj9ANNCBvQJ2eX1/y+sK22fWBm11wbmzQSSKBD8
b/v7iM+kIkO9IZp62VA+IXcBxIZRAj1rAsqqyVpAvQje0jsK5xuKtlKONDxuV656Wz1H/AyABcTg
ScffuiLfOWxTUxZnrsZXNVdKINPoxOwhIPwm1LnS3N/hsif8KT8rwp5i5vBZJjPEd8eeH9Wqr+Zf
dwdR0z8k4St+qSuBLHY2180vodDLY32svsFcWSqTvxX+GzSJZoz8ZHuDu51NgtTCjcQEjiZkcxZu
m8uU/Qwf87BNlgSm6KROKOLbFso1USpb2H4lXXaILMH40hl3o6xCeLoJlyCjWRm9XC7tpI2PoaC0
QeI4sa17Ykcni9MpFRZpPZfB155ayeSmuqwL72duHS+gDwc51TkQ09WT02u2rNYcZymAdT4daoCB
SMrh3xMVSywPzMYktuaqdTWah4oBguf9RNeTNf/0iL+0X1WjXPk7FR3UuiOd4ESTvvkHXbwGzdTA
9/QCmrYOrqZozKoj4lUzE0mtuieb/b2db7jf5NjRXhXcVuSPEFj9iwaejSFmwFIjGDEzs2E4b9Rs
vVsw2WgGLxuGcWVNgENwVx0KRdyDm9db2SRUJZ2kqBqzG5bbpglfWLiCiEyRGALCsvY8fhUEk9z5
9MqHLI6moUd9SSTfmFxKnIUgyw77+D94M5qi9+LgG1wNvTQ7OQkk/PggPK/oMx/kntGCqQUF0bAG
XOSlcEaMT7NsEpgXoEV7hcbtfUMKLXdnhrsSO0XvcruSChooA6ebAelY+LIHel0po2pQ5er1zDCt
40iVFmD1Exe6QKsPcXb6v0uT5nlhMB9AqWL3Pg8V89i4d9l7Iuh2rg7HuX6jC6VJJkWbutTwW41+
cyfnwi6kdD8fV+lBJp3w0080FhwTF57kTayRS22s1PAx6o/8Hi26gqX41xwAP71EPeu2LtjIRcFC
ramVY0p7hr2p9c0a5T/i+HdInIdVwmjcLYsLVMKJFIOB4RUbS3Vr4dnu9AsUOdb/+d13kvsGMJdp
6T6dC3mWkjK7F/fb5ngTB5DJ+46cBmC52KSm7bbJDDkAZxhbllK0CFNFLJbBHDi30W5hTnkv0jY9
oDqg3/oRNVLNIUze7YosJK5LCzn5lVRn4TlIOQFF62LNWr4jyAFLfu3s3fwlTZZcCMMTRxQ93Lay
CPm5gELd7aoLiYsSZUX99HVlASvisqOlW87ikvm8c4u/ZMP2vgF48crlrh3+qmgHuqWtH5CUJWtu
gIIRezHrOhKJlVFR1kRL5Cmz3r/GX/5zmXm+0X86fWdphur9SoUSeXpXA6NbKImTPSL4t/xVW7Nn
2TE78KPs7MPATmIFf22uwIIdv75n4pikXpj4CMw0H4P1FF7G17K3h8f4shx+37gl6LamltLINeXM
VLEWmCxSbeFgR/nok+DJNVPrbLdzedKcdtVxlRgqbCyAMa4SlRjBbhCqllqWwutkTivZYhhEMkcG
rnQqFbYgT8W9AZ+qFr0JqDVYafVUJ+68lZbRvqx0K0pR8xW4XmdQGwwn1582ceBDIjqokUR4uiSN
BlbeDGzweoLGOgyDvnfP03eljZUlzOb2dDpLCPXzyYvtSw+yfSE+orEg++K4s9779K8XdsavbArd
fhUxpBDLXdNrZM8eYUoP2d/BWsrYJuR0mYliuayPYg22heN8zW8zGa8LVk/OHANXKz1PMXP0VATQ
3j9l6zbPlwEIM5sIXyoFj2r9HJcC1oKkHis99DYlYYyRkrrZeJ2kMCr+dWyFRERsh0mIQB27MiVj
FZU9HhtzKY3ho0Jm1rA2oiZR8ZXv2u8HhMqLWg/X8jC2mkNbDipVhPyWS5ppilyMVbRIBfYD/+B+
kFhFDYDxDQ5hhxwPCtwXbxIOxoYmffTuRCHFswRgeXUszFCjNT4KgRIFoiWaWsikCvxSuBd9cu6e
vWhsMB67t5Fr9Fg6NH8UXuQrRwdpjDp+HUsl3V9hLedAFWzNm8PhRo1P6V0GzyheO5N6crXs69EN
4XYBfk10877A24uU4XVnn/nRPfKE49+vLKdQ1e15hIaaBtZCRCD8n1f0cPOQi6QarVPIf6GVT+zm
SN36xWf3TH+rgpbT/Z8DAgSPWi2xa0rArTTtvtMkdACs5tKEK2hmQEsXPPg4d34v3Jw1N2IHa3zt
yMm2r4vBPeRcfE/1cyGmA29sPejZTh1OD4UgQElhMJlMU8yOkM8XWX+NAJMVAfhwvtDdCPwfNjUn
7UBZ0eFy52oxYzvOWwn2DXzOWoi7BR7y5FrJyFd4560KQJO5rw7t5DpxbHhfL8yw4L2f2hxFwXC+
Us6SrH+u3pqVYZSTyiVcqraMYs8+61B1xB/eGhAjaE1n7DcORaAdiEOjBvZiQtPU7mOcc+rsz001
463gwJZHc7VUwDUrlTfWk9lcL4DAVdNguMVgVAvEeF1IG6ypRNVzlQD1yZvwu09I/swbcMRdUTBv
0tKSJtXtcPCxBNJtKdQzLyir2w0gv9Q0wFlD+UOsAxgxi7jOaviQEa0g0JUHjpFszF24NYHCe1D5
mB7sI0A+ZSi54cA/rJcCJ2T1vwZs8si6kBXT2KmAsJyrnEOUps8K8mDcs39wuODYRjaI+rxTFsaD
BGonMr6qiDbE1KBbEJJXFop0tgN+tXYaqDsD6YcZj1CHMBV9rki+mXc3nZgB7aQFXSSYfGBln7+m
YGSL8pVryNwFh2PwLS1urdjiZ6c0OM8fU7kMeOfRglc3z+hCh2L1N2028NeBQlBbdBgCu0Rx9bah
LvZpFPOnrZ7kvbyt+VFnqGKn6DIlsPCj770zpYu5DS9+BWq8grA7/6Za658X53c6Cf3Hi6Xc8pUP
BKJSf66o1CFDqYow4dbNEFP+jKHl/WokmJVX1Dxw6FpYm+9OneS/jfQLTXAnVo+wU4JJfxIPlG4i
xJ/fB7zZdqeNPEZcMGG/qGwpFxEjzeKLHSkCAUBzGCbt3EtUtT/eyDtxbBG1ndW0aPqORCa6OESi
a71xq0OU/d/C7812cpkCkZYMaeY1D1VNJmrtOJN0rxxNjQ8xmwiMxJPrTgxC0xOcHbUPfaBlrYHw
XjRMVBBb8pwdIHkzbB5IYTdPBNAPQnjvO1T60tJ1Qus4KDwWJKNqZ2fvgqH5G9LEUw3QvYUBzenX
zkdFg7rv0ykSjGF6s0Us5A2fo1wfohyNBhvqYyD9qqayIK/yWTmDg1M46FC23d86+JPWsdMnxOxy
LNNdIkrmb8j0kYdSu4Bpwm/uj9Ck3qpnacxv0wTHEAzIG+NOPgQYDdPNfDEEsPKfGH6h2mHYRxDJ
efVrb3jhkeWrEP+juMKsl5EftSYDrLyDIHpAnUwhh7nLout/xkp7px468xOZiLD5X1shsb7EgVly
q80iRTMTNp1UrSLjOn4SLFXv7i0HlA7JZyHi8j1G8TXjBYX2t1VO7AjN/fgarOmIKSYKipq8/Qqf
MoZKlziulLWAOeC07QjvJrxEBbG8i1k27gvgpCGJzXJyH1EfbxS9wckkSinXL2d4XFTBFfuVXd72
iHipO6o3bIdii5/o4cZPP8NVgpifoVUyxU43g8nzB5kBbUr9Lpw6YO5tk79nUDBECzr8MRrR3Hi2
GCGzgtLsJfbLARIsxPDqV/YS2LJlHj1dIookZ3zeLqzcAPdjG79nnHTSbz0SD/YCf0tvl9H9LCu+
1wvUKwCpBrPZlF6WZ5z+lTAeUZzT1voEnA8NwUDsRtKqQ/LOIU4cagDPNIFNsUxqk2fw5CfXl/os
lnhEfzdOwYmSXdLjBJjy4ttzYCZ2uiuxdddIIb2gjDJdtJbGvRY5rILWuGa9gGSXt9sPm6l1Pi4y
kndDM06r4v+1bf283IU5pcsHpfh+e+QAZctDsBsgi3BORO+8mYiHlJZAoAg6uRMs5mJo6n5IgpzI
xtY9Mn0b1y6AqVM+ukhtgyRSZrumPvFAN/TUECmURkdc3mc4xUYtIlad29awW775W3OfsdLkLWoK
YWgmUSCuHL3UdAlUKTlimN0z383sJkwGVlWWm8gnxHUsXltY3M4VNQeJq3D+mzG2VEOls9HPjSOh
AaZWZ5yi753JoxoT6Rbhy/0Y1eCztjqcxEsU0gw7ivuqxzIym+TpbV6ijrt5o2JYzDZDAarcza+E
bIwcqG8FAQw6BWAMFX4/vXjjUVb2phrUc/vEa8I5df5sJMVlzgLlmQoBsidpyF6tIakeqRrYNdDZ
hGlDaP+wIdtphKZ9Pg+fdX3QATrhWuxJlnRmSESRuUGmaPSmZXASla2pN6C0KaFfAdsa9xPhLQkh
PQ0iL3SY+16vANCR1MSvJI6+Q/++9GVANpxbK9lkrn1jOMlNl2ouxPBBWYWVtcddqRvINbVZXCVb
T0+bfRFdq8YMBW/2Y5xPGRoguVhK6OqpoCYO+FActPUlL2KwLyZM20vvMaPDea60eQB21d9+/pSK
VaYm0EZcsE/RYuwAZDsYlcVpNAj2HYJR+eYSkCbKbeW+/MAwczZ8j55rrvFXvU51OnYL6qhGYtU/
MKRO+YImxp/o3ggM/BXATkTv6tzQKrnyvQybBDlf3fcqv8HHW87jQ+ZGcpsdRwkucTL8Q535i6HI
mxEhoWdUfwQ8PirQcb1Pz7dtYNGokbOnNyz7iy51TlnJ4CEpqw++EkyCLcNGMruv/jUd403fYxc1
USghXZ8KqN183UddQE8te9Ijfu2wPRrqKr6lkeos9na2OqQbXG8yb7NK6JaF2wed2PGPWO52esN7
/gRfzkFIQfOnGoRdrydChG1TWFvt7DJx38y4omaSe5B6jLEozv52Ke0UXc9J4pwZ/Ojxa35K1UWw
1a9MhqiDdhiYNgAw1dI5hi2/au1GxinSwqD/ZHCtWm9XxvtzaDtNgv1+XRvPq9cCAl9J0M83GA0h
oAPYDsRSUUH4KHRd+AwH7ddNrGhrnanO0gnqCnXSmk/XPEJChORhwA4Q7iFtVWWqxn66I533++0x
tvolfETF9aUY8KEluPqKFavgbUbmd9flMPQHatK735yubyQDtGL67fS4+mhqO5aInMfg+KLMR6LV
hRxJI2FiPr6rAbGMzKvh6T3DrYeL6CSgyIWuIxSrCsx7nieq0eR8bYklsx31w0qtsMUeJf+pIoHh
stVD799O/Bx88IU8/NELV3F5vU1/d9+drWmWwbh2YhUqbWFTtg+wGxM6WZvfORjb8dxYkvUAF7fP
ED/NRenqML6UteUiMTJhzYrlKTasHw5OsDplAeZWCC5N4ylR43/p0om4q7aVoKpjSoYgphLUEijH
608EdK1EufDrUfqDXtocr4Gknc4LghTyiNSrQsknV2GrsmS85rFl8jMQOoH+9ef94CEmWh311qVT
cYDXbsFV0O5QYG9Wu2doCmhiJ3o/iUZtnucx8LSi9v0huIAi4MICOzSqw45zX3/U7HQJID+4copK
Efb2lvM8t6S9gng4omKBQoDKqq3YyQf29QDNhY/X/P42sMJl7P0bFzvZ+z1p82XIES69td+hd89U
C0RqkKQNlSC2fxIMLZ5LhKGXXjLDnQPXbVkOWNvucIilfSlpKHwDJeeUpoegZMMP1MFP0PrY0Idc
GVnYwpbDyI+zafpOipo/MUsYubqp2Pzr7/cFNNOY/uNWJunvwwaMvD8tJZHIOAYAJIKP2Y+PmIQi
1q4mdFop+RNJfoLzLM7cQQCq8SRQZpWpj9MwmqqlnWuRErv95SlKfBmf2XYnB6GB+twNA8HpvPDJ
U3V4YoIQF30TpVSk6XadqKga0IVijcm+AkPum7bgCK6xMeHuSCaDrS7aL2gRXGQETnmMsikdDpgc
E9TjFuhPEsszrY2SXAs2IWF20kFFcSgrDnWO7d8yfSYJMJX01P8O4ZcuWDgnwBqxk25ilgxzyki6
VWQPSXfN378b6jY+JpY6smeyINR2oEINvZ2vKo5nPqBaCetzt2tEq9W/7bRIAl8A/bq9u8a3EwaR
MCKea25Z3PkJrU/yJNLKY1gNP9o5Ba0fvWoAw1Qjr8IY3Gxkw9MBKxJwVKTwCzNCGc1ReKwn6/Yd
Xtp0WsghooJnVYy/wQpnpKFsUkpXcxe74xO3ZRZmySFNaniesoEkkfuVKYSS96mlpPp1TzQnhk3c
zacpJlUcxqjwSagcdb/E3MIgyCLBpxXJFZrm0qVLykhKuHr8WL6dMDjuWEaRVWIodhyivSBV2iDh
cSz4cpWEVf/7qGuYt9GBuG5PqOa9BvpYmAdathOZhpFthAtOyds7sUTCBXskR/5dn8IXmjWsea2Q
l/Sw6O24vvSPuAaxtzfvcAXV+UTCbNxXDSekQqsxzbGn2UPErAbdIhlQZtTyY4zzGYufUxiy/A7A
pMW0EPnR8iSrWk9HJccFRcyMfr3tqF0YztbBz/p22Ov37OyIl5kKxPsTUcG9wnIwJK+V8doEUW6r
sgNwyN3AmS7h4NPBJAoa37H15EdYwLb6SMniwbV5DAMhRS8KmVfepHKo7GwHcCwdL6n0YqEKewaB
ak5+sTvoYQkV80DE8rrrXoDFZfxdtBjtcwpU5tGvxvrmJg8yD0kDJ1eJXgmFfo2dhG7UJQESeSws
OiC3u6Atch6GngguEe+y8J5njwoYl6Id097AFZpVZTzY8SHZKWMBLBKTqFoeKbZxVr0To5nvoy47
INhVo5JOAxbAiHzgR3CWAKRA+oUNbG6f6+t13tvetYvj0hujWxIum2zZTbtPPj9lAP/wgG1KIsjQ
Ob0CAxSxnhOKJ6eSmGt4y3WvC+CXpXQmQoMxyZhX4zHulSAxNxLMO9DGagF3T6O8lpd41e78r90R
ASN0mglm+fw7tBRa1Dwq2bEDEVRilxMptm48Y1bNrGiCiqalLZi1EDXOamqJ0Wm0egzj5BpLdDjG
JzGM8TO6NN4hKEIB6HH88Octu47mlCMyoTiN+Uz43pTVtdXZIesP1rOY3wM4f7wbRQgCqc+9bs4/
qENHxdnJ5Hy3WQsBxC4Hl59b3bWCeslXtSXuoYnukHvPzyg52Ousj4emI2V4sm44S7IAW63RW5cr
6LtY10g0hMec0chj5kcKoL8FPm7NQzL0ENoU9DjbbIuMi463mU7fzNqhJEwCA73r/7XiBlLdFmyH
u/ztGLEQMbYPLxVpxPsAFlOS0DnLO6hNix0KWhMfRtcf7UT9Mlo7Ys7k/Y4rx9ur+ZG2RdHnDLqu
lmFWTEmXkmcpbvbUECyIv0bNuKx8qfyaalTPypJ70SQS7q2rGy2j4+5/Xv0+kbdIm8LGs6u0QkL5
p2DLkMYygBE0RKlFOKbatNVEQG1U32HvuLLTApTI+t4rMoiCh0YjxExLkzJTr9PZbqhfdiZm8ASY
HUgxjdTZSCQg8mbHW2oyUZvfdOKPEmbNMfBKWDS75HVrGdOj+DYO9re7SagE7psMK/TJLvXMy6aq
7tPAQm6r/ShUrsqslKYti6qmSHnPAm3c+qTbtJDG4M1mGS6k3T+3jCgwAjVM+n+NWZAKQEdqlGhO
bwv8zo4r+JutEF17im75V44mHdxiYOVNrSZi33fkAk+zzRwuFo/28UqAmg4OioTlW5pYlKZNxPFR
yfg9rqiLPBdu9rNGFT/sbJUAIIm97r62VHhVG4+k3fpmENFtPI/qsBB/htO3QqJ0WbsVFsa5sIqU
6ASoy7D/kTjYzjsvBjdLUu0jbU3JWPy/yzC1R18XdgSf8W8yeVC9zm9L6yvExmL8WEIJEvVXcyen
zwotGJAROLWBCgTHaU6w+YiMjOTwbbIwYtjkah3JbCks9LRTtVkD+plYOIkBOvCvBiFP+6n5amqL
tw5swz95OL8lqfNCXI/CLXJz+sQ4UdzeLw9+bDgto2Pb3QU+VmkXjA6VpyVtQr1MACOv+oHwXh1t
rAgBrWoIfBkCiCk5VJ3NRBrAAHT10scFlJDgXFizLxD1/HQ/Kkz8qSpfDhDjsythoZvxTxu+Ri/D
FFfHAz4z3AY8ppMVX3969rIgdJ/HkqOsijlkAu5hcnyE6Y/aNQB20knYSZyyHATxiGUH8uHacGlB
v72kpChJG2rtG7kV7ERAy/0Pzvvxqt83UU2xF2lHJFr0P8Au9mtRmFfQ5HGpM1BwgxjsFeV76BSU
vjS0g/opeHVAji7T49LkCafd5SOr4jfdNH7zmlt21cKu+pv8ftDBGHSSRfn16YlrWxIoLuwrJE40
MDkgQfqSO6e4RMnKOsV4C2ENJUx/jQ/7nO5ljm0gQ9hqIBZDNvpFpe/aqRZWyZB3AQsusgNV0bgJ
7KJdRTmyaJU+q21VpDYCgorJ+DO9/wv/+yM1B3AbbvKXY31qrFqfF3khF9RTkWzGN6mZG1s9os37
4a56+CszNleI5RZOHCc5A8MXMaOn7dLOJvAT290CuYdM2QR3AvXt19qBt3sl8atJLxCdFwr+E4jH
JHFE7mQvu1/aaYMPgsS2SHYao8gQLpVhyvz6Fy2Tga9FSsulKPt3EDynE3YAmPIgZ5wCaKSgYJsJ
fnuzispIHJHHxdq+kxTAo5vs4HqSxpRaglc67RufRCMntUnVFw3nZy1AEN3bUahSAU+uDRtHH+Gq
xiVgB+rx587YhqfCmQlsugGQumN+6Sv4fUOzGXPo1z+DMy8EoOzG9f3MqjVKudxHIfENcaPIWtgq
RYztj7QvjLX6k92bXwfAMvfjISmm3iXSLH0OMfieozpGQO2RNc2VkIDecTiaE96doe0dIr7C2Gaz
onH1v7fYF3ohqDV5ZMlcr/K57P9DBdf4NApxsOgcVSqXoD4qWWXhBXZu464pgcdO5y72MkvyerhU
NEPzMEoyXdAEDH9RD2vCyGLN4YmpY/9evQnSJ0KMXCfi80w3RxClga4kxC5BABt8I+WzLxz56Lxz
Smrim1D06yiUhgHs8NG4nWXiCxu05HFZqb1u+mqUKv9eETwE6ctXs1xxT9nWqhwNUH2WDbvWTtQG
V8EW2XK5FSvpRscHIqME9Fj4vEM8nA7biVtofGH9VL/qsoaSP61GwJB9IvZSlvkOArAR3vAOHs2p
cxQ4gxf8cZXsSDsyQfCFpkqiT1aBiQ3SZvFu5bkOR97p6XMLVC2rxtg4mzOnMiuskjnyKLxYlo/o
l/6ocr7yyKBv7y2ua2A0Y3PSLOf8zoGTj5Cr7NQs96KAGN7rRTttr6qBkWXdRGGcPC4II0mOMpY9
Ssan0N9k0Xpd98fO/XPC/5/dexFkQH41xhSJ9zIfMcHYnfywYZzM8/ThPoqB+3HT59xvdIQygXgi
lYsDgx9raVdiGRCZPNCG9d+/Kx10sQa/WM/Afi7ILT+l3WStNpIFP67nz5wyY8IqA9Laq+h3o0Lu
e1oFev6MH5CjGETta7W/FtTFTpwgMbptyfAGMrcXfXZUzhvwo0ue+VpIRfRnxczmKqiolKH4dlEB
+KlNzcBzhXqU6IHkMrsizcw2IG1kEHsppCB84+9Fd95EoJd4bcnHqTred3Juw7adIg0YJk8Dm0rf
p2xYS74klLfe/irM47bZ47h+WA36eZEvqrKozfOD+npI1zO72QjH8jBmCmMBCNcUvrn9LlZYXe/Q
+M3VBX5UrIhRPk/3xc7lQWX1QyH7KJYwQykhOk7E53LMDTCVdX7Td1qtW1pr5XwGQutMpjqkH+el
WxcW5KokSzuDp6nbUdJaTgqdU4Ya24nl8ni8FncxmLSDYX4oJ+orqkjKEzq4i/RA5GJp+hQqgvEA
BF3QTFWIYVq9/1aD6XUcKF53jQ+Inl3bhNiMzFqnIHDQCxB/l4Ws7l5Il648lloQ7sIiSd6L4fXE
aDI1srzjQqLRDv52DcdJ7S830gNUuWeQQ3HwswanfJkKkfo9lKpZyUg36rYo94o717mablbJmRXC
TBganIyGmf5QMrFsN/gcZYVpnewaOTIp/QSWvXK8x42lckqa/oaYL+byIH8CbUtelO9EXp7VBrf2
DYIOToug+pZT6RYwX8Ipd/YDV7yifr0Zavive/NGXoFZnflWdjIakfrQwiv6e2s0EQKlUjX9DmVd
kp5O1DjAisltyxrNHF+e26iML3u8hOa0Iu6GhQqF6cmHQ+271n7wTGUayYQt9witW4XDitNYcT5H
oOmwgGQNhiPLjfgOuD7n5KorzzvCE10PltfEHqAEEOmnZmbI2x/wdUz5ZIHTcT3qIW4fqVKNFSBK
MI8T0SpkaT+0kYJ1NToYxzJyDbFtOzpMW0QT40gd3KK+H/Uw7N24t+b6SzxfjNx+Se3X765zz4xr
xV28+vRxvKJK4oZgwGaN1tbI8bzFVYSUkZKMMNLjPkdhiU7M0G/bprUC4y/gCZfVToc1ijqw8UCS
n1Z3zUhGrxu08/6pZN+CO2SjFPnN8preHQgNbVVNzJQ3p8axG1gfDybhr0Di/kzcHBtbcIuHKd3/
bw3uaKfrdxfv+x9b0ezKjqGFQlg0MKiDK2RhjmllcJA4e4pjVGzb5giXhqYilJCoC5b8u9sf7uN8
3iGm8/HpTZTZGAT7cX2qJpavjEUSwxmjT3E0vbWvCUagNRwT6ArtItwFwxcxoT3plIzpe5lb/vtu
C6PxQ6t42oRmZjnffinemk/wtnu8SpYQcwauR8yezfc5e2U1mV2JPkbdKixeJh8b7b34qGAwP+PS
Hc1QEnzNSJPfEQ8nobv+xT5W3TigLD59htgc5NLkIFNs/vi/73zTlyDQcg6BIg4WPM854KVucs3Z
ca1Gr9/kmnzcwVksDtzN43RDP/5YfNz6yo54Ry+V/DnlZfBoBY5C7RQCUqSaIdEbpgTvwgxxbjDW
6lTCzaltcwpm8xdkK9+a2AndUNjd3cXIZVytp0lNR+PC9ldFicQmiztehZj8YaQ8fCs/eiYTAsLH
yi+VpGl5sRHWQXCnTY7F3Sty5vaZ4lFffWE9Ev/kKULabZxjzUNVjbjJ8vEdusvQiLWwuoLodw2r
kQWAuPEuu9NGfQdEzRQyghcklpexgQABgOx2pjLV9hXVoDDirzT/XnrSdBOIwTbYCSi49AmJgLJ/
75ck8quKPgXVjJcfkaDsd/ul02Vg5afFptieTrV8HEQXRfVH4BCqavf5/QJI+EdmVFMvGaXw4NcN
4vRXGZYauaEzi8E4BSOuGP1TdsLIf/YBNtiJpspnEcyJYE1di/FhllFMrnlZ+3FmLObH3/Lxt7Ep
EoySWc8LlZYyZIBKM1blfSf5o4/pKX23735AyfzXN7DQphEsUb/QN/P6sykhjRn6EzK6RjwQ0qzs
LcaE5AA9F6V6mCcxrc0G2APgXfOfqAxCU3iqUs5zz+BPFNJItwKs5yfbyPE/zB4AUmHpqrq3xnC3
x872sv+Zmo4UPxGBeZgN6VCaG2TeM7ulGtrFc2Az4Q7TNbeEgj1JuABdJ85XySLMB0BqmG6h+t4M
krwhFnj9I7DM9kxbaLzi9aAD6MUmT375IUeSoi5c14V+kmiYgMNJStjeMG/iGJWPWz2+ceaw1anj
HhXzOf+0I/qkJocZKxHdMtBXSS+gu9EUGoSREQvCeRRXrWwnKL8omwKimXiq9dujxUctfk6lPghz
YSsJewFqft5Um+In95uHj2m33gS5BdB+S2xmsKqXTIRkaOzKUzEkRcf8ea9MKm4JsIAdqO+y5tIC
sVG2K3G5pA1VYMnpYXNra50WWa4qcHkYjsWn8x/hF9DQgx4GQZXG5CZIgDFPSy0yyev8UusqeN2g
+UIsOF9OxbxF4Rt1RCxfUS4+MnjBcdA6+XwICjc0OYKzkMuLjbi2Ex6cQfZ+4KXfIDeDuO/zeA4b
6/Zq5ugIFNn4PC2a6ojq8Vm0DDFkSc9s8TBd3pPTP7fbnhqsTpRjaNDfBobD6hIqK6pLgDLMCWPo
E+8CqIB33Zc48n50ubJN91fWErcTu919aj3QL6X2TWuihSnUYWFRGN71EvKmhXUOdlG7GqNirqmE
saiXTW3ZhtqY6cpRH/FD7bduNTxUSkPowxd2BaY7ihxYgb4nQ0ySSZiCNuiG/7C9+t+uh3WNHM06
55MzZOJAvUy4y0lHEcKQvRC1/oNC1lgJPMEqHJ0ax+adUapYSCneP+RJR1lVeLAtyVd7i0Pf/Y7n
GmZr1ridRenY0RkRIbqxI2+5UtClH0UN01GlgXXXIPO408Sf68AC0GwtZ3d8otkECr2uFWQQmjMa
r66aypSIkqip4iyKbzrpu5s/GXISzNVmn758zcUuJt83LmK6lLrNdIVkVUOr3YF1t9RSmlHVI+t0
vQbE+a6G/w5QHaJcOvFOPn94InQwSx64dMtAT2tI0oP1bJuiwzEQyULrHHnNlkW5ql7vRshiG3cJ
SnE45WDIDs/E/+XMrkoY1SGoXeO3rd8F/Fn0RfDUUqP12LRKm9LtIRzML61l465qPin7/bTr1t4w
ZlwH2PUCg+wWNtmdMlZhgdhjnAdoxClwbt/GpSL6ECFHmOtR5NdfzPU0f7RE44zODx1EO70IwvkM
Ch9EKSqaNVmyJ4QS74GcblN0Bnggc3ANYIl/HBdo+kwOvV5U4frHXwOrvHQ+SxrksWMvGhs3HHqG
oGbSRnW2AfAqMfju9lYMHapD9WTYSYBr17h6dP3pLNadQzFsOOkfBlfomPUbuyMHWNdaCv05hV1o
/LSInVBkijhd8bpiSRMNYT7Yrf/z5jSdA4jvFt7w4WdMuzWnJZU5OJcC25rFIcnzUnzLFB6hBdUD
C+0XJh2k9cnkJHv8pahR6ZlQeqIPYsdv8Pk7We8frawF1myhJAJUR9LHimPIYZpJhAzHDBjXNOZ+
HckMUy0cxjEn+15vaNMvJvzQq+PFWPtM8oYM+X6LUDVIbq5SY5wSl9GXhov0Jht87Lz8CaCx91M+
aMiToPPGzr2fWip4A//bjx57TRZzy2HiNgN76QjxcVuFmIUS+L/sGzOXyLa6Ap4B+mT+UlPEpMsL
RP6kLqa+gAEAClN8ulXOIAHZxcDeJ71J/12zEMHZ2fFGkos77Ng/y8wp0a77JohGKdljRWqyMHvG
v75uVs8SPpGejXEpseATcLIm0N7hOw+f+IBPr410pPnPGjIVlDA9H0hwtfkCKsh0JTqgyN+rIVXT
59872IDVO7NsjVPYg1S14N7yHRb6hX2qMG8KQL2wmWiG+knWTgn4bXF6zPaYm4yl7XWgIVWkaY3z
HbRi8EXSp3Hx8b/L9Y95CwfgBNWo8r7sGqwKDiFr0eMXadI5Iw6ZkxmRe44ZEzwuHXfrRqr1xk05
EFtFvXX3pI69K+1fwapZ+zSlWWESm0ZN+0lgN1/7eFZmFR6jQe5u/R+GZ47jrB5HXCUhZC8KoR4l
4hkmXLjKdCTSmv3agPsOfTbVL8YeRx2QDgFcsAs/ZavZ6gO35bXH5PGd/WMwZDvL6r067R0bsRs8
vaj/5sPjcUDTe1ExMSmXtu7eCCTchXNM5bf/Gc8PeGZtu4nUywoBADaJWYoCViDmshobpGXjSCHD
uDzzc2kihFq+8E1tWpUpNg8f1SjNIHSDJswjRrZiRo0W0VYzRbl1IRTa1w/0usfMo2jQGrfDiOu3
jwzznQ3Zg1uXPYhYoBYqn9nJzCt480wmJbqKhtbv5lveOEVzbq4v97Rva5dcQEF+IK7LJZB1mNyg
Dn/HZLRO71rjbhz41hvLTBCdXasoXeUoO/NjVaUdUDeNRnMOou4UrTL/JoSjgkrrxaiFsu2AM/cR
dzn72WX2b6KfwktxL2R+FCfgw8zJikP19dB/P9JUMt+npNuWsy3ugM5TF0XbqbgpwimiLSuJfDPh
kQDiIvC2QIDI5q1IkK67oNbjzsfB9FOOAClZGjMADtKlL+IhLmRdlw0K5kckBCaGV5lClrJ7gzLP
Pfi42XRE8uMaSKjjyNYE9qFgG1WY0P52Kr1053tJceN4bmuKAxUTs5rCujGiOuOGqq1K1yIAtpaC
8bCd1NTmKkjx6/h6bWQRvUwFDd2Du3vsMI6EQn+RVy/kIkQ8OgxJQsnPZfDlncnS4s02l0D2h3Th
aYIGJ62WQGkMQ32jQCD9EfAl33pxOlxBYkO4MommKqCHCdVpFz3FQ8/XyGJEpKLvyAyK8fFC6CIf
kct6zILmJjzeenBQxqNiHK6sWrgKKKsUQzB0vR5X4ArFyW8PmmCwsqy6roeHoDsmss0ffBh7PF62
DofHJtzhdkx5VgrvKZ5207d7DFpptD8mFm3TAk4feoUOuLsaiPSRYC1/zX04OxqvSFUsD6JM+4aJ
3ha6i4o+hIGcS/9tzY4xI60Vto6wohxuWNV14n6KVXD05i3If8gpGwoAcAw8dSuqPudpwgLiK6/w
shE+mVCTGSSMYv9glbXOWKN+broI4GIgV/Cf1OuxmhBf4JwXHsAPt0sIrfnBiVufHnhyKBG6HMva
wqjzF/9JPhpsFeNAGcYeFJahextcuMAY16AKWUu9C4cNz4gXOpWBhF8fen4SAd1VyniBrrx3/N1H
4Jzs+0UxV9ZJII2W5XJtAqbX0ALRx7agdBnOxSc03qJzzvjL9r8SUQm5d/ldP+5tKN7Q3rAfHcIw
q/OqkWVkALqtRDJvIpdTe2cibTbEhLLmwov0kJtkXAzXQo4TJco+8kmfPlFCEA2fqf15Lx9WB42p
+ZmMq/k5xmoQ7Vja8JVHRBRVxUrt1F6KXizsLMnHuhmH6CLOqejA3m4pp6BEny0sN3ioqmSYLKvL
eRRObPWy8EpAZCBQXErWhi6YDDuHgqr4FqBxHjl3vn5wQeyd+I6YWIM2DZEoiCCgNlgmhJOxGGOP
oiyVKL0uzyyCKf9BF6x7nS6cScT5/DdZOS9lZRJS6Th6qyyGV8IP9WX78duBw3zqPBQc0fcgJK8R
YLbrGrHbU3VAdmWZ+PD/G7e/f/Wzaf38cgGOfBUjnRNMNpnzGil+TGJTsFXjQZPvNzEDZJjwm4Vy
70RNTSJ25JkWWBrpzRF8yicyOJzRDfXfM0rz5/FNb3sqYpioTmms+WQONx1e7Clul47KuFzmLm6a
fqBw7t1RFTyIpiO/hk8BewUIEXvzuQfnxBs74I+Y0uy5R2ejoNFjVHyU82TtYzfTcq8rUmvE9zVI
Ek3AAMJ5Mm4r86PQ+cguHVhNCFV6KOxQUIpQk073ZOuxIOIOcWvxnB6t8fg7XCeFg3x2kXupPWdb
64PP3xdjfgoLbjoj8b2KaQHb8Hta4BZhHGSkchbv0gT2gQvceWjvp/ohTrF+mpK/JfRM3lLNXBuN
46lt3cvLrC6maDLy4LlbZqE872rxurecRFmU3urodfWEAVRgzNu5Zt3w+r5WygRGWAAFQ6mxDTDs
Satm4ja1jd3nae0g6RcExxhPupzK3edYauvPOw5yGdkTwXO+s7ZUn3MTrb8HhTatKOVdzOicH8/d
sKrKplkSkHYPFj5Fcaz3evEPwV9U1WTM2QPnpA6wxIXlUNActHWGFAooh+r9OinwuRmqEvs54ae1
BHwR7tmQGyM5th0UBR6E8LW6VLZjbL/g8nVG5HpRzk/n6Q3vkZGDGPZpVCe0tG6S1UZB7O7xL2bX
RM3qzsWtHtzOzTw/vb14UC8L4wx8irgKIPYPu5iCoyLXAnlQCWxDi/Hb9T5iPldMACG1G+7k6cs6
kYJzPEVgsD7hxOE58mAC6JFhIA2DWcVTkNzSoTdCreoQq4IoqY7gVJjxksdTEHqxilqVcvAMuiKb
sTH/sHyZwsBCDwAy5WGX1lQC+q6SSrxWKSX41ivknO+5o6clcUYyoJgrQcgGYAIzPfCfdlbMBen8
yzSrCkRYn+ql2u/Gmy7JB/rLbzKcwJ107TdC7z4LwS56jQFDYP85Xi2PhFxnBpAVbbQEL2xRU/Bz
KPxR5CpwpDQYsoCJzZA+IjGa5IEFKxd7CN9dRagketHsylDUDW3eqIyUbZKsgVAw1MQziFg6ui6O
QQO+pBYUWaVP8WaLCZr7aGiG/kQ5xiRhQqSSjOJ2+wLc+Ig2K42I5bC8SUR5pwrBHMIauYnl28DR
/1nGMRSNF8WUjgfUtMkdzGZBUfhBLahtZbPP1Foqk7rXBSTKS1BDEFDFkGL0zD3FpkkuwiWJGl2H
vpBuuHTRRvYu/H3USnhmVEgU6CL8+xg/LZ4/AjYYEAIN+BTiMbvzlxsHCDyGwTdl3UxiT8JWcfzX
aKrpFrSmiP2OxUJYFPeGd3cZFBIznqAyOD8avhrte5lMuPG7Az+ZrGMiR3X1Y34DDqotjHiL4hho
EjrPkTu1n0z82aZMTgz/x5L+SC1cvKc45KuK48lMXm0gTW9sKpy6s7/9KqrPZCihuqfKmZbDOfQ4
STeQsC42OxYLi1lLDVjS34r9eKxVqfUZP1mdgm3Q2zscYd8UAgdox4elk4WU0QSaYD0EGnidEWRw
+DOzBc5XSXxgUkYtgjku3yla9oa9buEQXwSUYUVR0s87aixdDPR44J4453BB3IUrUTF4KYj0Aj01
Q5F+YcjtVEJ1A+jrCYghBf7zWT5ZaWr2U2Nxb6wtfCicMNRT3i+76S+0JZ+04VO6um7V+W0IOH9N
oedTYM0eYcKVm5O11LGePLVMbQSkMBMGEZCINizSLad2mL0pYUKuNzsY4iaRyaSDWErKf1M0+FIX
KKwm0z4OOs0h2djkKYVzrXbb8XbHeu7KCKFYkfIvQF0qIQV/6shoElHYrEQJzhxu4VdJFmHxUOG4
wbA4E6g/rH3oLjrq25g7LmaXpjbUFXc0lu+8b8uu1r5lpgebhMkhwFEf9UqKOfN90jnpBP2jgnft
BRL+I2pXhkU05FIZ6omM32DKbRwZcWAvQUrAiKwpS6kVSqkELM8DZczxzzmoyhAMOvEaYmnyv9Sf
GFa6XKa6CSin6l55A8kUM1hIrV/g5jCaJ4YkYR4o8nP/Vkb7+M5niXEjlQ4jmY2sIHFJjYnp4i8L
HDypo+HffCb/iudoV1bbiMEj2WaTozQ49gNWL4lN1KS+T6azrPUHChsCbNEH9G7/PnG+qPfSLmfl
w/KCUC3wilXVU4iOAqGnp6PYXfew6OUyMeVe5azY69/SXX0ErdfDjhorI2R57dMl/9OdXnFq+Zvq
VDCEbR3EflcuVR1LxCgcGt/1ngqUusZeynafaGRbLYhBIsfXVRzpBaUy/qmBWhenim+hL7Ad1bpY
pziR+kRf1OT4xz42NmN8yBc8+IjEKaeAaCFD48266xdziQwdQKp0faHuphLx9/oJxfDbV4uhgdyc
PUBLmeRKKj0bXgztP0iIepjanVtCIUJZtn6cw0eAEZ242MjMzLqqOby20CKjloydVVX5RePd/cdX
iaFBT8TPTXRnD/RP/dCpZGqMdhm+z4REZp5nhTQE6JLEUthW8dybqP4w5ptgRgnRq5WImtvkcmCO
Rr60WH573C9UiitRvuqQQvPlxiMBNOsz57xhrdWteC5u3ovFn5BDlbTU5Ph0G1GHIEhv23e6eBVZ
UWJ6xkya9j4yL0rKUaWvodk5ZiecFWs+IQS+q2N6BzSXGORNBG1YhDIvJslFh9OUkxCTcubGa3Mv
mAL001qM1CnCq/r5jK9y4b66k8rBznTG4FrVGK0JDBTfltFMyRbMBcFHKjvkXqPJV0DYOfX0tHn9
G2rxsYuoSLtldrKVbh32/sP8/T3VbzrYEoGuO2qCdDaBofB+tK8jE4/52O86EsLjijjL/skcc4HF
8AZ+jRaKsZeSBigUE+tQDWLmznc+zy1JRZd/CNEmqyu/UxMfx2VQt8CWykifEMQOheneeoMIEBFQ
eTRe5N98ItWDHrCkpDqgGnzIy/lLkzE5rQAIUI/RfTAGrunIttTkIhlW9YbVlEXgLMKzmRD1uI5m
jZmgqCn2B8dZ9pHZwWEkXP+hLkO2OV9GgIqNSarELXWVD833Esj/v7MvBiT5O77FJzMlQN5QSDba
HIgTxCY0whejISjIle2f7ZP3lgDjfTtIoYyk4/aqHvY5szhMKdBu65k44tXhxsLCMpDq6WDzZxTw
mzT6LNXg7Ybe95grqvIwxLhT21LanUW+JjZ7NKdKeMPrZZb/bfSB3Nscz9zGsO7c1tU2mPvoN9EI
diyUqMSABuD8LZvBauG/g6Mm8zaxqFrP+Qvea2IuSehF76fAouzGeYnxJbKi3k90KGbhpt2PLNcf
cq67pJE0wr4YpmWq46NAoRp7mNvkEjaP+H6Pyl6awSUosVdmjYA/5cdj3bklfgbciHevmqQC/fwq
3tdTheHLCzvOAAbqg+HWZAN01K3Mzt9bYaKUSPDnZL49ywBkfGWw71gSI+UvaMLCSx8oR80kp8n6
zF28GxzjDC7iFtxBdwoz2kEaOnQbKz8/JWBHE6QeOvs6yfHJpmDyfso8jcz8srBkMlJbOWAieKmq
hhkmL25kJXrupfjKJzs26gQ0c/1A6GlNf5x4vq6qZDr1BbYj98iZ8zADBSY/rbA+MPM0bKfg4FP8
C6LjSXL6Hsse+rIICT0JfRhM6ss/yZKKbVW5JnJVs1dYDxGtaV+UocuoP+2/VN3EFzKkji16Un33
QG+nKnwrDKMYSIwx4RnoBHztQs+N1hrF4nBX9ZGTsukN4m8b/oVF8bbold9NfYSG8dQu+iAcXUoe
MNXJuEhz6Ml/Hqr4E7nnuec50hM0wRJ+fK4WdnZyk9WJH4gIpfclvTEGrlyqFyxXUwm7dbQPRGnH
6c8mIW5GSjVZw+JNDXcnSbZKvXAGGfgI0JmUg1eN0OcHX80rwvzpEOLTZpbKDJETYg1lEsJ9aG4i
gyDKBv7vHPFUyREijsAKtaTY/0Rdl0CP3bzcGZ1wfQ6lAJ5QNaDFWOKU8gq6kJSgVWAxfUPtmUzE
nsYPOGjabC3Yo0mp4SAQ3DqsHc2EK1YI6x+xdocazoNoxToYeHygqqu4LsnRXaSlIaTGlX1W6AFA
SF0sOyFiE4CBJPwgHHszob9jeCFVMKVyE0A/vQgg746agudzth4SB3TMgmZXJHR998g+XO5Uf52c
1VtKk+QKqRLj58R+zm1n2lP+ef8T2mD5BU+T+fh/1+sQLMHg2p74peYj2UiuZSjkO/gEPVGd3qKk
vLTEJAffMAUlEboihmeLT3iLCn7E/wHAADgc5dj4XOGoBFU7VjynsKb++HlX79CodDBcne8pGscu
EzEsJwqMnX5r4DayC1r164AMKRUD1cQHHbBobEvMg0dk64WKhcW0VSbdvJxkFNv8DbZhPERO7b4K
n2VfUN/6/KN8koxn/6vHVay1bmNF++lkCjo/5HjLOlnCi+gdtJRJCMaa/6cycswrqtdI+DieeaPS
qPndnCpE7pVakkuaImvFaIIrtlSQa74BrLh3TRx1qvaf1035aLeKvaxcon31WPznP1DGyT+cdY9Z
fRtOtYQGqMreXyfHyAtzHOPNqJeLeNRrIBljhEwD3sp6gIqK9nzwZK4QClugYXlL8xEpVnwr+xpX
eJ+NQnSQhp65hk3HYYa6pQPmjxERDGVJWf9mtY7fJt81ozCC6zF/QThbG8vEi5/vgKGQJKNoZqiL
QRnWeH7Cej58D609Sip95LKvaa88Jj4UBa/gfBBXbLMmJ2ToITa8+pOa7M/22CI6aF7A8GgLVYPO
NhDp/i8i27MnloasTpRUhghP5LHpoaMQ7I2J9YlR17INu3Z3TtO9zgxdzyixM3lCBzGKb6DN2db+
ebjE1HwvpKVOoibrLj4MyVOqGB3mGVWzaFtu/DBWNwZMyTZHkhfVFI1GCjKpPhGn6hk6/URgGzx3
QXMmChy+JrohLU8dlts3bcQ7GyyXkGd2GaVwZ4JhVCtFXGBM9bCXUqlz09AKaMoM8d+wIE6QR3mM
CS5lFar9MYYKbuWkXU/6XDHVKka+5ZBEhdn4n68aRsGqSyzYuDe5ZIsnsUBH/AxW30vLt8mtWK/J
nnqWjzBz+9nZNBEXuMzgwIEQpctd4vaQjV//6FY8vswJErHBT7RMrxJuB+iFo0Cy0xLzB4QHzzZz
mlnfO3rpVjXcTzbxbaIyoHOk/Z/CD96mHJuR/WviS3Fe1676MaKi2rUs1KdlCAKcb41hZJGo7uS4
COSr6SDsHUd51YoRGG0lr/iitrjh8d4UvvYCEGhZgYqDDeKdY3h3dscVvTWl85/Wqjo8biTyTzAz
MjiY688P7e6dvorE5aLx2V2CDeUNXmpyYXOinPUxClpylw2fxml890AP1dF0d6BgoJM7aTiuXw05
cjq5jpLbYHTUJuj0x3TEruv5KMO/LlJcgK68mngeSWbpBgN59WCJxeDHWOMOtlb8+sgcuaE1Sqg/
G+BqL5s+jMCtzAwuld6PnAPEbq7r5TCT+7xoebE6aZgBrJ81IOy+UfY2lyPeEEWNpDSRVF0nqRRn
a4ETC5GVzgbEB1kNM+whXt3ruNjCFVWiHrpNa051+a+++t4FvrfKQtCJgG8IWxwzh9O8VPD7ZpOX
BOIuT0xzf+mP1A28lzNrhWUESmLaITZIzqFStqHzONvE/VnCuIc+LVJQEYPqrbBn+BhJQom47WWU
hUGpVa2jZJCsvkFuRYrGvgQ47COrXh9MPLQekJ0xgxzznwj6HnTpobMgqjp6eal/aYgKEkMdI8WH
HUcZx2kN8dvVy2LLI8kMvEE9nTdukbyxPBwjwOyX341E361stKpr0UvzLwh+V8WTkPWsbNksxUrR
YobR1phvncB1Sms7kTk9sXzi5Q/vidjZ2OfiCNcGnsv2Y5u4xAcHVzauxOphUd6IJ/tjBXMoiblF
7/Z2sLCrUrbpl0lv3XU2bciOsO7T8YmyUKo0nzsz9pKfCcIPltY3U5erDknZ8YZ1KOMB1bQRXkiX
iF5RPJIktyArPGfFyDBKVaTwdRmUFpwnAiOnYrQ/FCKqXukt7UEWe1wFWzk+pPzGhDGeVf8SUYhB
FbzyjuF9G+Y5MwHAkcef1WO22U9tvKxQLsCIpukvxfMJoxgCyKogYJahNmn73G/Ckj/pxRl26ahy
Ms3TO9VAax1AKy1U9zxBrwQIekpYnviA4sI6y4PEunrC8OW3+vBIMNg16Y6OOIgfEGl+z16IDPzL
mS3gkTi7YT5KvZCQX+9aTTHbCfFqcBQvuSZ7FbUKuUrvm1IH23WUIhaZYzGdCIeeMMa8p3m0OSvH
YNVW4da5NlHAuF69uZCLLERkdD9l5awWvapE83G2QMtupUwovIDKhIXat3jPF8voLG8caWBCvrSr
++50lz9Z2gT3rVpiC4zwHpPPiEtb2UcXBDwG57Kf/25npY0iA0WEGvVUI/FytBcS/LzS9Fd692Go
ayCB4+B/rWLHG0w/GpE7ssfaNFf/GcoihK8QDOg2vu20vR0q8MuhhmmBtZVTt5aNzZvBihxrgOje
gN3kThrJOoz6XiuAsKM8v9DieZ9wE3HyXfD3yKrXohXQMTgmBSBlfeRnjjYXHFsd5SESD5BcwDN4
tjtwsf4zvnMDkjHV21Ngd4yQrkUyR07i+IePj4QRHWyX7AiGzjhVnwhYzDXEkmwUc3qmzhN5/SZb
XT2KS18lcPg1BzO9telAnggHTVix5BLFCLIrdjJoHJLpKTMhYm23is8to/Rhke1wSiWO0QF1aepv
A++TkrnVQJ9+nE7VlJeu0vFwsJmKwz2j+uDcWjOEXEGhkZOQp8k07oRWmy1LKTqBjvmJKZjBTa5l
9ZpcDgsQiUszNfqSgxCoXGoBiWwSYKmyJnHrl1MkmhV8zhyVZSPSeFgAOgHVOy7mA7ug6IZ4oJMn
5Xfz5+Oy+WQVITjUWDOnLMsYzqdUkL/W8KzSGTBF59wFyLjxIdR+mQARJJxlI9+UcWde3n+9myHT
OHsNGJV0k3Eq86zKau2DDHTg//J6pjG5KEno0QZvOy+i17f6VnlwPk8BJxJcSmwl1REB20UfuZIf
StBKWQJISX9P5A/nXQkxXw+RzYQrci+BEzWXWw94NlDVyr3S08d5k1+VSgeacMv94rFhb1h+Y3uH
QKbJssZCPGICU7BrFrWkjmu6gq3jFKtmtt0J7dWWJWmgFjohrdffq7eDSj17ls/BS7f5GDnxAw+G
cSyoAa3yvdhJ24XkuUS4jWfAap8lIPhhQHzO8gn5ErPsFvKGB77f8ZD9k/cBW0vcXQalNfsLlyHm
+eJMMu8RC79D59PhU2UDgQSEDq+CGu6T6BqCyZD3YdhFDNJ/H4nn9yUCKCsFML+JQNUxiLazjsXp
PkMddLf/sE3IhXfhPMm+UOvm2sAsFkmC0bUHvn0RrO07S+PaKSASB+dx+/QhycpEoAKgT/FKfzc6
MVX9j+yXr1HtPTPL1k6FIbAucaefUNZnyeb+X4IQvCaKS7C7lIXagoyigWHp2FJ4b0a3QIQhLHrT
C/pSJRwhbJKO1tUlwBc+agSjTspyGfarw5rGk72K+OTQwxLUewoSQtZt0cO1yfrq/l9FXYqXb/Sg
unycnp+8aSBmnuW4NKjp5eaX5MadhscXSSVEw5eZXTpcSRSVsZ/uV6yWMNDxM03YiY0B0L8YmhYK
aDSq7Ahwhtrbva+7VuKBwi975v+Hc1DBoCgKUR69fn2u6znARFLD1qGQ4vjvVudYtG7xSHla/Dxe
rZfjCIpFvTqsl1AKuW5U3kN1HRCt6UIiGZhFTgDafeqGQvaXnC6lB9zFbCXbCeD4x7iZFTlNDXsi
xU45Nm93JYOGXRvLtUvR72c+ucdR6+6TAxZf4ICpWWqxfZSsQWVQ/LrYubyG32UiVZLO7O+keumw
ZPY3q+ouMOU8ZhtQ5WyTf1wjlx7nVvu/NUKtT8tVDRQ9Ed5aleE00hGuLKjDuxaSsbYx6NtDW0YY
FJzmsjhUy8DwMcGyAsSMYQvnlNf0pBpGlHhs0NCRhsrxmRwcTRBet2KtMkQf6Hx8ZEE/tA9uBrJx
jWNlo+ugSkcmE4Hdh/9jexNxU1tsWlK0o2artuR0vTG30VHNOCziHIAcY7hvID6oWwQZEq5RXJmm
zixCI0rvOSvxnLwQcyqWHpDg9Da17PSki3oTqgaLTw09GGSdDnkIYV50IG9ET1P/jU8lew8t3zHw
eHq3S8ri9PZYBbndC6m1Pj+aEH+EJgYwlQWaMpEh9ah/2rDP5L+lTal7U/eXm1G44HCl31mk6nID
L1DG9RxfG1fDfiE28ACQ28bMulJ9EUbBVEhBDn8Cwyjw8VuXzHXp+/81umIkPdhGtSQlxFaceOUG
DAKmRvqQoy252+YGh0q8gmsvkLGL6NQGKRXTQIeGgX1nuyu6BN2r4jND7f0uBsKvcKybYLg8MPSp
QarLE8gCGnEK+bY/Jb+i3ryGxyZGeTzMScTtcLVFZuhNDQw78YyeeHYnxHgi7JGZZuWG84vVyg61
RjVAizXhtLHjmzLKGGmMUk1NlTF/fjoRGE3lC9U9+Qsu2JBYJ61mY4Nl19zO0xDKEhZb0dFrhSGG
Svwbts6KietlX3Ljsa5hyr3UC8OZgRjiktnyqW5Et/FybSOcH6QCo/B4ycGVAdmtAaHrGf9oDsPa
DrBJMJW6yuVW++Vod/Cl0Fs2+KlZBdTGpgHcgQrA/VeQLNQhf2lYbuocCc0Lv0gMTLA8r/Q6Ee1t
a5ZIAAChURDVk1ItjPZaZ6Rwc2VhiBXb/ST+YjLA2xOG7Yp6Z90YtwQKD0aiPYg+NC8VFQXQMvTv
tqIPypI4Wa2dFcgYlfKg70ypGGD2kvHTu4Qk0uk0PZmC2ZjCGJOemCzMWavrNPx6qDZ8OQ+6Dba3
rOeguN0kfRIUpmDEG66VfGmvZnSRRpwwbIZPgC2GXxZ2hDUGz0hcPff4dH4txJ8lMRtUvmTBM0gx
79K0XMro03iILY4hKkTDsSZoJU6yzpmpiF/MutW0MDKLqKrKO4DnXir9D0hbrynBpbk0wATqqMe9
t9S7Uau7s1lqNorWk+59RCvFfghwkLK1M9sH3RaUztAqavSzm1Rx3W8kwSG7c/5LFNtCMrv/BvuQ
NRi4e5PbUVQMFbZyAcmDZtooncy6CuBg9oHmDv4tHchRkw62MDCgjbI2RNYwnmwmE2Eqp504ZRzz
+3KHiL7XWMf+xFNm+48gXMp9Cr+PL7PHdxLHPT/ypyu+4SdJGQCdijNKV5kZJo0+GtaV1kfZzkqU
Zi6WtTFUbt7IvvmxgB1j2+0VWursLVxj4gvP37J/fdAruBjejt5qPXlzmOS5NKeVxaPzW36V5U/N
NsnwVWct8/t1368/+bGgy52KpKY2Q4T0jnn3AJFjm7SHdSqJ9tKVMUXZbeHpjc9D/nyburLbKOrO
5tFk8ueMa/XSZhxKJOCZDWE4uh6RgRjIhbvPNV6IARop2eJ6UvIyDI9PlGDUo0CBeqcJpc/WH5xF
s+Zdj/gj2rSXueAqW5tIccmP/u7bCYn3onYrfCm2a60wy4M7AftTG7DrDJjmw38u/6jmCgvbKH4V
5pbSV8ahAlHtzAtPCBh4+lCYCPTVQR2CnWP9Gvuwr5M/o0Mr0cVYEo8RnM2r+bQpLbS1OXehdzri
jSsbPFq+vYnCCn2ZT3oKUiAiqTBq7TcldbWltVYbufkCusXLpIV2+kr8s3O0d54yqVq727Bwf6up
Jk5nLOv+a54ZItDL1dZ4fR0xGBeDBkHrQPT9hCfs1tLPqIi04suwHlpAdtadamB1MYU5OdqY/qoM
T/tPNOsW/YA07jtnUMtsVrUzDfwr/gmUEFcpJj3f4n7CUF+SDJpiBKtz4BTi/na0Y/uiQubBcEmw
6rldBydvZDCEptnr1VhFyHozTEqprk7nq4xhllHKbjaKHa8dQi968ZRsv2ewHyawnppSxib1sIB5
/CtdfUtiKWm7eN9MOfBX645s13IEPlStfXkNdCXHk2TkLZ4YRdczq/HRklHfZyc4IzT2ssYFF5AL
quVMhjHQ7zKzDGuKP4pFlLLhxQR/xqLh0o3TLQASNn0/6LvPmgXMyS6d6s3aKSwC776FJ81MxxyV
99+HPeur/cFMI8Y08wWmuJD2PC0vP/wJ6Z82WPgXWFIKSSJWZPxZHVkrTmQcnLyNNEk/H8rnO3Me
zM47I1UjpBXBQfU1Oe41p8NHeBNHaGzg4NfhqSYzdSl9nh6/n8Vr31i9wVBOx5BSYXBRFKRss6v/
4wtZuh6Pfs9PQy+LiuHuLsWO5bzkzbBUsKfeamu+Nb8gD2V/TZh5EVUvbDO0KMsZFYp4V2P5Ej69
1yKRwpGMHaBVwKuzEgpsmMFSvYMzeJK1xGTFpN7VVjErWdU3G5YW8pXjBpTuNC3Dtl75OUskvVJB
j7CWUQvWMTo7EZxPPkY59Wd+rFi/dSwBa4U5P7ZjmUGApkVvkbw4MD+8SHgMZU37yEKvbwX9wf/Y
oXIMX95grTg9JDNXQpsnhEUj/eJd19ip6bavcFDmIeaYA8slbhFMKdZCnZNnxBWiEecvTTmNV16M
NSl25jPRK+XrTe08c+DMKRO/9DjFHDskI64uQtdnjoL5eYa5Ei5xqUUB/pd+P4h8azZ4uoGwbOgW
b41c6Tow1bEr+8qwy5PgPdg9FUym9cfseO9r13yKyItjUhNRn3wKb159mBFMEXQ337ut6WMcoYXQ
TY0R0paMZIN89nPKvn2Cura758bqoX47j0zQUwesXu+X1xmqDTC0YKAT+ltADt+Y1mrSmijlnyCQ
LOpYhKA1Yq5OJ2Y6A7HDRisYkYm6l4vACm+vkHK2ZDiUAWHLs9tI0nC/eLYdRcLv4kwRU5eFqLEt
esxR0iYNclDLhklG44WqsgieMLFp1MNSZGK7hyBB4w+W1siz+2SGSTthYRvP260vyBPTmWj8G67d
MzouL8zpndSodcXTDYRgkaY/eRTabT6WGz1Nuwm1ORBCz5NKtDXRXOe95EaMdc1i5Ykpe8WQ6+Xy
/LwDqQ6xCM8ZWkiW33Rwgx0tiCXDH4siX3gGbnVug7ZBATfz7IjkreYYU6Dg3hZ/zvfrJhS5wO8R
KpUEXtzgnJeUP0Czq4vkms6uEZP+KdiCS0bYV5jGPdvLCqBJ0Y+B6ygkjrc6Kw0GjijLMxAVAPgs
qmor28opGSSIKLUJ9cCvh+cjDGrDMq5zwDQ0HeW6JLkIC5WJ6AMath/mjeJ0Ql37YBPW8CL3CyJy
QhpxLpXCP/O6noGcFfS1l2rDuaeH99DiItFij3RDyCaq2zkFOwq7gxO94svc0quCd5j2RUrIOYxX
5BkrNVib3qbFKLrQGhiITgQExj+UoqT2je6RJP4PlH/VRkGeGCrUw30lrChWp9A1VA/LP0txDXyZ
LfgbxubNP4HxlStH4XRG1bgG/39PUmxC+2EOKXWj3G5BHBJjfS22bjTW+Jw1f6m2Uc9ZTQmKFOHU
Y0wGc0PY8orNx4U6n+JFH6/0Q6tDAy13IBZ6X1dukf2gSNmOu2HFsq8OWZu/j+BJcPHeEza+xGtg
+oEuaXOLlJj7fSlhyPwjozc6apWEZlGTLX0yUoJ0et5XdpkvL+CfezI5+drK1fNe+uCSME6aQ4D5
IODVuw9lDoJSUCNrGWVhvP9P2N5GThhmq7DvioB6seIzj+ij5lrRKUpp3E5FEnegIC0rt7oi5+jY
8FRtJnoT2cZNj+vqFia9POkBezyBUS8YN1hhKuPmlshfAyRbv1gBDBypYgBBwKtBxm39dC7ht9Fb
XD5fznkWH5Nf+SFrtnWihQZJgEzNHzoG7ozaKk7+DwDpStEv1j3y+R9euUYiN1x4HG5sry5vmXRK
q53Cy7Qb2HkFV3IZlE8R37ymzO6pyfCSbA0J1R4ou+KhQw6JGBY5abLHxnKKwh5YPNQayVR69uAG
jTpFl/Yi9lwTS3NUwoTeo0jKQmbtfq80UTDkz1rP3v2BexuN78yOXjU5SexTOoSm3qz1sKwjtInv
5seREhs/LHefj9tpopW1f/68Jn2wjqnN1sy//FbZ8EmhMRnx9SLFarGi1iYpfWevAEoTU1U44AZy
Gml3l9fguaROIahw/rUmRsl4oKS53m/CN8R0qCZMBxehoE5EIHfUVIka1bfQihqe2LtmsjpKcvX9
AHjRl/qZSoBFeaTrHZ0TRlOV9ypU/x6YEfpzdLb6WShR1sRJUYWZa3TpIECfddifn50vpA9iCKki
J6XFUGeDPRyg+3k+MLnZidrpaVlLR3jjay26tXv9MQVdpJCEcnYWJ/3p5+1UYNGLWQlhOwr+Mj0D
khDUkdijaP8vOJkAI9QV8a8q1kJ6rIe/QUnOm433wy93uMZBncjD98Dd6g+zlogMBnWzgr5jojyx
Ucyo3ioCYfQT2SACLauegMQSC4h2tmQlvEuLbNDJ3looLATF7IDDQY/kn6V45W+01SOp/I3/7C30
qlDa2n9yOKMZSAYBF0hZYZJLA0Heg5FPUjhr27bXwTtthhhBF6BBkGgJkW1npFlYDcrvnSfJvZkY
oOU7XqIKrYubOvEKjMN/WuMdr6TtFmbYOO5e9MoHzfTT4qxfNTGbwEZvGFuaVMbfsyjZoOd7wP/T
PI3vg24WRnRcwcminYum5TCjCo0ZY66dE/VRi/gC2pc61qPOBA9xRArK98dcJv9xLlrYWpo6b+Ja
j+TIHqRdhqZdPnL2jzn4GZXSZ80DEBFffA41l68fp1sITxv0jbyMxk8vFzy5GuZRHHfdYPkVXP+0
BP/NmCZnEWyQiLiAKT9FiZ/UHARtK1YiAeF9P489N0L4mBSRQ807pyG9tO0kiyB0xjlC8jIvRA5o
0eLpRspnjp/dhJvqHUUaw9uhd5+0mxU0p7syU5c5A7ghZBHFYG/x3VpoA0mam5KkcjdGSULL4Naa
/BTuoctcJeqRKYj03QOZP+2k4GovfpX3uH93RoBlNFOIveOYjMhE+D+0Z+h9+WhHRj6OlA/2CBJm
sC6rNaWslr/Qo0yAOdAFditr5e97Js9ZDqfKQaB9OxrKZ9uoXxAMykvNHKsF8uCn7XlGlLAC0HDl
aFKW7e+kICF41MVgIyAFRStSxx2xwfk8rst4rr3U9JgFtBXIR8U1jgaGDbLLbJQ3DJyoWyS8ju+0
2g+NGY7909z3Hu4vXlH9fFo90MB+icILhp4UkfxzeoTuYgzPSUs4srHibi5WYoICiYrYz/VVJztz
d22gWaHATWLr8BShK9U/yPhz4c9QgW6a6VNFjV9H21ZMwQGyi8+w7F/FQIJ3vyyKgllN3FgA1j7b
T0XTh8kDrdQhzV5p469pf5eAKobQqlDmrHWp9jXBFplcoobKYYmrRzsX05PIk1LTKSi49kPLkFD5
x/SPGwkH4IBlQy+iWj1q2NDWOfM0vOUCc4saaFa7N2VSpWP4qGzYa+5DlS3Mf3VRpR0mBnBGkdpj
dn52s3m2Tq2n6BSsMFO1LJElILKQv8b32G226Es3wlgMfk4fBvHIAbC5TfBlF2LyBylKjmudhjYL
bY3dREcdheNxoLFSTDezE5h2AMjZXQTAByoGRNZKf8d03MJSLz2cF316futrezyPXaW+6Y3UEdzg
vJRY+CuzcArRSvHMH3jxTZgJ1nspNFmpH8DTJJwNAwFBmlwr3eIG5tKLY6UFOZF5KRfWccbZ/w4D
bX+5c8AQi6A6Tu2qZCWbD0tYk7sEo6jpWvGXCuE8XVzSm4/j/zseN2GGGoeQfqOlZfsCScfWlkqs
ZMbYwk+y/SS8BunHO1UFE6VMmJL+LaZJjM8mC1zuAyDC8LpUGjIyq8PxlsieYfojoHwCf++XnmrQ
S6MtVlIfDltjb1LBpPqMNyzrVR0ErKExvXaRuYXUxjdRbTHP9BPTUGSZ6wGNJ7Jitk6gSUZLF4FW
bRBlXakG/oK0E+mY/mjW4RB9lI5/pCKn34kPYyUwwdUqV4JGhAcnvFHDfLaw6LHyKFFWpgQVp+5w
CGVLA6gif4L24xIxZ2zIMjoAm+CmoyMkdyDSD0ZBoy2Leedclup54neNNP58j2ukbNU/JFAfqNLQ
w5JQQwbZVGtoEPJZVn20Gci/g/qtGaX9bYAsvo56Vbc1cuZaf4Nn1gwWYi7bM7kRh13RTcNk/JdE
091Y8M0eV0Ak+cnxv/72oMMqSQkIINgLzEaLfb4qDZfV37/wy2PEGw9+2raWJPccnuuy6cSaJsF9
AfLg+Uecxrd3D8BNpBtkr5zQJSrbo9s1fJzt2WvlkauRdnEV/lhfGuMUJGQGZoriO+5msd5nwasL
LUgRgtbopMTpH+yC0SaB2EUhwnU2ymspzyUMpayA2jqaEo8DC3jE/nQ7mA1r/jHEz+M4DD98TKf0
7OntKQOhAYQq4Tvwwa3G5b7h+03rypb+A6ngOemjQZQj31DfcVkrx6sux3jPU4G2n/FcBZ9wxvJR
ydoevU1tmgI3Qcs0M3mNBb9Y7JRqmEg++rzY1Fvz/z7Q+W9W/h3J+SrCHrwVLxKDOrz1SJQfzRJc
k5/c7jxe+hOQOZ32IJOTqEediN+CXjGY+0y3riUdcHVPKp2E02XY9oQP/LwZCs+kF46tpx/eqQqo
akI+pO8+RT3neQlLfXq94HRxl9UXmGw7XhPdQM3JSLe6WoPDjBg0rokJF6mqhNOOMocLOBomFYxQ
P1Fj5A+MkoVfi25eB2ovRv/84oYsXLl4LgMgqEJixV8Ci147DtBhQc0LRQBLkoUuOdxaR7r6ocZj
qsLubbu9YitJ37zGGYCDDK6anR394MDiu4b/2OoC2WsdWBjejn7rgfYkTj2QFW1AS2jOWoqV5CyG
HSn3lVEI8oYJ9G0zki3LkauKqeme5Koe8tA+01cVSj5lbFfb4V9/6CGhkDHvngksjx1qU83vayIN
MRpZlHPx9G8VrgTUKjh2REbuGMRxvuhT/NdTi2i3ypIOMAlx6wbTzD0YH7O3JOrpNfrYiHCtXfGA
k6ddvCn2yuhkpwpEgA5yD6SNorDLnbGKRgik1bPiJBdNZpLPLPSdoMqUM+EzBOMzJJWWfaMfAZyq
KZyQnzbA+EU0fs89if2zZoTxwx6A6GOU73Zmu4BG1G2+OPa2KH0Qy9vB8BXFGnDfyzxIEOw0CXzi
GxczOgp2gq+SAbNCxJ7FEQ+7ZrVQ/9LLK3CABEyrfrrDsb6GlOOKnTPiLehaXlZzPyehMf/Xh60g
PPI/5gliQhsR/mzWJPDSyixUk8bjXPuutqvQieYJAo2SwQTFUxzPlq0FFVW/rDiu2MJyCRc/R27J
Da21aHOyDG7Ea/Sli6g5zwMNdST/i7UgNNPkeX0TSnMHH7RtYjYluSWB2V/wbtEVYhIweCy/G9mj
6LGZTAkQNWNQv9WVYDPmJ+zqzHeiEfGu6Kfeq28NnL56wM6V2MUv+ikf77huxFA/1ZQHhh74p2YC
Qv4lDbbl+KpJJIX31CEJqyrLmrnYjjxIfzQ+CG18nSdBu5R3vmaxzVR0nE9h/0uNH5G3kZ4HuiUk
JwJABU3gLy5aViX59G2Ghc8ATI8AuvBo8lLEYM9A+Ct7rpr1oVPAN8i7r65PCHFC9hUc1kWPXvUP
T0wTkGNssP9HfWxzca/ox3dcVprQGuec7UpDZgj8J1y3dBzwsXxLMqU1pA9JH9wGbJYUL8qqUk68
+Irr/Xw6MpfOnn/Rd+iHyS6J9r6Bb0nrmZMSwTM3nUQyfNGLNNkQ1hJZz+hK+lA58mCjrc9NlwqW
dVEVfGV6qd3Uj3Yc2tnuxAss/KZbjF8XPAdDgazWj6E/oP1moPMQYCC9SIGrlv8oT9vnpa3gk8PH
BMPt4Ayxh5CH9CaJvZGj7uE4Nn+wTZysYXCXOryLWoDFVRg6gHpf9VAJFM39oWjk4+Uk3JaPzlb4
zQEaObwzFbjBhj70rWqE5jp7+8DQsdQpqVNj6kyDZHP6VIzIZqeC1y88tgfKqFbdcp3nf9kZ6WiN
FyqKrl2syzfFPkgXcK8U9jYti0n5N4NyOk6aKVVy2r9CGPKQ70lL5eCwwz5vkBn+3f3KfEuPAbr7
BU9KZzNOfSUbc2AKyK+VWiZRLeRSSJv/I2dJlK+p/ay3Bj5WAudj40d1gVLpbf+I6ZLKw/1qFzcN
63n+QkeTNkUFsrywElJXSzoWQ0VrnxP0U0y8l5q3ZlQQKzkQrTwjgkNkutLJWeHIfEWFl+GBeU4E
KyUhRUxzJLzy7viCLH3/lOjLgTQMO++WpCIjWSVBXu30KCgmfrIv0FhXe7WjgdI+SQ1d7Hf0f+CV
041K062rcR4PmKHqs68SdAoo/j2k4B5ZaHpdoHEmEoRkhLtOV6kslTNMtoirMrSLDltiewR94+U5
xnySnQmFjvGvclMCXOeFDOo1dtxnqeZ0GnnWylyQTmckYgvE6sYcO0qFhnCds0Ve/bg7zy74lBiG
KB3EiSDEHFAV5vsRzyAV9X3DLlfbwxS8Rnz6gAwUOgYm3O675If5k9Eh/pzzjL8ft9Ba2L1GBs2U
QHu8oznJk1fJUKQHokz8WIEOtlO8pJHpqFwfHChL3JVoOEzbbH4B7Wd9SSlGA8t/9YnhE5l7Kx4g
aSIUzaO+LFUDDc2zXmccMiTJKQ5rDyntjdleS766odwp7mwVEXSVkiZdPvo1lYJqWg/hgU8GKcJv
BdyLPJQsxLCSg6QTq/vLOjqyMx5OA6lhrkQBZ7sCCaNs7pvVM/1CibgKODgebbKqyRI9rEjD9wPq
MfvbBDkw5TpHJoc+wk0US17DHlABWifz01W5x+isUjFpjzufn0p2Z3h1iIbw2hpiK0jdR6oOrVaa
v9pPUl6eKNnlx7kF0TF0n62sYmhWQo6xkE6dAJHia8ycTiUsBwnECYhUkfIBDGlIMqlJez4pGzzb
06MAyoHMp8LYw3WlWvrF6SyA9s4K18I603YCjsCa4hT6GBbwvKuOaWxunelWpOKqXFlG6qLj+hQJ
2+HExcpekTmxFp7qUUKj6VAjetjAXcDPE4zy5d2bl8L/rQPWXP24nvwFEmA5F7Nl4Ym6cEdWxEIG
XKXoNAmByyxKOJOt6RMhzGAmNrHuUBvc1OR/90FQQR/d3PE8kNVdjCuBCD0h1HHadOC1xEpW1Ubi
yYsKG1pNL+TlsGis+8z7KGrftcVS5rsl7U1Di8mIydQNwBXRg04iNVqTM7ZsYNIqvWj0wug6kZ1O
c8peu7zEG1MFIJ8Zv3YrZo4Hj7u13HLbfO+akM17rs60+271kaOEQGJ7MciGSOn+pFqPqRajm4yu
INuasnqTB0/SQCcIqGSXG/3kBR0KhIPcQyZIOtgNiKdZ7ss9mctheLA5ztt8xBBY0cJ0E/yyg5XB
3pwBqPyVRNkf+sjkVFFADbc9n96y9LkArHWrMNmi/UkuYtX36LKyTiJD7+02/OUdqest+HxeecA3
gqaQrXH2IrjY2pT7iwXMX2p0PvlwLL1FWl+WSThnPGn3QimwDuRhZXzqB/uL3Carz6Df529AMkKO
TuPBBoy0gdhi29e4MA58+3nwxsD5ETk9IA+ju5Vkdobw6ho1W/l4PPOtQSw54s9QOQi4xfVWIIm4
giYtDOjZMCFEfoET51KWCCKFiyyKBc+zQlfIVR62U75ZXsNxIdMi+J/RbRm/yZm6V7J6pUUF7a51
ILY4ykoExK0pFI+2JtyPKwrA5QzffS1QQWU9kkGxlUxE08llpVA/GuUkFxWJR6dMIbcVpXDMrZhv
Fcf0BX1NMeE+UUepQnU29bln0OtbOTdRQZcx9fhF80gBQ+3br7QGisWROcRETTYSCTHX3MlGnAju
Wx/KvQ7exRjk2pup8FGkmz1xsXyNAK2JOUvb8s+tHS1zpqWiwfK4+21sx02XmSPOK/MAebpI6QMB
1rFTjz+w1TKiHtHd2PRnkI5qab0b692bnd/gXtnhTIxKG29Ia5dlNxoRfPcLZ24NNVKEuejgk3Rn
zT3ioRhuYD8aJiyMs3xlLnF2cAX8GTzLTUOfMaLv6BQKBJ16AnL/R1PbeDF3gzd92zE4k2v4iDBa
HWgLcsocZ7cmTLj9altR9xfs3ALXr03TIn21DJ3la0tzMKrpFmNqLReBBWxhH2Anx1scvugZQFJw
PAdCtMiule8xFeHAmkJ6bfypY/KIkviMDyaXyXk1fvjT4A7DQEmIisiWxA13LkeJbcsh6Obwfhc0
7QvOAk7jjiMiwyBSRR+QRoViYBelWKP6j4iQTCXEs9FLh3ud16pc7m63AfpeqALYr7DmqCMQJbhb
dUOuokVdSKEgTK8CKpqwe6vUJr9T6hE5ETb8F3msKFmgBhfBKMtLj2pdXrZT2rc1OsioarI+wTEL
km0jF5eNR8qeiGWZ2sEP8MnhKh3pelRJGEc2uUv6rCjmLUk7jJVwgHh+ObYaT19fQBl6u0AXdl8P
+XWCgU/ORmze+6/j/SCH5HV4O5W8UvUlbd9wQd0Zehunbe4mvCZ170UeOX30fF4lMadYKAZKy1XJ
aF1Ufy+QQQ2gnU1zxSStrF7ioHpCnIFsk4fakBeN90RXFD4EZF7cmDS7yyYlO7HVtJNhq5540Yu2
ue88osJ+Q3Ym8usheFUfNhKgB6nXu1vqjHgneXjMsgkIPneee5N5K8KLHPabRPYdHvwSjiCz6n4e
BP0A/M2EllLaSR44n5LVlOhAcHrmF2BdGwISaKC+3sP2cv/uvFiUnpK2T+Gu+vyxiVTaOsdEqaW+
ChqwMViswU/uIXOIjjS2xsJIRiv1TlVyi9K66BcJ5W7mQZWq9OiENxfBZADtartbm6HIVqMBOEqN
2aXqjJwfMTiZoNDw0vxN6u9Sm6Tv0za979y5KSoMXbLeeuBsz5Yi1V4fzDv2afznJD2KYXcaDTrM
Fe6KNtMEV6k/TCDlvBatbB35AGs99wd8FYnGOG26VcpChcwPtfERfiCGb33NanlnMEUS0MBTi5DT
XDJhM5WPl/VR4JhI9jsw3oyBPXc7XhxGmMN5xnIiHYw4iPS9tm9OEo0CZekekE1oen60CZDlyDRQ
incthLUc86gXN6hR406WTgUUctmRXbKo+FwHmsnlK5nFZPDPbaUc1KhdsGxTgQQmAytPWIrUr1Ra
skcuwZcnQxmO8/y1xPYzuBStZEHPBCbv2e2RFITQWSHzHH/sF/AduV+k7iUyB3zP9CY8hoasSSku
en7GqJB18fhT3c6p0H14CKa7fVX8fI6CfMND4NYOxTa4bgOIiyonwjW0YmfqcI5P5i/3gR9N8IPR
rwgO/qyJxXVpL991QJbfXrgyYHkCnR8kKklS3RRiVSZRLbfqMXFpEvi2dcGEV5Xf+QPu++JH45FN
+4agp2nHlPuejW8tOkdaOISWWrOe833pRbuAgrnkRgjGbQHFfdf2gkYwxf6CjfSS+69nj+Unuz7v
qnOGvaQ25wy71KUL5/+4HIwSb6H3/ulkgoSqnHfHU1xjkXvMwQir8yqKZ1ekqwT+TDOE7CWtPYjh
582YFZbMrWRUbHn1mwO3yiT1/2sXZOqRylBfFlsZTBZmZFBzjd8NCjYgtI1g6S2fG+uGbOzUOXo0
842hd0SLcCSYJpHfjWJInpY+ZIEd48PBRbjGkPrWj3cgHS2bJ071ZlR5I3+NmobiAXgSreHkXx2B
jXoiyqwghlbyXrU7mKbIJEvj5VqBS/Qvc6Q1L7rfvAHwtL4BjecTKZ9f6shQxs0dRvISz1g5Lysc
tJxVHLuCS8Jqry610unLZowMhVkVzADErzLv5xXulbI1Kmkx4rOQuC5vZLMGx1vL/NqXWPiBE/r9
Ri/nfh1fOE21DSRPaidoUFaLsI8LiNXIcL4oplQy7TWLeyZQkG9ucH7HkPM6Cjw7HDzJ/422XorR
P9WB0ILVa81k1PPGgoRbX5KiJKWfdQqGaQ+sYPTPkBzscWufLtcln2IpX2bdtLnw26PJHlVOZG1L
4GOF4RfZ3ZCVwanGtmJo+q5NVCNOhfZXsysN4kKeqm3ENRso1y99aGwrYe/3FZu/CnoeJONm95RY
/iH5bvsLeqCvfLXP1MkVsPspm9xa3tsp7iqjd2W1J+n3HNSfCyJgCkW/JY0EX6YrQvcM1/mQF9MM
y1WL6SxhULpbCXlWaN8VwanHEyUxDBJOuufbOU7O7wvvJY+4DmEHRzn3D2euAqNTpCNKQ/FSeo5Q
CSOlS4JsxUGDiTSCJyLBS23fRBxFrTuBDhIb2t0/pFFcY2AbWsJqNEL6IZNRJyrZ2JTikk9OluHz
qCaApohtZdljpYVX8CwnHLWr9vLo2/meGU9s5KirYifcZpIfp9aHxmp/LQ4TrRDY4WddSyT4PPrB
nC9EG0qS58ucgUPz/yMq3HoOVLg0YBy1CrnrRhS7M0UrCcCKxdKFU/WWC05eQxeT/HfNS7QgdbXt
dTOv+geis+ieYbyIgf2F4B8bTdZx8DzxIK9zU845MMz91o543KPQO5BjCJpMsDJf9pb+xSZzWpY6
iQP8QqvqT030s6vxP0rMci+qREOIZ6WWjEJ+CjiRwQQAteUxxkcr/2d5Eq0k0nc0qCCyDCfnDrx4
m7ApbQ8jj9KHkz6RfYycLtBH3uFtGH9K7mvdqXoIUFV2GIURbCKDKBAJorfQHC0axVfyr+FcVx3H
10XkOwZf+pWHMS6xVdQAKscTDFvP8VUgL0EhuAs8EuQC7CtWcCiLsg1Yb4B3j3yqM8em9QKmjdZw
akde5ECjLSaiHSZN7j0YN0JyPWUvZ+W+y65blWmnbeCjXhxMT0013yAtzpqw2JgsgY/TF5t5rX7O
biBhSCzDvyVlijyQ/M4HsIjqZQkpxctqUtjdAoQsA4lAd6zgL/7JnlGLeyTCPmr1XGTUi2jSzOc/
nRLET4x2lEPBp5jcfa3WRQ/tRZxzjZ9UYBvUV9mDCi4OU5+aYpmeRIF2nEOyOeH132jtADs4V04w
0syKgC2pvX9nJrd7JHklpGjj4CeXxAS0uR8tNwyijmLha2tqY9kVHiRM8lxNgSRFAJfojGW05AK9
khb0NuEzZsnB+mz8bDxswB26kArdf/IikaISSauYyFqIMWRXMLkO4WULmTfUf1PGkF2VQ+JMTaI0
x9ntXO8WtbUhHmqJAWPYasAppXHcHytTwO9Ugyc75xu9cCXngYeGmNcedjtvy94k+Qg7OfY8vNQY
fQTRp8l6L1ZHJaM24Qc96WQz1G2Uk7tlGQjRqpSGgOZViuhsl7kN73pYWqztk2istN/KbFgtJ9fa
xbIVeHyZl6P7PPURP7N0mESTCiRSThfD/SHi+WNVmAJh+xk3a9u3M1feBbtOfenAYLvALfGwAqQO
2F4WXX0fE2kjgrrtxeCfxqRtmtlWYMUsgiSU4e7gEh/d4wJOdNXYvCkf3axO8ienFB2+PzAzXqdv
iEi4kdoEKx/vpNLq5Mo2PPs7soM1dSXHI0KcNSitelOCwyD295DsK1EMEsjYgsM8CkxnrWvm02Po
QTKBtB+22dbvy6FGTZhgUN8f+Qzxj5FxlNv2wYjBtwJ2ZC1GcvqwCtf43gkhPpmzO3Bm+iu5CoU8
KXjXlUpheX4rQHZVW3++tgQpLblNi25khO2GTDp45lY5YbGj0B2KVNUxZncEbNKLdQ5G2Y1sPuag
VkMJmSPld4dMOoyWG6GTaLsPrurILfE9mNeUaBLi533xEDOLhRiM4Ag9hJB20IIyAZdeQFVNVkMD
s8N1o6Hmy/R+i72yaZtNWOgxEFrlpsXDFTEj82C2fNe4SBImdKDyBlxGqqFJzzcHtLOmLRw90vxV
AZTlIfMqLCds6e/S/HbEKjQhp0ch+omOmtBDkX2WyLU/f4dvDiZhjkbLZIEZtS0EOhkb/+Hjnuf1
h626Gnfgdal15ZY5aYoFGtREX1VlT0NTN6J2jvYMwND07JHWrSAsowp/sX5ie7zE/Abqw4WPxCe+
Q11kCSDMnWRLYCkDLIp5CoQvVUPlWJ8Ed0Q1bIfKSFkHkx9Y1wISzM/+0201dmm3TLJh0qcdtDzT
kdD9T+DYkNgolKx6oxOVO7NdBNuq6s3n+m6Olj91F4dwipvPD8OcD8yJNeml01kTdBzOPvhqxii8
yziEGGstabgSZuVog6jqG+OvRXESPqmx+j4JDCm4i67byUwhZdb4xDyyW7Lf+ACKkl7VOBpDjy/Y
y1YgEpB7xrWVJJFk/rYQKFqu6uFWmUFU8FJp8YhBMEEHt2AO4/tdOQDiqB1fW6C6LX0LJToHnoFp
KHc/C4AKEsoJ8UjGvjrkWgpeYZaAYBu6lUTCOJ7cOIeW0r73n21wNdc6W4LkXZrpkRY2palqWmB/
cp/A7/hzxrptcZMjkyNcUnn+vCwY5IMm7m3ZjKKdWdzzfCuGdzwYjxn/DCIW86h90mrhk6a8sq3r
sD313u26j6398D3A2j/pOvZ2bEjukSeaamkjxwfYYgSLRtJx74ZOH0yDnGR7q90NNgVg0aE/r1Rp
fDYgFbo4iaqWE54NAJnHkWFcaFFPbgT33N0Z1TTE4CcoFgxulSeLjNmu89Prv3tofEEoaIvr4Xud
kQR3rI6sP5XVW81f2OrBG5TXWi5TosHnEkmTCZQkJgREF8rTrZKjcHZQQ+9i3+Etz3xE9Y67pfYb
67F/rnYajuhcLFdEGB0PJRmafvNSUqTlma7vUSIPUJSr/2ba8MTJnBM4fy+dA7AKntU+mIzCy3WM
AZyIbrW20xliJpdeHt24cBE/kD1DE2V7F2J1OWY736Prdi+lnnOQ4Iam6M7bw9hhgxAWQcYO97N9
EOD30WnKyCDY0AgO7om8ihOPDnomlRoTEIT4eLDCrvWgaDF8PZQeD99MWU01qK+FeByLPRMM/pvF
78XV2px4jml67GYMaARKc0h5re0ngCz+nJ9R97sd6f22PHlHDUllR2E1txHICmtv1Bpntym0lhKz
tzpCjozXYcobHVc8IdiGFDpFCwbzzi+/qD4O3lfT//DsfkuD//FntZ7Sw1GH1GlnoD0j4GqtniZn
aTQcvNZKZGSHkbUFJFCYZXpSjvwHywuxXkgr7o+4RWI3CD76fYnOvPBRQS23vI4EuPN9gO+eGGjR
b1OEwhFDNzREHFuRCxIrs533Xs5Cr5A8YLg8B3t+kGMkwQEm8JQCgitSf8NkgQF7EqjnP34BE5yo
y4NtrjsXwXP5R8nmRI7qjv+cZ/lG1UiJTI5YaZHcRptyAOE2g2bL2e5cSObShnbWGCccI3+S1yt5
E6XVUqkcZAnd3o9wB/u3Eac6ywXyAB6CY4/tOsL2qIvFRzVhJD/H0fyOH7gsOQeNLwH51Mr07gbC
yt6gJKTDws0W6jlFb8oeDbag/QVMmCG2UU1RYuwjWRsFW8+NPerEjrt+KvfVMwkXTvo2a7Yz4vsI
xeusdaW7EN6RpvkGzA8uxi2dsl/Tmm/lf5fTLiJmhaiKor3o0xxWmq6oTyRPsZBjszIaD1W3Ez2N
JYhGmnZwAL06my5C4I7crYkrVuk9sdJFaufVaiYsF5MAQFsQ0XpYUCv5JgARbc7P2c9K10bUptwU
5gGiZJ8EgmB5gVmKD6ubKKo67PT5FM0PubmwCLvmiQSLSBGGUsfE4R4gpq3nRV9leATQGJGhB15G
CsPT4sWnrSgNNlFUabu2DvzAbtUsZ/1s5s6PlrTFl9Vt+D7AjJ2BRi8SKcAlMzqd7QPnHma4N/Yf
5EZrhEf1NyflJN+6rbtxE1NYB+z/mcsDnqpfA+8F/1229G1BxnXBBylxOn12f+zfRg2S8WtFGThL
sba7YysKitLx/AZSeRGbEiwFm7Ch1kvXpu7CtUgcEFEu1GMCJnr+jE0WWwLk1lN+sQF8N5msx85d
UHIxyedz6Wn1Sv8IVS1TeNBfWlySrzIxCKO150/rh5pM+wR3oOsgGSRpyNIDl2m/brrhwEAxD4qY
Rh0iT8nThpU1HMqfzf4uvDz6NYc+Q805GnEalQo3u1+/FjI9kJEADqwCOEppcgY4FYvhi5++ck+7
z96kfAxARuKUl0MtRyxKeM9JTA92HQk8BXowwtgzCas4HX6k7CU54tdzl709VlFZqdkQpZpUDL1i
ioaxvd7jpzKuefieiPPp5csuP4uK5f3WDa/nFKJLrMNk5LdmGkQsosbXHEsCXxOozn0fj1gqi68C
brH63zCBSKlIy2MRnxv+0/KhEJ3ZfW9R77O07v6VpfNDahqqrL/qlrY8TJdALJOyFUPp1xMDbyOi
htV1I1V2f5D5Hz2ZqNaDweTlVRZeva8QWDErwbjUZv68Bl0XBULkoJqokqEr4hISGUZkgvEag00x
hfURKZCNzZGEWCQA+JV8+UalR8TYHaJqnpDWuS2lkvZaPYUlMW8/4ywgmPFofylLfLCSEX9c0SS9
feow6HvvAWGTcoSSeQamI8hgJFSOZMyjSMD67wW6gZO3rAQitkgoXtaoM7L9plaJACIzIyd8inrs
OjQl2c37U0rUZPAg5OrAxsq4dcT8rvH9VTAW3nC9YbHMMoTs6Tg+r7En6d5eT0riBjFjJdqKCJ7a
ifI8ngRMfkEKvJzRIsUXrXbKl1jNqClTFpjNWqV1idzKh1sFGB7jycLtWsXlbAtUCiSSJdbyVCEn
/jFWcAtmeh83hMQGj407ozk4pOZPGEtoTqVxd3saro+rxQfbbJcamZidOsE6X3iIzfKUYcv6atqQ
nqlYdHLXFTMKaxiMCmmqHjd8GUurTZwlJ0fXdyE+Mu22i/lwrhghJwm3Lxv7UyDxZDpOd7FX3oaq
zWvnvRpX8NgvHveQLiSN8s09li6IKM3lFHqGVtA139f82/bZG+u/D6/hFDhVKnMZRXOPcRcSPLIH
rHp0Qp6iO5nfVWEcNZ6QAZAcZCTvfDC4B9DTDdtGOastIEsk3IarFacat4q5XsJ8guwhauZmmEDn
t3/orlFUhdPcJ0YArnDmOcFKr1eHFhUhagheb9YA7Ll2BjL/7KIqCGYgr75u9QHBEu8inuJKcMCF
3QdaLSMtIQ2wFK4v3BCX7w2z0i/ZRDpaPdj5PDTOl1frfZPVLjQuiaHJuVMXW4zXznpjazfVZWxL
6vXZn+m/u/AoV06YVVgIZiE+jBg1yE3jeSR2uwfoAAGNkuIOKUTA/7k56YGfsNMSk3IkHxhvHZBE
n0EKc7JLQkMKPm28aCOtQThF3BAjAo5fD+RlIL0vW5D5Njzf0Q61u2HYVFl2FnAgVa+5ucLXpFRS
JcB22ZwMYizEmjRnrMxh6JUE/yJSbRsUXaUJlVlaA0U3+x0OpJQeSnruJLfkpJgfr/TtXNDFA+Ji
UQFnb9KV0xzkCWRsRCQNkFN0P9Uu1QP65HBShBUl2Oj83SU1xVeeUzNbC0pYh30bAL3XqJLnblAr
PIQt5U7wh8yF5EJIqBUXo/0vnbreiZIc5HAX6/5XeoV2Q5pBLCzX1eZOjNwqkn5EMW7qTymuaFIR
Z9bOPDxcLEiNHmmveN2oHNS+y4/AAUhISpWGYElEW9WQ1wREH1VlN+o5i7zDy9qe3I9euJwACq6A
N278SB6lnt8yvcBi7bhsoQ3zDirSLPSdkw6CDgz28Jg9zsH5mRbUOwO3AWezOoE4kk94NhIgcdSm
cCnIHWDWitxMrCd+F6PDW4asvX7zQN/oezSbnTUoPo10POSL5gWwuLsEcMSUK9skJop6EjnEbdMy
HTkSCPbzXXfpPXHKqccU1Y8ifJhDKOWGdPmmPdhdygTPhC4KFpu58z7HRHsLSo1kDZmTmqMJiuw1
vZmkF8wzfpc+SCDaIqOUNVMm1JxwrVb6ZVU9frK+ZXxTw9AIyJj+KdYI58oiegjyOP9IQw/uFLAj
TcZhcQnj26Rdn2C9yLVOcjDODdWks+6DtZCCQuOZZoXYBNEYeW62C6dt7eNto4hm69MODgQDfy1g
b/DG2RGLkMxO4eIawmTludbkrlyuWtZXDB4C1sixnvANKPfAst+nnmEGqKbymCKNxCStmwZfl2DF
OAStoFjgKim4FJo3olUHwOq6Odn/8xSMY2+ecIc0sG4Ki37qoNp/NvDMeB0pvE/5dnQHv3j8WHCv
fT4IzJz7Orrb6zpntgHUMV2tOFvVvYsLtzPTIqKbSPhPyOp6ZQYmf+QaxViRJaQlEM9Tp9fddcON
aMeq4+E2/Vwikq2GQ/wySbooe9HMfdhij4GSIsU0JJloYVdzUj4kusy1elBgn91rSV9nrU3lZbJ7
7iNC4+BKutNvGqq2mm6whjLt9YQNoBRhP9j3ts4RmwZVYmDXo6qapbfFuX0BIyotKHk7FSZBDx9Q
0R9ETYNT8Xl/ps0804MX2AoFSF//zWtufxOAG4iQMxr236JHUpWGfqKcy6myWeG9VL9/UJjGA81d
oxee3dU8X8ZaMQRUbkgILa1kwa+R1FP+eM6MRdjh58GhejT+j4oosHSku8XihCY7PduKWMoS3bFz
QX9hsf01fNJ2h9DMhvEv1ehTMWkRDBpi94iNsI2hERiqpcRgHVT2S2kCCnBPUung/3fhrKCmwpiB
at9+k28qCw2Ztu7UV0WxPkKvWqoE7BrE0E/WJI0BkpRh2wpPhyI0MF6jsutjSJw4gakojUtcF/V+
rEIn/jXRyENtDwhrqu/Y53h4t93vTKSuo/Cb/dFxbxXs1vR0D1XLQgHUNQ9nfR+BUfDgJMoZwbuM
MTHqtMXLL2dIJh5MNPlUi6jUSk9fXir8B2ouJ972y5l7g6mjP7kNdfdkyfx3HWXspoG0czCKwd7K
ARWcrLaqbEsJKyHY5AWXI9oIS3S1SGghjKmBEt3vSzDQn/TBP3PEDyi1IqKeUu3/sfUbV6Gorztm
FosvaifQ2jRsOK8+qboEb6WeU3tHXEZLa3KoR9IJhtd4nJbxIzFLMwDQL//IFqi7zMY7OPOl0URM
AUW5ztvBghwaC9rD30Td06U+DJyWooW/cMmdpdwTakz4SDc8lgTSOeIa74WNjyXMGcrUlyCXklwI
orDMIoaforXZ/JhkdUttIR5JhSxwI4Yz82ki4nLq1qL7+/Y3PZdMXfpSNV0kg4kux00rCz8AF3Fm
aDMb1E0L8v0VOaNfAzxsTXgPH9vfUM0ml/ZsSWTXyFRHsQOJmkH+uvGiTZ9bi1ZTYuHD3pz98aEy
6Fm5AJ0bqLv+dtflzunEyEFZC3oBbMAn9MCL3se/vcknCHbzfTyf7YlAM1VguKefwos81Dx0i0C+
3VlBzLwT8qvoGF649+gDgcWAouS6dfq6Eab/tgYacdaKC30ZDuKTmzAIHkuIxyQN4ZBUHMBrD1I9
aTV7zSwLerFT8aCwTVqczXgZinjKSdoCIIuUXVms6l8BJLddCDZBwFVyV1F8A/hoTSSt3I8/1BSw
YvLd2PNDna06mVnn5HcZCtVXYKK4z9EPrJqtgaB6eB9v9p55c2dw9QgTwNtWT4BaGtyciZiiTBQu
RglliQxy7LopnFYQ98jBZLI6bgoXZSkeptlBPUKz85EtdHXpNYq1dAhUK/WyoG38wox+OxVijCEY
kUPG5Pps+f5gBRjP6yEmMu9QL5iSvoVK5GTWfzCnEIOwz4c/Y+M7gIFsreUaRyetOf9mdtcPvDsx
HxOEIDwlXIfNk1Vi2UKibxHbGoSUjjxmho9jarZYxmJsw39nxrBOeQMCon2qCwlmUrNRx/Ur3/j3
Q2qVsrhw28MEOiVqKiBpBRUBrBZtpBQvVy40r6ao+5tJQIyRX81kvtbR3Vm33LkzvzcXS0DLM/nI
MFh3lXGFYlZUCBoajNcSspcjy7hYKpP7STxCqv7uGs/jSg6JOcJ50pDax4B0eKzXAgVLqgRwe21u
j8706N11gq2Sv56j+49MRo50HH/QE6umNCHfhz8Xq0X1JC4p8c7E3nvxgWyG9rb0wlQCUKHAKPA+
I0zBOKZTGHBjFefyJM0tn6jV3TYOjumVM/ClR6pN0iV0rxFjOIF7pxPULfVsBhI71Y4JmTkxYj8V
8/HZcw5V4C7LiPy/Fy/QUYbvKX/FHVTfUAssRGo7IqKOSIr4v+SyhjywPCMy1outJZ3xvrYJ8tVH
BJEB5Fseo96y4RvRppzLhOpmfDy0pROo5e4mTbGtQG/1hhVXDjKRyINp19kC9esvTSd1HH5SKzU6
6gDu9pBql4LbbOsgUF8tT7uQkmoN5rmDylnY+anNHNksoG+a3dkdAYzOxXLziskW1PvrDckJSojL
Y17p6aPRWQOR6SxncG+Y2i2ZQ5HblHYIDcjgVbKk71gk1cko+VeEl7pios65Eyp5TQ08u9zlteAF
LcreABUzQGssc/MBfhewcmNFogjGBGCQe69IBHkeU1jFYsUMtqJggFTCwRqDNHLG+Aft18zgpot5
YoQTn+xqqRcuXhAc8FkT0sdb27GqUg7BQjtqX3c1CXukoCE3AeMJpz+BlsIbFwjEmordQXxGkiBJ
2P5cD9Ft18EaoX31fZG1JR+XrnQW+yPtJoFPjNzCb41Caj9KGxSftocHmqVe/U7JW+8EYHW0m0WV
/YeaMdO0Tcj2FV330r3KFKTKlPfu0B2SsDAzJ7SfF4NYLdJgEC1uk+UbVgk6mt2XozXQoPoC6DXT
vqJ6Ipw2M6hCbhg/pCYTmyugBOAhu0K4SRC5gM3XUL7k40sbHV6uT9zo7O/m3iqel9QztuqhPEVZ
9tChVRzGWpLaLlb2LiNb6Zfi6I0goA3unqkNlAK3QJJnN5vu4CsalyHIgk8zLuH727Kl5DyuQ5wn
b6kSzlCAKk31gORjbwUxakNJcSbuXpcwHrdMeHVfNAB1NcPL7QFPkjsj+TZTqgqE8t889uMNpjub
whbGrtXz5+MAR2hQfBfieTnrmA3hRQka06rFwYvXjoo/RQDsvyeCMFi/rD+BZr3FfJxCM5drSVUt
RFKBqsAh0sowA2uNh1UDY0yva6qwzrlMFbjFsBqOrNYZEn7y8OXkp3fDoz6WYIoQNwI8IQTvtG68
KYQXGPGM14akhiq0zPcAOVZ7SggEM18wI5WQtyU27TnBDr1x3Te5ld74mDhCYq3iXh9afsBhRUTP
n4Oqz6sPVexv2ULCwwJUwq+qoQ4jnEPx1ANKuerPfhTyKpYtC9F3X45PCrP2KqFKsy/EAJhGdnu2
GYCqAQOMhV2gDYD5hhGj6klKtgt1E65baStU2A/PJLURlHWH+Gn9QjfT4cP7hOv9pbqxxCMF+bHY
7DnnNMVju1jm+/K3S4wS7r9KgSv//moSZ5NFUTWbq8W85bJylg2lchBDeyFCEn9hOwPpQIxBn8Gl
C6CyL1/VO0sunxLSUpVweBOC+YH+pb0uhk1QqpKWsR5dxAcmJMwVAl4KoiH36CLYeUfJi/9DknY7
AQDaJAyVLdhqCEf4g5wPH3NOCvUz56MyVCdA6NiBx3fElkdGI+ziP5+YiORyR2m71lqhdETML/qL
btbOuHKT+Hw5QIci696p5JjLhyoqSMBOAmmf1sxglb3Up/mjyhZs9fRQttm0cLeMYRfoUR5zEMEO
D4rGT9YqeXyjoe3jc/Fu+lsaB/+x0UwCKfhaRII9MzXwI5r4iPQe/ASdcbD/abSnw6Aq4XfisaBb
XVuHXjK8wbuqWGThvoQy6eyblyIXlAx9Ljxmo5Xk5ilkGDPaooOETxRgSciRKVXLCTnRGAXR+zgK
AlkqgtFNJEb2QD351yz+S/LnadWNe5SJXpHKwHYh6M4qBbFwfPtG7i6qHgea2BRT657S7MgOwUf3
CrtYlrbk8sdzcDp5vM8jyFpePVSeWdv+7l4KDN0tSNffsN33+VsCHAcw6oxBrAi6HizUMDSUaokN
L+6qgf0xldKqdJod9H7WDnG+NVrDIWpOoGmjU5/eCtpIa+AE1ZRNpOYqdtli0pCwbt7Q0PNbD87T
xXWfu1GZn1G5d9qMU4/at0un8/JCtyW6lJFFfTGf4WZiLWR/MIIPMfOQlXn0FXDZtI2Er+9iJdbW
S+OTDQYUDQ6Vk/u/v7XXy1nmOMBKRhFg7M8QXqk5uaJvW7oqakKoy2nhl1paxPKHtZp6svbZYbs5
yUOHaBAZBieDAK7UgVXC1XoJndkO6+180Ej9xaNW8eUXrMw/vSnQ6KArH2FjDBDXbV9okORXQvdz
uj0l8Pr8bFphXDiWiZiU5UY5Vci2XV28BMsuuUpW4IZqNICdYczs6L4cxW/vRhkCvb9sFqSkwg8y
ShL73meo1nkF5FEZ5I5xC937vvp5LSpH5zR2xT9VpMNh1D0oR/yrwhgBHt7xQ6/XLXzSSNyLhn2e
sxnJ2ztMsFKSA8O1GjSlMzHg8WXrVmmWKzXPrsSM3hRW7m+wXkD7p+mbGNfZ8/0I2ghF/6Qn2WKq
WDpV8rPnHDTrXDZvdBHvYMhjCpsbac0SzbSJUKg/gLXmD48QcQCl5z13gdaoUAn/p31R8Uafw+Y7
4K9Tzqw0THKnuAuKvsAKVl8lGOPgBjvOsDmBPC9OTcqG8WxuWj91XSZlG0S05MUOoJ9MzUibWlgM
RsLxS5YYGZ+kLEwbEN/KjifYsVAFVQ0ptvdbGE9IfURZoWij1AlCLmP0EG6xOzwdO3oCDBYpLtNh
Qcj9hCpbf4DvXXDezmo1U+p6zYdHjcdNuw9I9le93FY8xe0DvEPXV2p7kZrxiobiiPFutC6BOFjk
wY2vpCF1Mepckx0i0vZzfS4gWYkpERl0Cxj1yglHF4TkSrjpGi+e7kC1/KXf7oA8rzncher3BsqC
0bsWtxPA5ftwMNKYbKSxHI2iJCSXdHggSsgaAsy3RXMmFRWFR8WhVSSTKzSZMuURRY6bxZgI8iXM
7NJ1jT6bgnn0FYNEROWeX1+euQb3uNfjLyKMjDJ1sxZczGEZ4Z3PYuRO8Fg3YSWq9wdyWeRN3o1i
bVA/YbXSDce2o1BonAwm+1+IFC7m+riawPXLHrw86s+BvGmv67YAeHoIB2DFMW60A9/vx6JscQOU
3XJd47Ese5D0hd5lLTaWB7/veTxzts7fuM1FjTq3pAyGbMtDDsJdm/a5Qf/q3L+UoX+rqomkKtmL
kQst9Db5Ot0wnawVWObMWkajRd6fqjr2sEr3j3IvI53Lvvba4AVf4lzKMmC959xNrxb97otcQuoJ
IH0zF6tZf8dSbcdzAsFjjZLlIt8QfiUrFveEcy8N8II4bSbmc/MOX+PrIpSf+M2q7HyRE36wsMml
7+Cojj7R9JRatEFxpnjfpSyb6W+7E5YJPnkrOxOgjf+y2Ln4ULk4xooesh1y5+3BR1NXuyVPnAcA
M8LK/ubr2eSrtaRsaYwvPX6y1cub5AsBFAue3RYiCqoh6Oyn0mex/rcmRN0HkEcoqY6zOj12Bnpf
BxIadqp4YdwCph1JMlUyQmcoRqKxn7OkKroJm73PkBGlaqr1BjJ2q8hCwKlE1srj3Yy9WBu1SSm6
oQnOdZRfo/hIf0nV/UF1FRgGdrerqWus15/kSQIJq0QYa572zENeaQCdZ7Fkn/oLfEn9gO6q9THg
lQ1pMFf81HtmiR3eIld4KycdbpGMAF6jKOdl0d4eZiRNjRPXMNmAc+INaKuk9L5NHPmE/wk7FMiv
OiDtoh9SeDQiobCEFbbfXlSyXRU/+WUkK0ypBaiF8bbyTRoNWuCCwrKdmIPqgSj/XiQ2YAHWuljB
h6m5TtPxou8v19PUW3OmIEKeKhWBkxy0OHLzMn/cBLF43A1eviopbHyI7UaKNX04xFe5KZ8VETdb
TVNo7XvDN18jBwcD2oji2u5rllZombOo5//AJDL5Kp83INUXwpvXES6sVzKYllLcbu/EGvo7SWVi
DAWqvhFCFfbodZGT62nMMdEjVGlWIRTD6HaQ8qMYt87sHFVMFZu0qaU27hNJnKwrYyC+vB29yz9V
NhFnC/fNoNbVy8N5DM8a/l9+aKQdNNcwBk1vYDrM7Hn384djeA2KZOuGU3LnZ8y6hrLwrFzpyjRG
KwaHdwgMET2KOxKWIl1obFMQR/64FfS9kL7E7krXCJoj6t9uiYlmkVu0jKV9y/CgwO9RGCkLynUL
uK+1HdyjoZhS5VBqO06IfRBv3Iw3M3Hdv9yRHynv9oFG6cPa+zdJkiGr56EykfuPUmbMbJpvufI4
YRXh4j94DD0B4r/KiQ4rmutPqrLge2wd/D7I/70KhURTxvZVXifApCAQiSwhbN98l1kawnqtW6e7
Pn51J3/DhBu3ds3rPsyyZLr9LGJQoxJYZL1qK9YR79rd4frivmwmLPRWE+IMX2DLJDiCLOhrBn9Z
lybuiRp68VLC506asfl5hnXqsdnKPDeSvtcVKi12G9WLyOyu7B6U0k1Pdqf2tu25m2DBNiF+gRz4
PqcLEEpCvUnzV9qY2baQ4d/2R38p7Toe0fFTjJRmcs7wqUV2xzNSWo8N6cqojZW7eq44A6m+92EB
w6CdIZaEqN8A7xMZ1SknxOdBE1FGz60Fo5oVNItfWKKWJiTHek0lCv5EgwhSNRwO68E7cGkhP697
HgeGic9lv2bla+ioTj7MJvrLbZmy9ZCkWTexGWjIwg6IAvZeTnj8H8Wl3Lvzt5VY3n8EzHu2TEQb
TXbkml5lm4J9HTIEFMfwNdxu5wtev9T/2+CGSR3bV+Q0k2FPm2Glms4cphpJA0DJBWkC+ccIplUy
hbWSP3Ir7d9ULMcz0D7IXNv0yFoXFfIE/RSy48zIoZYPN19RSN6B5CORJ0QtVTyqIuM2XjyRkvOC
8SePG3h/C1EV8jtjvUSILgW90dOipsEp6chgTSVc9/OdBCsDwH+uOTQ+em0jhD9iaz84E9B6h5sw
y5otuVCZT/pQLHMmGuOzENxaSO+KgcnR3GmXMAQwTwn6/dyUNk5Bmdiw5XN38gFMMSYFOhdK3Ulf
IxYg5OCEbX9v4Oi9xFZT0w+nP0L+Mt7zg32spl/+UXh+NtBlxejmbwuWunYfmxKZy2I5dJ5HSIMN
Oy9K/Ol1MPInunmpGnB2RsfuKyx/n7HH2CQ4f1qnwdOB86+zQbWJHF5PNtYLaWstCu0QgsYeedaO
AsqUVjIqwCgsvP7rzDHm7qHL/08B9q2xSI6NDtPCphdZRgu/3cxcBfu/AbiZ36TlSXetBLquqlMa
mlSBZ9fQo79B07qklQE68AVXDLmOihX9R9gLsk2Q4f7Ae8EAnJyOlJCuIyR+P3WVqegtsre+No6m
Bv6WsP6LewrLBvrkj0sEl9MG+mPGCTqTuUXIsalYzHKVD695S8jzk5HjR2lx66QF6AlsRHZsEFSw
b2Sp7uBsj1rdt4IdcYJ20bBjhu5XqxpBIj1lY2eXsMqotv+ET/jLIZrXrbAi2vZg3F8oxAerhht5
+nNCB690LBjcymOASNdkMpnLdlqtJDMjkdM5lWHkwT0Ad8x6iv3Gb99K2RfoS++bWafFkWLKDGQE
yhXW+YOe8AJRvp6M6TjA/6mIRadteamL7YHUhL4+jzKEGA5b1i5gxNqQVSYCAFhWslUYGo8vA9t2
vfowO6G2RaWdjuAvsmCD6F/TJy1bai7W9nBTJjlvhvIbfBkXRZTpHpIlwSLgz8p73CRulLNaGxNZ
0xU5h7u5TWmtkQhNfNAjr6VTxRvV1vu1PRgDEnEHmgvkKdLwfVVvSIcA3hRsrpMaYVGuFGPjh++e
EsHbhliagbUnFmvk4D6IkX7/nZl1C1NCCfOPYpPeMQZEAR3nzjwfbvkMJUfs7tVP2US8U5nVvykM
f7SVJ3sulMRojjXJiYg5rOZ4eMcDx17icSKfEmsJGy8tycrMMZK07sDddjgtx3IRwLWXALJ7y2uL
CjuKlZ40xG1vzpfDknZDbBw/9vj867qwBrdwgvehdAiC6eVsFtg1kVCLVFt6lSPqcFWqdRgXrQyC
Zv2UCPE9Nh+duJ7eKbbQxImawDarV34QJIlEBSPo4XJRQvPQ7+FTFaHLFwfBYMmxyhn4TILo2Ef1
jXjhN1WCT7eQcgzvNsut3SU8xvZbdbu6wT0BTKu/Ofg2ueVjBbK2y+RJKjErFK2NUsvrugae5uSi
kKIKdcV4zp/QqQD0nnCEBmlDwxNtw3ZWsp7Qjdw3JsmMpi1EDyrJUqm0MgzhUnu5ZfxTe+HiMt0x
C5TEswr8aDPdX8jaRB1gZMxfq6Oe3UrP8osPfqQxDM/iIPlYdUnbIJ95+x1PBylvopuQiF0m2UPt
DkFycOL7WDepV8XN+KN8C5YrknEGhSEizYPpkE7t69ideYysWlX9cSui6OcNp+76G/fp2Nah+1mY
u70x87a9q/UKheHbJprYScJZYaeBE7RgJjsGZoEb2D9uUhmcYRzD/TMhGX6lHDk3V2MK3zYmxJeU
CQ2MOm23Majd/f36uwyoTkpy4zWtN/BG4RfDdFqVR2gFZ/Hfg85qes8m0jWk/KvEpLgv4AwZsMem
EhcQr+pEf7K/5lydWu7X4tkb0vX1LvxMAUjchq+W98epZ9mxQhw7o7DZz9r+m/o/ndvvDnzC+m9X
LvKH4ZJTi048R2QNBNEmxHukZzT2uIWt+Zh464WjHKbHhcc/PyfOs9BP5MDkl+bU4AfxmcMkvssd
BwWakTy855CEYN/F6ytLPL7+OliNwXvIafdwQuhIXUOx5491oc17h7w5AxIheo8U5ErQjUeJfnlO
xAay1CI2Fn+afpDrQTQvunwQ3L//QZudTwNUk+E+X5P/xQX1KtCX+TIP2TVbN0LWSX5gBtLksMyG
lIg8lR/iQTzBdV2+lkD6w+EPQi9XnQVOsQZU8/8YBbpqrotfBftOBcRe8AjE1QEs5lCXjyEMQY3i
zWruOHsXcoX39mzLy2yAj1erx+yV12vIjxN8HFabEGFHPUR+Zz0I3zl8VjY4BwDH7pC3FEDgJ+5A
5GgEMNsLkKB//2geX2wVTk2ZkWVBCcwYGTS7zM8UWTanPMt7VnzAdBUktdQTpx/05rai+VVBepgx
bWk2/f6kyiVaASFlTc8RYJs0kgrMM7efbD6B96HYwanTSBlftR8JS9anWgqsfF8shhi1ybo/WKtp
ABgNf/re+IN4y6Fjt4ylzNIgNPGgOH6T+yftyraEny4COcwegnZFyCdGO7DUJ6+qdIwSgrk0D5lL
kIE2fYRN4eG1D72CXSb5RRFZD2MOC3LTC2nVu355oOWuTREMeBn0RMr97yG6RnlO0c/14JyndRcX
A68xy1hdZi5ZhXB4wnfIcRh4/zcWJFP5JV4uj48LVEmS7aRbx3rG+wk673i3T5nAP0SiCw4izYSc
LVpT2LR0LwK5aHXSAaIR/ADJfLde5Iu9+bbxYM+xkIsV08MHsROeWIzNuB5ZXBgw7Lp4j7Z+L4Tf
R/ftZyY5c/p4n8NcrCnAcJXdCvsF7jlKVypNDtlEZlaNexjsv2Jhgnsifl9BR+CSXRlBfv1SDWwp
yECjP8Rb84av6NI5eRLP00rmixmz2aR7U/biV+KadpQ3KHd+SvATabT7hIa/C7PIORqZG9U8MYTj
2f2Gz8QHeB9C2Uc4FlAJYDze+CCyHtZVk/Yj70rHhufGKktTHRnSMja37EEDSBifl6eRMbbOuhNZ
RsRPb3zjrz4mj6yNluM/15+GcMeVU7cQN8rfyfbxSfp79+CuOTNlpaP0alJ9/qHNovxRPFluxj3o
5Bd8LgTwmCxFMuxJeNwgYu5Neesm4ndE6vteZOM7VoquiFvyDlvN436PV/if5XSBIa6XlRLm9KwA
8jl9tE7KuwDE8UFA+xWdduPqCde05NxsX2aW384RsGlz+b6kyiO7xwrMoaQYZpWqcpauMDDsuU1N
jxnYrTnyr4CBPgERf3lHfR7/zGlF0guX8zyB7CnhFne0VBRJeX9UCOR2K2sjxCeZlPBkhum34AyI
R2tZXAFNPAIHfxEXlYyVj80rFF8uAYQoY7XKC2KPu46m1GZc4sW6NC8AKEkOx/FX/i5SyN9fV7DZ
k7oIOZkf2L8yfIg3nGTEP+bjBxenMKPNuXbVwzpc0z1RxCa5kExkiAhfPt4ZouDD+/dQ9mdd6yyq
jfubVpXHQMSSUq0Bk1yi4IB93DWG0Xu9Wk6EOcXMMVXPjlqsLACE7bQBJZDt4CU/vc6jOpFA76DZ
oMXlMe7j4+HBbMvHg9F3klFLfvlTJPM94bj1/KvnGZ7gmB79Jxv17LRNwjW/WexsVJBHFs5xH51y
UIey+WV9y8gEPTevPUCgC19K2hCs1m4SvVyFWpWjj54UbrEoibkeXxIpjXEXxfioc1BdenLe7j1/
EeODXEcfhV6V4DjB1bUSARJqs9EkDDgPzAl1AX8vkp1cKvsLP04aQOy2Z9FWnWJURiuRHW009uqm
bs9GwxbpgnjyVJ/90aAtweKEV7n6Npsp+3XvOJbgdCWeQPGWITqdmpFlgIEgPXewYd4sd3ejQsRW
tL7MrGoAJB0RJ6lU62eFGtAvSjLqtXbw7tGlP9d7PkSb0O6aJf5UPy4xGCvvjxJhwqB6/63EjDtc
wADpvDTUmr9ifZkd6s+FGoVkeIONuqtZtTe0is95PyAZWMIBRhjPhhORBrYIMkiaEV8mTMGmDsMF
NLoFhTJlFI+VHT6NdsVOdk+S4HZsZPBMvZSd2HNwq1b3DGW0XM3F7zMEcON5ZWVdbVBooTmZlP7H
/rG2tgW93YEyRgKp2lk8sb2rQ0imzdle+nu8Ga6hSKuFf4f49QSTTrbuhR6KcdDp0Zjb+Rk6eerN
RcQj1vgx2KzDa3Q2QobpxdH1vLPmZ+KXjE9wWyVQ8stLK5OkSvoQaGgfS2RLUDyTbYa3y9U4ZW2W
9ipTf6d9O4HzL8XsSv8lg4nHZ0M2bW3X6dXB/ht9saW5gHLNfopj1lYjHHhOut0b1FOFreYHpngu
eNL1SgM00H7/4ZF8pi56BEurgO38pnO+Dkr3wsOkjXoCHvdNn6k5J/+AgR7/4pyDNVHV/ZeUe0F0
6Vw1cK/nAJ/dkmIjf1q/S3moK7IUuWnF47cykb3z5weECEyqTF77BO2jDby94qWBy2ELh9ESacvn
lT7HqRfmJVMubnH/FFC02lfaS2kmkqX0F8S+w2xgGkYhgPcBuuyk3Qbyqfi0RkeZqYi1FjPW3SYT
u5hiBKWABVxIpcbRiKGe2e0nCB41Tk7bQJLDL9nidMsYW9XYiim/b5UfVVrbNd7o/RVahmykGc/5
Soxl2I10xHppMnQDXyLf2gO1TTfZLMgw3OhvLRsJeLz55GPcWjHWbNvw97TKXpfCEqxbBVpREicH
tLxQ/tZUsG6r1NMRfdYkS+hAHohRgf1J9yyJ82wyKnNMYpxVj0YIkPAgcitJsAaG6NB67ILBEDJ8
14ZLR+xckJZPyGv3vkZlNJ2H1IN8VM40KMpzAQ0RdvOGFKIB73q+ucqv9KNLYIiyeUrjG0VDrPf2
waKKRGatdllt6mwJjf821arHGkcSUmmNBSmY2qjuh41pF8RcgH4OaUR1wOTTB71wvp/ioZDEQExl
zCF18pQR8XGkVss8kJixXFduB59dgI8us6ZfQLj6nEjWw0QNheL5ZkH1cyuFA/oZxz0lTtoD42nT
n69lKZXPn/8ElRZLy9JoQEkuqzsAUnO59sDwHdKoUUP9MohRQpheAVj8a6H/rJXvg0nYt4n+pkR4
dx/NxeRVCjIP0K7yy3WP7REGXoiWEX+qnuj4fzCiaqOkPdfnJU2d465GXkAHP/NQvfKZGeWIUmN1
FkARCgqDNmOYXJueqJxjzb+qQewxOISa7/5MWjvQpgHwfpRyhBtfpEqJNvy8CQ4RFs5QL9hBm0EE
G5vbXTrYIlnb8cgwpug0OH05zRAnu2+pys4/4ij3da3n0L7omBAXmtlvqfqpcbJ/wfiXxao3LOJT
RF12WoYbZfB6cHeilC3QtoB5IVbqES4OiutBccoJx8CxxnTg9ZT5azzhbwd/w4sI445OmFwA3kAu
tSj6uI5rcFN8sSVHaB9ZEwVTQhWstSb9ULd8Q7qNB8c2TAXJkW5lgp9qux6jHhCbU4yngxgI/Uo9
7HiTSboWh6FugYJ7r97SywUmpUPm85wabk/ijReX6MUib1XNr3X8uUC2q+4qTGLE1XWV4F8dlfR4
wElGiat1/6J2vv9YK9AC0htcX9zj7kTS+0mwUiX7sCwMnqu3KdZKpCpLpkD2T+z8IuZPgTo4mZLY
xnwDHBuKaAnN/1cDdKqH0qaX5SKNg22HRYISg5HvVI3a9jPF/NVQTbb4DJgK7ku7UaI1brlK4Tce
twsYCYErZJvVAY9WuvQbYn3O/ZtywBGXQ8ATjp12x7mI4KArTQkNzvxuBNDehh8SsoV3eNeF/5IM
BYVyyzXoelWhlfouJ5EJtcupr9Q920zqEIDOLVoFqhTNkQAMWVzmCND6BsDYpWNWQT6Yg2YshDV3
csPvSwwtTmoxau0prpMeva6maeUuI9biBBD+pLV1s8oFu+qrB5VJzMvbYndEHAF9a1WvcZyg6G4m
CmfEKwLL7xdpDHR4LsGFEclGvK9GJDrQyO4qZhGdxIHFaWXpSGuqabZ/SLj/ZUynnVJ8Z4xyNmp/
vCM8FX5qv2T1zpJNmEvwzP9R/yxZwFNFUOPB5IbLecG4mrzZ7iZUMXdjLHJqldIsAE5pKmeXAvxE
g31VenKJteiGdRPtNsNVwFIrMprhVa0Ws2Jb2KKLreg4Brnwm9w04plEV40XAWtfyzo4PAoRJp79
bzyBoco0on8uVTh/o4GlFVZdwOTC3eELAoPj9GuBIubPmo9yHqvLwncYTpWBo56LxX8asKTVHYVu
ehutRsjcIH3tIaRpG8J5VMtXpuqBuL+AmJVVJ4oiUd7h3oze9JXdUZtorm6shAvymTa2goFOir0x
NxQzS3Px+P0+eleEo3Z1EPOmc4brjhyj5biAhnOqnBYmiYPmGZIKNigtEhYPUegOBjS2bjJ5I4XD
7TswhjN2oQxmD1qvwBr5n19UX0YucIr5u+vmb2t84VmCFeRnCYsbo8BJHbmy/+Joe4iUYV3fQaRr
nBRjhBkY6DzrM58JgfLwR+hfZvBYr2l9npg0KuRPPX5GGqfwFaxdgyRSpEdt6KOdlxp5iS2OOGAw
mggdD3aBpizEwUpv0o/uhws5ZUei2wGAakGLaRkXBN7ofU7iW9ERKnDnqQQqrVi7FUd3eatG58jP
oj7DvWLQuddGHN9VuemOblWJMcTv0qUZs7+PryqwjHui9RHQ4cz2inPAlGUfRs7WO2kwUULm9m9o
gTBD6sHUMszfUiBnA+wssJiQR8ycFhNXvNyvuRjeMMFJDPOJMs0JFe4ssquAxOFQ7qmvcpgDDAuw
D3XstiH5CMs1XdATMNArQelhfUgM6R2hBLrnc2kmdSsmXZYqdPMFBjyUphS6OM0A1UEu1gIGlEsW
LfuQmsc0+8ULnBdwGsI3Hwu1p93L+HlZ6VUzrUE3nERcgqJg5bnV2ZDRmXMxdX3N1+MkiMGFLY/f
+DPeYDkdcrH1XslPb5FFa6zL/ALzlRKEYR9otfZ6h2GGQPHAhNwKYZrs5klzAnB9IHycjD7wzuI9
8VT+5ZFz/XP4xFoWNEB7wYwg9J0DGDM+rmZQ+1/Gg9zcPT6rOyBTOeyuFVBRu7dXuPnQR63x59qm
CsPj18T7bTAtwbzocsMZ11QOlhTQedmI38B36BSjynsWDpU1RgGrj8tjAMFAsFn6T3t6E3dl25BI
fi8Qz5dbXy+6c/Fkzfl3070AbHSLzZnyn6PsIhR+8jIi1ounHObIiJ3PPUeC4je2muoZnFtgGstU
F6SW3QqcXZkSscsqwTQCG+miw1PqR1ejskO4SOgYzNWAQEQx/jzmMu36b1W1300vaxIwwTL7N14I
i8lBL1c7uaal8nuNTmaQb6eii1zU83K9HKcPA/PsjYJPSkGSmgRt8vVX//gJr+bOscx5T9TyNHA2
MkOJPwf0FIyjnHuC4e3+g3cJj7DMyf93s226zUdNSLLjGG7pi8JcGfZa3Dm4+Mt3wELO7aB9V4uM
R2gLwH8pkVe5toPLwYckNsHL/uY95NnZBlYqF7BUFbQUWCmxBI11bklZjfe3Df8cs6J/TEzohMt1
As3aUJvSyqItAwqdMS4yLk9WkT1q175PoO/JF9b5I5Iy+5oDcWAqNV4opXqt2l0bB1XGqdxtP0AG
GpgANI4O6HeFgWbsydFDQlus662ppzSpw8FBp1HRFUyn1hSLpzBgmCoYd19wkoS+bGL6LO17Lj0F
StFf5dwDvaBEweYFk5a4pwLquAL9HvgHv338T50LNzxBy29RT9f3l9U163fI2kvVFiXT/NPvF50s
L7FktpARGPyrBVQlfH/RHJvoww+xYFYT1gDrgajwD6AnGha+9P66I/F9476EGTFXg4VvyUuvco31
T0Y221hdKX+uBT+Gvx+MrwPBEsaKtRT8pnR+oGJ+eD7TvP3Xn/mGYwUulJuL7hLbPmcAQvx92XSC
kA5IwvowTGm9XX9w/ftAHTynx/Av7FNKrrXl93Z4TKQ9+8sv1zoQoEAW87Bv8Q9PRiev87YHUwQa
WVRAW7rAmLKlnIm8Ss9GwHiXSWClTyJ0n4pUoV+iBrPKwaGRemMPbAp1zFct9aAkHH17HPrE3SU2
abD9aOUfshGRS5Eejq+8MZEPS698HGo9z+GefZHkOMBo6Ld2nvjahknPm08vWpuhq26QSl68EFb8
FNY+OyuKgbzY024+Lt+vYOxPWsvAhp516NXeqxczxLWrz6Q+u2laLYKnjoRG8ty8d7B3Z+ZNbO2f
R38NyoJlKskaxq7XLYByuaUE0wivn0GsgMT5ezflOtkQU/Q/SmNaIM0wUqmKdWa4/d4N87uQiA9w
3Sd6Ib207WV3aZRccre8C0ZBNZKwLBdBq/pF1MoOG3jsDTWv6nXnavLAOKw46XuKq9LbaUV4RZ8S
4OzZT1JdjxOteUpemluRZmWL2AOLEhFjXt3HezAmTVj+tcwaxfzIj4U+nfZQ4D5E2e+6m/FvMJaJ
mD4zX+oOpGXqwnPrrKLqHICKiSGH34t00EtOv0e0xRuSSC6KYNr/K0DJ8pTsI7ZCpQ1l5UIFNJug
p3U1Nf9Ope/8ZLl8E1Je6skIDhJaW8JzXF+vGNDHLOj2ZRSyRPz8gcjdSrAc2TKUw2Nn4mXpIFW4
p9tbxM6Q8B7YxTrap51GKKzWrBT+ba0nT+q7vKkGVRTHeeZJBw7UWtwIHWhGW4xwsBP8J3QE53mK
fxItwlJJYVJXjI4RVLvmv9s4JzqbkSDLqMpPhvDqtA9FGqk5Z79G0xCHXAxO4IilwA3GkLuNiRc9
F2RDW8VwGYBRj1nNaQbwoEFT2tBrYLRNMZt1EDooKNonDMd+sqpHSjc2Zddi3MliLf20bBNysuLU
2CWIGA9aSKCFWLla+ID4bml91rjjsac29zIQsIAqap06+9NNc5bDpmTqi7+Lzbyp8pVB3MJKUu1+
2ipPIaVE90i9ZGbKHjbn2j8COjmB+y07EQ9zS86aen0H2lqqTLOt1vklzal9895M7reOKv975duI
qnM4k0bQSN0cZBDgsrJL4lQjm8qCw7oMshEdJO0xqjaDfCkaV4CqO6TISD8YlH6DgbcaeRtUtU+1
hdTu8vMkQYa0hokl8FKTs9ua24uvU4Fq2KZEqtd9lklV4p2keNhrURDbtVHIWJ4Gocnm3BI586nm
HyyUOHkfOvBzEypDxBlWhyc5eG8p1/Au26+yuY3GIGtH9veCWZ8FIAjmvQst/flvFEdERf7efMIT
iA01NJeqVM9AtuWEQoe1nr1u9a+uK9sq3pbz8SM6Gdgmd3z4aMKJ1LI3gtYgiByyvTNEBGh21XvK
dq9XITm0LJrqiVHl4a5p8mG9mxYG9zb/vtuzkHKY0Ei6RwmASkYY3OSCmnv8DWLsj4fKqt4x446l
7okPtE4CIuUkXxArAjiawxyx7qWzfqA20QCefjyxeNV0AdjPxEURfDWe/7sTGcRaXgdxbvWQzCVw
7H5x0mMoE5cgPXJ8oci2DIJnIgcFPDDW0t5wpgbbOoOLHhwjJVBM6E+ef6AEIxSHf7jDBmUT/QRN
mv6688qQx/JWXApDScem5L9PTl2LTsPovF4H+j6veSTUl4apxUNUlpZ+IIYnGF0D1jiD71vhelmX
a+dXLnRX4TY+u6BTwJVCiBXneSlBM/aKfqnKjRUFJyiWm2WVLNixQllZEFvFBWSf21QFA/xzsl9r
9cgzzRmg9XWaXxwerErFIMKiFk1GbYxtw+u7Vzy5TlMdbLQ4Rbi1rgjLBdAL2YkibcQksIHsbiGI
mTVrAaHWvJ208LjwJ1uB66rWTgDuk8Ps2bdSqmqbCpllKWqzaUQtqa/IZYGAdhFQQ57K8POSnLHX
pVNEC5sSjqYRg8SgPYEj50b2JRE/2RIEJdrwBR9bfRX7Ld3pSHnoLQF1n+WjcbLkNUIyG/abxKAk
plZdkXlH6XYr4jRPnFyuro9rrRMU5/hq1VEP8PBwabphPcGjqPY+tpX9FdWB90FU+nVlK8tiQblD
qQYlB4ip4VUu4wxDfwG8F+w9WYbLbem3tE70sNL5IICMpD0noc383ebvuIDhB9pkA95qiQz+cAYE
YzIOe5VVQlETPyW6jTJCFmJY/eR9W3db6qqkArQWSNWkRPt+D77kjgq9qGMZ5owgnbZdn7VYp6IJ
GCu4nD15xe9rFw/lRLaiUMviujEs6HSMVxHJ/SL87nUbt8Ux4FaFtdveI/CXzYSSvOIvGEtjI+Vr
PiImwyml9zQYtYyvgZyADdOHST8SB1dH3CTh+vx0wP3m+n9VJA97Vr+qWZoZ+A98d0ZO5ba41OA0
ZrX8zu6lFfVH9/w+mKicZxuNUYTkM4O69tXlYAfvtEQveOzWLkx8asDHJnuyFakVM5CSaW0CJUe1
aQTMe6je6BPiCieCZ3wqbA12Ni08LmBbOV6+QhN1Rz6bLO/kytVGUjNGejrENcYCcNIq5RXDAwVw
rdZyolhRbI7KfC56Mrfh6uNV4Z7ak9a1jHg7hTIYZNob6WpDBld7AJtaRcLqjDsuzZP2+6Qo9K1E
06v2jVS0dO+XEdNg0PVWbSpJaUfXo7Y2ylQljbBKW8DBe+Yrl/lslsGYYvnM6tKiASBFvI1urgHs
bOkQbAqjCVAaNcpndeBxiErdtBcgHARhb7PVGGjUekWBRilh84ItsGTHILI7otZS52+g53QKF30c
ETigQMdCCmzG9tEMOKns8RBoWpCe5bPTK4J+qG/kjBnhry+2iEvXzsEKymyADeYLkARahNlBbXpp
A3mSKDM5WIZrCokYx5w6E2DnAAAYinWC23dl+e3iLHt/qRDeE5ojCLShXBBH75/OtRD1HOLvrNmJ
D8RIzm2vU58fjeCbfJIi5N6JeeMxjvQQIOU3RpxR6DKndW/8oMl5CxPbXUQJE9OVGjaDVoNGgSwi
nX0d+oZBsFiHcLqnYBUGbQKgUlQyyu9R59YVMCl9Q/xOax0nU+jvc1WhjGx/wAdkctAIfpysvjF+
IxppnKm83o/2pXgbvRWBSn1C1gwBj9sPzV+UEe5rh9n1bZBS9ioOXNufcOHII1sFpaSxy3EoGXRF
WfoZvg+6GDoCtt7zpx502qBRo80KcJ6tbhK3XwEj0XgE/jZDYKj3YBx0tSS0Ux3TIONCQt6PDiRE
ajvDE/1QgGj7Uydj6wgSZ1dcv+pWMfKThqFkNUDaghniOVl+OJeS1Si1GCsN5ISowvBQ6Yr8CHky
xxZcMC4rTHHg8wJN8E2E1P3v71e7vV2/2cZidpm0ntbs4c6qZPDa2vRQuaoeyzlt0Tr2bHrkvhqV
4azv40UcBXCIaTRYmHjAHqxyvKGiyhs9GCo7rvsawpk58Oh+daR0QrMB/qzu4tK2tK2jzvU7xUTH
6u2RptwL2dre4C935K2M6ErGo64teQdBqKMu6QJHDmUUjtUU/XtNLYPqYQ8Re+5Qihi9SUXWPbvj
BItpQ9u/TWnOMKbzly1vRmEx/sy7qq5AZU5CRKecx1jEXIm9B9nL8II4r6nMjtUodmpCofcI3ymC
gpymUqJd7qYwFn1BWO+2JMGU2yyZ1FBIdQDjFlgNuobVOO037n36fOyLHD6g/5Jj/2hdtbaqL1zk
WLYtvgiZsSFkG9VDt6Hifoz8uG9Q5goS6rZ+JGF5+XblEorLNidN6dHLxkqAfcwHrC/HwSlbQuPu
zy6u7bMY7//JJT3okUDjNGW/5pl6pu7kn29iYCpHt4fDJRJN93jYLP0OX/0ZZuHAPhMO37GnF4il
2kOcgQ/re8qo+tQDSAYIAiHHTuxIl6X9HD6ukZSC7KWtjwbVQJsFqYG8nZ7tubITfk353H0qS+bM
+EdXBDwgMATBd4mpRJ7IbGEK8tpJrluF7T9wD9dNjpLvSG39XeU4nvi9HrrT8VyOuZLaJdBc2mUx
rsac7+whfR74jTL07gsJJcP4RAOPQF0Zd1pzwJ9wkck/kFFyIakx3eD928/yG8DE4Uw0b9ZirgUU
3otuyjzuDnBXAvdIOMcytTIGKBhbqQgpkmEuNs8cGdYRydjq1Kv2pewMj4O6QtSFiX17KG20yK0q
dkUxYzUaKO7xVGyjvyP3U1/OulFlE5SvQJa86hrkDnm6ZljvnmqiuhWs8584DPxHqYfgDxq8hkyq
tlDQm3vlXn6nytqHByNwbQQSK/U2xgW+aLYmEFq7PB7+qXi9ZsFXhSQ08v1YmuizipZrlejjgUI1
9DCZVGqz+zimHaiOW2qTB/kllarpojtgAz0D9eZQa0AzZCG3vYq/9PnIO4vt5Fzan1Emnb3HumbJ
S6XLX1qJ82TLmkqR0CcgR04TV19plPwdMMXqIghedRZEEE7HMxjMfg88LPmL2O6SKjHUC8mnkg0U
V6ExCWx9Nb3xLrns2itdSADmQ092XL0OTd6uSAv+iZG7KZ/4/58imOeOXvn/TOKqU65aRo1Z5BIl
7tV8uuwndwkxatoFv7XnFfWRG/9i5b2jXyTc1XZv1cnJ+PpuTlVggYw3LSujPZLTVHyHZ7ZvTCoK
NDfk/+MYfNe58br/jVgCaPTsBkvvQ6Rkz3kRxRWzivYlAdeQGfvJUSxIzZKICsgKl8eaUXjqrsb7
bi/HKdHZOIweLIJtMcaZ6lANkeorRK+R3oVitHuUtVIFoqB0R5xWYoL5/eVU9U7Ma0f1cjTMZqVp
spZpT4OuKYn+To3pR9PnIdftMyX/O57VPfSn64wRUdBK3rwgtFzLKYUQXHyhXKEx7y9h+wZK5sfL
wRkG8Bw3jH5A3Fa9/vtQQHre3ceMBDNRiB1xyAgSmiP55evEkrpCFpJaw/KLOrsm98TA8wvtO73q
5hL4QW2+7o0PUEvt61E1X8CyQ98apOdF01bcTn0xdobmAGh7/gclsVMATRa6f4bT5815A5RIjYEX
Bhvq7+STmd60eduADQYbGrq53MfljrCeX8LuC1X7/1Dz1b9How3/5vIl03UHpV0W+dk1vIHJGd2+
lMs9c0moeRuThFzEdiPG9pfjz49wcxKf/vUj6/kVQMcQHL/rqGYOA/UImZAarjDKT9CK7OkJnwTK
fZdnrZ+zbBPsGCpypp9LuFTi7M5TOGd6VrWUn19hbKUXv5mXA9sJ7wxAKN1n29wSxZBbGv/lJIsc
i6wqN1vYxHutAbo4si6VaeiN1Kf8cz59fX5ytgS/6y24zclf5PcDO+pzqiPleHpwoZ088LQrMr/d
FTFrNgTiZ4P/qQejfR9vswQ6dqPt6UuE/ouHgX8GV9kO4UhyJVtw3R53ajj8vha/QdqHcXQX6f1y
nQEysfu3+2crI/gpl6mbhfsM6cRiYG4HP7jv5JEquM/5BilVIyG0rcEPikqS/L3nUUL2NARl7t1m
yIQYC8Tv8EikHRyLn6/z1z5zWoZFSzi5Kti4m4nRmufdzv5asJDkKvDZWGve1cxDGi8X2nR6jh5y
YVZT0z/ZzocyC6co8XjmffFIZpwGtmHG0VHKSYLqWI3Jw72jE1b33rymwg0oGuzdDROBdQP2XSfr
LOc66AuzXr7GIsmZK8yIfBRkQ5Mz3ydfBSh/8NY5LbHxFBpYFasj82JpA6iOggjxGZaflRh6wQyy
+YZ2U+CEAFy9+PCuPX1t/UZqRHgw3gHDRo40tMlVXMgcPquBd1Q2b/ZaXoPxfzIxy8otpXjnN96e
ZySAUy45nVHAi39jhZB3eq5lTKPpRD+3Ap8Mm1ZG+7aUY2buF8GlPueRU01q+k8mErQW0uYTEPyn
0hxhrFa/Tp6zNxjXERIjAi2iPuA0catLg7Pb7R5BDl70IwRoShqUluxXXMwCS0SPJtQS94pTNhxK
kzLJ+MJfu2B8iYN3qwJYmNsF2bjokO/Qioc2HQOGHecJdtXg7BdID8Yp7QlSwE3oXI5MSBoHKKr6
3le3lIa4S3Mv9RdkRcYOJME/eNIveyyOpZjzHFr87wKqSjxMULghbFbJcRHt8yYIczzaYhmVukDU
+X4ea+8++AuC9zB0CoT5FL561gqFoPRA3CwnrRtnhpOjW5J8M9BE209lgT6hwRV5O94jR0DDGmw0
wIy+wh2/DMxP9cuJrYZG0yUf8AFAjTJzgBrghdTZgFkwtBYsMnjYswqDUbixiw3HgAGYIo5sL104
lSlx2GlOlhpjOBfBL+ehObVo9/bwIhXz+LxLSBU0Fuh44LWn7yw3fEl0nJrJIM9RJx1fxiNMTqt0
QF+IPKKRIAJckMiBkvLXR/7xTohgLn+DEW/qCJKiFzymz/rJo4sY9IDl+z+3AA6ANQ6uiuPbSbby
YtSnAQvVuRoL5vic4rwO3CBAjVkjpi+iWf3IUeZmG139P+ntoOHFKmuI7W1eWF4M4mVpd8dTEKnF
X38cN6ayx02QHEblhmbfNFvsn/HN+JH92ukWRkRPrUYeDbqK6xYbHYG+HBDsf05y7HMzIUNbgabv
1DWiLV2VylBfYg1/BL1gpM7haLzCzwwqHDRc+cXkjn21kRFk4+65xW4h6IPtQl3CV9oKOfO8Dv79
hK0/ckABN+4WuDpm8bQ48lzuyMWbLtBcRs/5OQ9F7YVNv0zRNNfnCtHjHGrAsd4uRgUmAVFFDkwi
wnqlBbDVuaSMt/Owd1DZXro2taTp/kGor+NdSf1cvPhpDzPAssWkDeiYKm4X6zphAfgE6BgIcu12
78rZZdCpPze7dm14Fbdk3MRM4KwHI57rB4f7W5oIlwDs1f5pAdixUAgISLkwJE2F6nG0xjlGsVEv
vq38aiJ7psWfSlqzTZAzHYsbO+4xD1GLp/V1nL69SGjY2VWh07WjUa0HdWNixHKhkycm+McOU2Dy
YbfDdeB0OktDsuJrfboSOIcNGL+STUxX8+tjYpZEytDcoZqnkUN40FJOlfvgtx41GmFu6IVi6ry3
HfMUrms1ZTJy3mjg9qTH+Wp0yw9BfG1niprJdWQjgtiXJqjbZYRir5p5O5D7C3cHzZr0uKm1TUii
Ux3C0qbsgJb/4iJejqHIYoUCgCFPIE/x7Y1tPhhpdiVfutoBpFLPc1UOH6Pq8bFhLy0PRrjzWi4F
3BkK/ZgHL50P04yicAw3wvphR9kCm2+pFrM4cjbf20ShT4S62HE2/5BpNoItJaGUmh3elHcnEb8W
hJXtaQ9D8TUuHjz4eYNB7Hu2NaydjaueAszREnMdl0KcahyI1hJoalFKB3nu2v01tjk/tP2uCY0x
yfxFY4KTOGZ4WcK9w1K958+dn1dNNtA/4Fo9Udob8/U2ycqCrMkExA+cJQgKEzYfQCnUTbbcTWK+
Ym0CNNNvStnqvvmzy5bMYcwke2Jxso7Rx1BsgsGfEwSK+Izw5hWle0mgWCwvZoli4PRBtl6hVWhA
Q1IUR//Sh7Qf+QuZnQ/EFuRZ+Dx5je1EM6WSdNUHOmv8SXS7AvLdOAmSj9wulvFrmJ0o7UCLhyiq
GnqNm4SuyV0L12GHMXO6C5WGu9tGwBItSwSe7cr/nd/JbewSufiX9dxF32LRpddlnXeRlDIgTkrM
nETyCRxb9Nsg5yFTTYa3qutgu449qfsIjzdQoU9KcmhWgSZjTjNo/UdJSv27giKLfNqQPLACXdMN
MHDZ+lGelZ3jOZqKodZ2+VW6UMRvB/hN7FsBeFWrV5n/CeYvspc59LjNrhXawQ8wsLv6NL1rbnwM
NTuJ/Il4eDwWIZKExulllDYHseq55ITEv4zfw0Yu5McdcQcNSKRjCuCLf55sllQ33hWsyBnAIlmb
kQ3jFel5qzDlmdTSLrV1F0LhQ6OboqSsOjmbOdCFjvriOqet2B1hDG2D0qhe79N59BawLpCvmxe6
gFRChKCc+azk2fKwHvLkN3gOWxy8X3U2Ax5P7EFXlj6jUSHuqDjB/Y8bsuE8fUIqt97h44giv97n
2VbbxLP5AO5N8LyEqrGswAUtc05JYtmo8u+/ypGZF2ySg9ZHT1RiIQP6woObDzcHbRki/nLRuOKq
v8VXj09yadOdcHGJ9TQbh5W0noJ/IGBPfx54f71+Hm5q7yENM49u5ExbstC8mCakr1/kAMHV8ACN
19yHmIDZdN12QBnbpYCilaoDy8OIlhW4Lc1dbcxWsWyv+d1z4wTNv7/juKAMSdHz7hstJtvxN7/C
YQbi8m6cpxeArz1EUN68HXGuJclbfXxf3O7gAMEszrcK9MTnsHgjjJnbzu+a3BFJwizNp2VfVMMn
ldxONXyOeykQcAQiMgNHKlWHQQN/ljqoqPxYqSoRf/91rRP1uG2X6NrgxHpGyBDJ+/1XcmF8b0Yq
fXbievEmN25JuVEjqSv/C5xg339+wKwi3Lr0j3TNZFVzoMI4QR8TF177rQuZrPJsGjbYxdM72yhB
0Y7cEhoZrukkrAkjiVF3ZO6aeo3Jlh2ffifMwLlltNywqQzBq2+YRyy3a/AyiEMP6/k5CxEhNb0W
j7mWpPW2Cg5Gjyqg7iXaYQIEsA9kTGVbmOGPiHcqGmHBJ66iiNbtppjf8US9SJ7eylG4435oHpxE
a7+mHJKVHvPWbXudMsM5d7jZsnz35suM6vpdahFZ7XLyiEzxGXxUfi3gMjACp5QoUd6jwQOH4fnY
kGzYRYbQQ4h4XRwkddBvNki/Flf9l4uB3G+5asd+Ril9ZPumaoxHITiVRDHPJXgnP2aHHT90a0Bs
kSl912pQV/ma+Akk2WSw/sUCIXnR/VX3DXkC0Xsu6YAZbH9kIQdxfuOKrRhbRcnEfPsr5OwdzDba
lCsd19/Sv1ZW+R74nlLXCUnQLGTtmvMHKMBAFKt8HjNZDO1yv/qfF14SosRIuXa9ymKYI3Ed4kug
ez2yoWC3pEKgk1qDjB3x8c40NZkRcm6DSCVNE/BhoTonoyNy1vygoLzAE+gcJ3xOPX/jKK4Grbql
Iy/4EGrFshadODX+L1nAfy3s1YF7p1GmhrSHa+WRTYGrBh1IzNrffnJtiu0LfjteEhJoJHcDU4j+
wvjtjsW+qKX+8WvNRfKu8pPBM6TpE48Q1fjd0y8Nl3A1c62lN0449S/Ael1m1Ip/gNauk5SSSTpd
opQRRN/KCfDWLG0YZOWA4uXo4k/ENpDCh2UVl9TxTKhsOup+4nJefyf2cVQP1Vjq1Y48VIh4d9RK
hEPmPrfYVe86aw8qEq+V10Uf7cpIGIkV3XluDzQ7ZHmRuv+cFuhfemFpn/l5QN7dMmDa0d9fI1xH
tvgJkDno3KG+Hf+SZ6wo5/I3YRi17K/0g+HoerkqHt3YmTyPzy7g+3DZwy8lm+2yE8MO2GN8abPP
g1vfoQxhi6JxnDqHfNxHPrgWiF0y3vlCcNdYdSmMauaXJJy3LJckKqp8fL/gHwHhAxNOSPKeCOgg
XSWoIsDHQ7aKJGYYpmdw33LqnPl3u0+wXOCb5wELtj98qxkq/uvKvejskKgoP4BG6jhQsmYA4AL0
VT20/up0/RJNOOuyOHInXbQWmr+NdR6SkMX7jKrzRW1fWoDFKpMOwO8h4CbWdWIeeF4g7pliXFq8
1Wt7yx0unpw5Yfu6Gm4Vqj+ExRZhJSzeYKYsSxcyWJYkC/KUYolywUwfBZxNhXWd2zn1342mhyve
V0zKffk9mztx3Z8npRmatVkWEWHofs/CrVlrUBeWynHwJb7IxkgyOnqif9GArxO4xguvkMG92YJ/
sZ50UtfosSYPakqea+TrvR7I3Ee/TCzfkqIM9feIsrkaaqEbhVlwoTf6D+gOD9kx9mu2t/VyvhsE
NbE26Ca7PfwLmb/gecNmWPdXF5eNWDdetifmmO+toQraOtTeyqyxbLjmuf+8yHRYgdccgq4xYumy
F4VszPO12Iq5dV4PhgFgCWJT1c4BUUF8+cjIPPx/YGZXOf3Ej1kuP0y79jsR5mRXNd3SvEWzN/0r
EwvsGZVl5P1sAkfri8WTcOoq6pgc4CurM5/JrUaeWyKaFKEVoXsGIPipp3iYrdy52X6GsdZ1otwx
dgaRPZMnW3La//H6zXxIiPBKQ0mtmWuMmr/t1sAl4hI0d/ExAcRWDJYISLzEu950NGyPcfXEJmhl
+ccFovIrjYcAjDjCtmeY8eWeyNNU1FVxkOMfS4YkAhCvih+6N6wvRZMNx3KruyECngnVAD8RGdB0
U0rF6y3kRX7jOTOJrqntYaTbmgdwqt9x129gozFelegVlzGepExB/ybFxeaBShdWr8KT8jSnAORC
OlwRmCeB3d0aolDmDqqmzd7TzU+UMARAFkvNza6gRszvlo6H0puLK4r5JMOnyignEES0pG+Hnjtc
KgA7oDBPXpcT17r+7pQxFAXhuOBE6lQQwhfQEnA8Nea0vFiV3CpufW6OXnhZ1yJyK2p7is4Rg7A4
4MWE/gxrNp49TsHVXYd28rix0Drd/m0eSE9td0/oGGxywBk3xFwK+WasPk25Od1XPxjvHknYOdYY
+pXpyD5UAEm3gcm/OaXH26uzzlAFHRZbJ9UoCeCMeqbdlD6QWGDGpW1LVo7eqTzanocWnZmJsXFC
NYT0/PKAbavCF7GfmlMBQY6qt2Xvq4Qu+1tm17QEprt5iW3MAo+OxYoOESgJiLDn7o0zX5X0Gl/I
d4I8GnXkQ+fvX2xc/1+yY94UGqgLz/UZ5LJxrJgDSIK0I31xsQ/j/eNoyK1ijAvIhLibHE8FHUvT
UZT7y9ajQrCI84yFj/s3eBtqMgHAtY1+jtK9IvrHFfDQepOs+sPKOI6cxmhvZD8c+hVwmALlT6ce
2jKZ9E8hqUjKEofu3dCTMBTFwjNjs3pWO2GKlC8JIiQ2T138bagl2FVaFx7romQ3VuaHBtbAuW0g
qZ5+wNMJXt7QDBB/D1H01CI1GqvIKhwS6sTuwV0EOzdwMjb04RQPO50gRkfuF+OVAlo6Tm5EZDG1
FMJzItgADS/lNBqE0AGSOL4pk7sPP26Xi6CUA5Iqr7yGFQIhUcSsanbJPpTMTw3y0jTopIWK09PA
v7tzS81lbR1UdFEv/fkUhtWNGPn71TMZnKaLLydMtYmOE+o5/7cMrsGlckPHWGqT6McDgcy2FHZb
g2/YavYE+tFKv9qL1gT1ucLGSKYcvKEMAls7hErlHj6g2pjdH3HKM7K899B24uOta1x5Py9q65Nx
Tg0lCNVHv7vYqIaBaYggNRj5dwl9g40Zt9P3au7WxYBu8reCw59F4/o1iQFPdDvCzDXaqmHRQofs
4fak26CFBhKHeZVnOmGhxk//xi2UpjNBplSio4pE5QUasYHL0PL3UumswjYpF0HX7OGAxuFWLPdy
3e0feHsGWrYo+GeuFR7txamxx0584yfbPoRnMxzvJlExnRS8hnP/y4+0SmRk0zhEDwyyv79soWm0
oB23HtA92wN2Ej2Bdz6pjfg4XoWceueJl8WyysCpEwfe5sjA7oIxTu4t/DdrvpX+1bURG0PrGOl6
9XAduFWdc44DBiyBSn79POGtZczYlxbfnOR5qJXvbrDY8Gm+2bSPL7QGtHdiY2g7Y5MWTyMdkeGe
pE/B9aApT4oUtxfU3PH0460cm3xge9P9Z5BXKIym2kbEqH/UO/vGWgaogAApsBTmM8CsqEyCKQSv
iIt7F2LuEVs569nAJSbJj7Jd84nRgEddeHSf7T+xpY6HS/Q3AtUvZneK8H5/nrLKT39m2FcFxRoy
lIdaUyWlgWxKZlBFkvbu7TNCghmBO+1+lTDNpWQzH9RcX0BcRfjbRqx3Grxn9pMzc9mji+O6lnzW
EZuLYUqT8U69LqcvEDB+bUKHI8L6pYjENRpGdp4etICyZLzGm65Kq4SMZB6kYzxwbl7enhOHArWm
nDPwOGvEdfi3qdxgBFZi4wQlBrqLK0UsHVbQTAPpeK4fWKBshCyXX24TwL4/4nouUVKX/35fse9v
z0JN0eSvPEyDXog0yOhcZqMpOombSrxqH92wR0iBDowgHzCzNXnzmskW5NSJbjHYI66U0+JflKIN
UAR51P6IByyvziEr+VqgefblSaK0DmK7kPicYaKpynergqwHjiKitiGnvbcJnNNpaNCMWINS+fOt
xlHP3sXzboRe8XqW9TQr+ToT9wVLcI3xynFUuFg2ECZioY8C8osm9XuMfs9JouhSpMQbTt65cLQ8
FXKvcfs7Blbu1tXEbgR3AiRtm80ilke3EG+jbgpwYlbeOtkXI9aL1+zfp4rFHpPw0bicnFRcbgW4
QOOSmKkPlVaeuCO8iXPOyX7qJoQAVVeezuJ4f7hqczCcC64yV3SyB5aSkM0MaqfQLB9bxiw4M6So
55xA+ziQGWeJC/IxvB/y5NWcYviMs2iJxSO8fRakrfpR/cZifTz0OAqaPav5kcBaFMZGdzSaE3uP
aNOP3KbYS94vK9mL6Q/g1lN91Ky/9KdjqnkKgS76gBO6Mb6o5WcFOCEcN3405ydIdzUHd5LGtXyV
9VkPWBUksRmCkbTds1KZ7jdc5iLvP+lvTtgLYv/FvxJaC/n22xc5PUb3p6VdddvaRE4PIAe5yFfp
2XlovVW26oIooCTs1hUHEzdC5ZrjMEfSUSLx8+RgA+sY8fjt3JifyUGpggyP5mOH5SrCDXyA6ZyT
NjL8e5QsB0me22FdatqokWa9FTVc96mVTtrhY8dKPBV+U445xshWwsiFsmw5qtNYuDr5tJDxG+57
jH5V1xrwV3CqmouYVBQOSMlOtruhR0K2P1Stdst14/ZXt66oWP3AzAICuUQIRlbLsja8mx7YywxS
ye8bFpNu+UwOX9RbRe9TVRwlCyXASKHT95ibK3MDKusRHvv9Ttzjhg3XmRCP3h+wNhcUjLb2Flwu
VqbnR5VrLY6VcwwioenWDmUcauuZLgcEZdMGQRSToEaGmvfyDFuwaSxdrntqJ0zdI7jp6yhwkR+G
mjS2Dr0lh3iUtN80F431wiHWaFGDUHSWQbxmJhF0mAgbVVS898rR6STl6ifSubuX+JHogUa0Ue6d
2+K3uuquI5Oj3NMSBT0A1lOP9iKlJmktRFI0DIpgsrBdKlXRLCMIx4+GEEIiaA+nfil8VgxsrMBa
pB7jZQtCoWXa8u4BKGSwPyB/2yT8J1k3IJseV3Pz91NY28z3BgotxI8v/+ScHwXidNGIXXpNdp3u
6sEVJ8aKtnlJSIWWCMne1bugvHafBh5XV+mgqtn1cdJlgXn8vPTCHn/CWDfl6WG0ysRHHqxYDbrj
zTHBWWy/RnsEF6VRfUChLvG6/17EQskf/b2W33XMy0Kw2Tgbqhd3X6zFa7z64wB92wOX+LeTgv1b
0zGgZzs0GCZsBP2ZRc/2F1CzJIPWJpLBEpB+Ls+WGsQ0jZAy0PSgfi/ba7GNYjQJYKylO0o1FzXs
XVgk0tQM5UFXKf5ekhkFza1isFlCFgQ88vIQa36LmmWc+VWM2E/+LrEZxaMCaGntKkYkyHYJVV+l
PUrqtJ1cLgnyJoRFh4pNZt7zhpaBRUq0b28PfwgBRHKlNAKmcNjlZFTPeueX419t9P59QkmqwpPf
syb5FW1vQDwQCBb2O3FFLwks5wD8NN1dcLMqwUBq6++U/ho6UxyqVJk6K/mF3+s2nqE4y8XFLgIy
TLduvCsruVq5fg0N8EqaZ3S8UirKUy1ETG6s9V5o/4YMunVH+RXwOnlZue6We8HF1+wu7TW8XnAu
9FA4wrBw5TZkjR1TCkth0E6TbcIU2v/euqbO1uU+4ZX9kPCAx5IlfTMyQFoJV9t1t/po5SJ574XL
9BvId7Oywdew0GsxHlGu2KA4uWtjgvb4JoF8RD8jexYg3eOkt2eJZ3/UyYWL22R0I6WiCoOobLmG
bflwukHiVWLFLSMb1CkhXTJliI5nlRTc3l5VFLcHHL+Dnt+tpU4hjuGTaNOm5RPHTwIxBC9iqcY9
qbdyktU+x7U+erjo72ioRBSKRoThPx9Vn4fanXWi01ms6AOAFAL8MwBkDQoC2cn4TYI0CRLpJcSa
gVavIXJqFCRR1l5EIXp0CnBqP3vlURaKfOyOHUng89G/p6GyifvKGzOCl+acgHn6AQujB58sZYhC
HbqdFccAJbq3LlY8KH1+DcqKGLuLxaHKoAEUMtX/e/CzAai8HKnptHZq4sS0KSVim6hJlkfOIaA+
U+Gzk0TFqJF7po29betGNJ2M/lVnF1xlBkI/3KsVKMG4Cmed8PY69TDJGOdVuGTU2jwWbvoKHIxQ
EHNw0OuSoPE6JPfYB6T/7fm8mpicuBCDiMtME4h8HVgveIDTpTR2l8TxQmBvW2LxEUJBac8CxpyZ
D9jsjsi4n6F4AqugAYJ0mpF4F/KPvGzOPhhEcH++0kCR46snL/qiIxgqMkW8KlVauslJuhzefj6L
wQBm8q+WykHYpyFj82UFAGUkOsvmNBzqRuCPtpIHCiVvLh5cdTfJV8U2xNlOKVBfH//ShepIHQyq
vzkA6eI0K1s5tSLXkx1z6rv9ytmPaI/DG77La6cVj3EFZc7sZoYpOwJonMsbNILuzhzqBU7Mmlzo
b1ab32o+xQ8/z6UsTqrhYW1JCIq4EJiI1xvVAnK7cg5AsRTMSDGjCQQ65NT0beK8wcO7HiTtrgbf
zTDDfueITyviJl2NPmdc0vNz2pDa/MiSb3p2TBQ/jNDejVlTRtAeJo/ow6HOCHk5YOOO/Ub/lCMD
EPcCMfsx1lLelpJPYXwPS9Ayfj6BUx75BY72J1i7gwuw0j9p7vzR1XODwt6rkMlZYIQJTBUPKm1/
bneT/5GuL0CZbNi6v33vHelJm4NVn5FW6iB7FioLOsmYIEF3XxUrn9hIEd31CNYEx3AN4X4qJbtf
pdcR1YCTi1ziWYD7qyqyGgmPX+Wj+7ugXP4fpgBdweE5kWoj7PRVJJzkkbInZN0HFDqqMP6paTbs
Npsclwu6zqbcQaLFovpGlrOz/4KZtlcOJ+fr64bUmXmhByZZTRrr0AasBWejkko4gSGw62STmOPg
VvbZt7yvWQLOycAtQCR7tHydalgOKNSCw8MBaupCB6bjy6jPmQbWKoEW2VC6E5b6HnuMLfuhLnZR
VB80ACvwFE7b9itcpnU2/75tmIDSDyCLikAP49Ynfu8Kt4OS1kAKqVmDkp8PtZP9bQFVomTrxaZX
Nvuu/EuKE3ROu0OETZeCzJ0ZwyBgzshSUbWGm30p8wM+5OjKweOAG46qA36fotgWB5DIwxLqP689
NDG0qkZX6oYrpNpBJZI9l6Qw571ea8uQ7odMr/4HEU87F700knXTYZWAIVA/AelEfp6hg8EnrT1Z
+TnDq6mKJb+AbICFfQvMb0pdS4J9VdsbhIu6vLpqxwDaBaKOFe+ziXszAgSdwtL+sVOZJpZDpvaV
cJy3U23w7hMh5+V6epwwb+xdRONbGyA5I8ammI7u4VgLb3Tid0Dxy2tHYnL+pPtqsFjg36/XdoFS
Te/3U5kLfF+8iULgCRHYWfmFRene+p2chWSO/52V4niOz2uiwWkMNcGrm4MLOH6tNMd16uybkXjd
xhqloNCtiRtEvW8NToPml4QOXJG0t0byU+bM4jGJX3mjcH0dTdPP1xrIXeKMcgTMdZt95q8EAQSC
G4LU2rIIqULAOVWc7FTMp+lmEg4tfxwRQjt22ySEZd3c/p0qCryVXQCPQiRWQ+mTyM2z9Jcq1KQK
3rUnWkW0oSVI0PpRV75EZl0Tuzn5ffZFlEMDNThCtbO/PMtOqxZ9DNDhBC0ogU/rNzTl9XY83ZXA
x0ZW3uXM0A73dkzdl4Dx4Ue7156l8PS6OsUULlxotJUnSPpR5weehkcKREoxvFrtK6DeehzCoje8
Y1CpImm4c6IkwFssviU2e7LYI+i5h2Y3i1dafOkHpQm6yjjNW6g4y8o3qFu7zJsodd3apA2adWwh
qHTUJgHpJoi3Fvgz+QVlLxAqx1FD5PEsgmi+AjIWsD7VqlY9JmYSVRU605DFrzQcjPrgeRQTv77x
E3USVllz1+ZufK8yB+fSSUtevEFSoWrdeCUM9rRgInFs6eQpOyT/rAT1GFjJA0ALyCfUGRSNkTFt
C0z0qXUUsuHtp9ZG2UBbJK4EavA+D4o95B47I+ZiGOeR2A+4dkE6h+/nKc5Z2T45y8ImTkvM5x91
EipSECX4ez5J2DUS1/rUIJLOFSA6V6Powor4g07Rj/gkUh3YVy7erLGEv3jl/nbAuwknqgBI1u00
K/YypqNPKn/LwRC+4+y3oV7GwSEwmV7xeJO+6PKrLOsgSzycgV8yxRsrQ36jcgGuvLMRxke1D3QG
v00Lg9Uv+7V2TAfd6Vc9EeH3AEE/fV3ThirhNcg+LQQgN9Cc6PPX5rt3BQoLZyPGIGy9oAr5oYM5
uDG7Uvf9kpZZtHX74MQO45wBvLDhXKG9xY6KcupJykKYDXM0kq7g2Y2mB+hvIaY3d0SRUxVcCvX2
g/iyhyom0CgaH9MKZYxTE7Nfx73h/P1R88V21qX1re12qXuGyaDWN6hLnRr/+NKkCeGF8b1SNToZ
SWLbKYojMjmvs/gEJL1acpjP8YDk1AJBcuU0DepfvKqHd44BbQDBjSq8Q/FH+83Q8l2oWNWoHtCa
7IE0IFanGrZu0N4nk8i7Z4ke21pDV2LrGa7/56UlxvwLRi75JOjnwc/QFMt1WJP04dDlmfUG2IXf
GntETziAbAiD0o/5azQZ0U57CHA/qMEeM+SmpVDH1x59WGJ+5AvKATYIbcuol05y6Il/pj8s01Mo
EHPHN1PKE0rd6t7HgdIfwKazMqOrUjDdQAPI6X5I+pL6oLNpz7QWlwRg3OZH9ypnw2LD83J/gCur
2P2nJ15coBb+CIkqIT8vWZVT/zEbB9/Wi8YssTM4WygdHoeMFfiVqsd2MrOfjSMQ43qmpWsAjIEQ
IZdbydoUyU8elCQrNJ2Xs9o4QosCSVd8nvNwyQMr26SqxzL6/gNvh21YlxqfHIUP79bny6O+3khM
qpxeYsn12nVzn+gi04w3HPRktTYrNiuhjMz3Yhrc16GrjofHgVa/KxjNf8Xb6AnAWWuSUCEUNBFN
Z2uzFrHG5VuI7qdMNdyD0ILoFI/dBEJihGNTSEWzTUiQ73Oug+YqW3C0+nsuQfCQ4z0jeUIUMvsa
ALjcG9eancmLPXd54JPEKtZK4I4vxIGhL/wdfGkgIV2KL2jiJzeg8L0RlybgXoxg3OnjytvoUHCF
KXqd81j3+17Clp6AXws7yqTsf/dcL/gCB4W8r/Fz1EQvJ2zDtTC6AWTSFeRagk3YM7tKEn6KjwKk
GbKk9WbnnT9v/5EOTL96acOvDL1HC5kP5GEwhVeFtObsXb/aj6ExQPFWY63aSCj3Wm8aMyg3TDKM
WQGKk7xFug+wuKWmwzpxR8h9wWruh3sZvXdT+J3KKy1138syxtTTaR1qBA6d30581sNxC7tm9NO5
VCoYMeEl9GEEeVWgXznnBX+EuKA8CgpSIxTrg9Q/gl0iZ73cyG2u0PaUQ6eSTAyLT7lPm05w2+XW
40mWd4hBV53mrMK/YRgzcBlCyXyTZDCM6nULwBIddfVCZ69wC7eZXrfcCbISHPUE9DnBLPsnzDt4
b1bJ7/lehM64tnAgeuok8pZf8qQo1KasJftUL+3b+RH7h6QaTrN99B0hZ7fyG/o/DqFPe/wVaEtN
k4N6V4XAOAxGKOTSix1vFJo+sOSk32X1ZyDNxcThNFrCMZd9Av0SP/MSEFrdrPS686ZCI1HXYRvv
MjI2ooV5Bmc7DD6eD7BZxi/C3wyAzv4ZmmS4AslIz9dE5KdAZU/SX/lLIi7u2l+kHjg4dHjTJ5qx
M/uB9xYUbXLTYMXxJiT4sAsHf7OBNzGakepQG7Fs6d+3fIbKhbJzBNi30CJatRSltV+SaZO+fGzt
AfSfEOnRetYp3mQTf/0lGYxIt+eR7k1yta1DscFJuV+qMyplx63AVcXrTqNAsKZdGAxDT4e5YBNN
517W1GxmS4SZ6JV8c8v3/Q9MsFv9Ay4iUaL8NCRk+w1sVjU5YwKETOkZ8NB8xihNNzqyY8/2D1IP
Eww23Yj1UhbNQahfVmxNVXPXc137rpAJAH4aOeyDPzVe2Uv04V6IW5lw7dzEdfq7ZgBbBcbylAuC
vchsa7T3L/SqstyaMsw452YAVXwr+h6ny3/3OqrsyZHmv7PL3seVumQ+G9FH+At3nc6CftCLnMLR
tGksWOpAhkJh7pr9+g8K27ZMZgXu2nKRghktO5YBBG5vig8etlhtTg4YRb7al8Hd3hOnoszLKce4
vos6D/mSEEKYoo6wOmq5HthZ5PSNt/B3MiNIk5cKb+6q9SKvYzSicL0AGAJiT79a1u5srCII98Mg
NswOFGEO4UHdwTf0yB/9p6Iq/FcDgsar3oZhw5sUvVIyJVTNZW5xQ6HJlygWVaA3/bRb8Nr+MP0y
psGhsP4ymB49oAPQk7xw+1Y/Euu/2BimZI+Ti+luJRTLKhWP5oGsvBEYRPUJN2VFhwZ1BrDAnHb6
GsFqkwenMjUzaWVw/VrMJbwGxgPRkNNm0lcnI7i6l8Tjmf6/ZcITFtxHgJcYk/Zc2FNPqxUAbgy6
OMHPTjA1cNuHHBp8b1TpsYvlcSG3yyudW8d03ASBgWe8u64Snb0t19PJDdfTunC8gyZQUftnVhsG
/GmJAE9WXjC1jn/U1R3ib0FVZsbuk3x5fsxj4rmfIB4P1+YGhiJQ4bmyQpwwRbck2+kCpXP3f+cl
o5LRlHOyj82FgmVGYTccLIK7bwtCmGvSEPxfCqM4U0gqZNMV0XCBfmVY0+LmX/qOA4mz3Xa6Z9/y
PpwAJguR6saBKaaGs3yppQQegNywwLamCyjPMj//HiTNZKAWuGzmKazQx+kes52/LhZ/9YVndBuU
5T2gm0kDE3p+iUIxGQgB2QnvUzglTCM0FABqNJpsxaao4yRasLVNOqhetO9XaUWYuQnSNEmcTDMK
byl7iE9y5Xi3+qAI9BiIZZkBkTSZ039HmpsQVYyHfgbUibcFyQj/GrFwLmGcTlo3zJrhNI2LtsU/
vt4IUlKvB+ub7c75YDYa0weS5yUIQ3TWwTfHUvWx3DaFrUpmi4EyuVcsdaUrUVF2FYjU3zmv6Th+
6lKoVMAFomFQ2TsjB5zaemIu9J6rtpALiApXYdpC+aBEk+dj+rCQ+7Bt5rqgGppR0pXGu+txoiWN
Xm1qcEXTG1R8V8SmGA15l3liBg7D0FsUj2ZTuIUYqDYAGntnJ5k275Z4EapQgbKwWIZ5u8kJRwS7
aLODtFLMGHanwnnRbHDrAqhbdqWQpgei3B2wTYqJ0gqKn7HfbKTZdOJcYgigR6mQqC8TZk/fx/Ay
IuulCowJVdggfhmYR9DRx3DoQb4XabcEWC/KNQgyMgpSUre4NPyhTbFIT/RBsuagszQB0huUXZwy
b34WHmaoryUtvX+zSDhNp0o+1W4wA0ONtnSuo2UgWQdNXaeKVn5DVtK+rnxNS0JJh96dnbJPzP6h
wV6fJkCPecqujW66W7ieeWvZAxCaeAosBaI3FBMIRpjE1loyx08qLKQhBag2dYRljqswexqDpiZh
UEcvDHhVqqB6B9pmp6BH8m5ISFURrq2rZLEUT6KpJVn87BM4PKAsYOiiwiwX2J2YXTptWMx8zIyF
cdx1VrHURxMC9NbV/Nouf7/oCQjl9KFSNyTNqIxjDzyX4bznOManc1Xz9nGOXpP/C91mc77LN9YC
fo/YjXqUKvzsDHsJftotW7+8WrgwuR8xAtJBxzq5nQDPgYXljZD30pzJiwE6lc3CTIIRBu1k6PC7
N+zLWsboB3DMRKSuiU8nt/wxpO36sq7B5+DFD5CSbgJW7nGSvvJ4uJHkkqR9hQ8zCQruFuSJyuwT
bZUvvDxoKi5NpSB87gEVqD6vzfMIXrXfDqIT8QIPjuQX5lu0Akd6bfTnAyYcGQ6nYZ/YWPY9LpPq
yBHYNcak0Jl4Kp5qFImzjJAbk/PueRd0WoNyc9IKWYEg+Pn2G5O2b8fo/eps50/YP+nfrAj5Q/y1
tdxf6Uf/b1GjoN4CDnB/GyyKywwTMwhz621TWmOKIs7cepSgj09kh6YzZm4B6U4+1jTDvbgFAR5U
oMQbyfMhzl9TJs4Sifm4XLNiYgCcwYSf6tPl0DsWgQNj7cr42tmoGh5y59eBXnG2e24tgT+3YFv1
5hPDH7syy88wRYKB5LU116MYYdF1RPwZnVeDef/AhsksmInJO0XYtpWm+mrXyUaYxw6YnuABYcOb
TqaQGrXFBdi4+FL1AV80Mnth1P/vpv+aUmCsIilQc5PeS9UZkPy+q7v+inPhFILVHtrNtRbcmWrr
eRLYulG64PRqXlX96jK9Gxy70x/sWHHz1Oez+IAu1PazZywZx4YwRHAw+xCCtU90frmlVBX9Ku/X
gnuuUBmxGe2ZRsU1A8D1zpZ3BqbRRy2TiY8SOyjwQ+IEcbA9jJm9/+GKSKcYVj75KuTspoVqZzkC
5TEdQXWd25yG6Fko5WCxUDZrGk0Rsfv2gPfuqyeTF2VPFiWYZn/IMJ2u4fqB/aSCPX0pr4z4Htdr
m4IgNoAbgoMKSgsNkoVRMPYFsAVWyFX2zU4IFVHxhEpwyDJvUdUoRcxzPmZLY3HLVpkM89ZOQhO9
Suo8elmDtS47W+XQj8g1jXc3Y+3OHmS1exSOwWd+32v3+EAGlhVQ0ZQSQ3Jx2KpORv7A7WF3t7Mt
HSFiq7aCBGdT4wrvnFSnJK0Ck/LLyqLDOnWQ4zDboygyKdemfyd6XqQ+/nWWLiy/nBxu+QiqnrMr
vu1XtgmgIeP+E7+UXpDDR+5Jv3OLFy2TxnHA6s5+HVgS3OUZn1NlhiSwczsB4Dvi0vfCn6gYo+tQ
dcAUtBOLpRp2PWOVwxF1NI+tsqtky4PWiCBnLRsVduz+j4B1N8D+lIjHbQjkrIAoJZTiltBX/q+q
vZ46zvL/8QiMI4bu8FXydGA2ZpG/c/s2EkyGYx/v4oZz9GZIwfk67uoRH6zZrIdxQ0VzUTtEFtnT
WAMyoplmyjd19bvNWmkaovkvI+Ndn2yyO6LXOp971uqxgdhi6bxRZ4N43FPjmPCtkfEfiS5Z3LUv
lwn+/zQwEtGQtpHKYuYgoolClQ8fOR/nPrLuji/mLH2czv05Bx0y/BVuj8ZHgrN+38tbAd0I6zK3
stnEeBQVGIhhKNDSM5xd43NogGVE/3J34Xt0IJJwyZsSW2r3hBS5K7xYMHxYQI9IK087Pq8RcXFs
BB47VXt/80cIaOjh5TJ6GVVTsWBJWr41RkW3csUYfbM3gl03ODy3uuqwMPVRDX2MDi78c/vI9toY
iUsPm4H7a75PXkKbIj2tq6KYpZmuFIOlmMs8reaImXqoc15oQCqiRx7ZNHlnNisAY0b7NDPM65cr
21dpS+jpHwMlDsuQJtpWeHqrHAsWMm3pkm6Tfrh1jjW5rrYWS2XWuipPIyd8O2FNfIR9APKt70tl
pSKgltuEtfg6cdrKNBnb2pV+xirNJC5GJ6d9qW1HNF35nw7Tx57AqmTJ1zduUV1ORSk/BjMmBQpz
id8xPEwQY93O77Xc5oL6Es+c0PVQzTgfUSMjiINFdskdORZ3sLNJ7D4ZpnalUsl92jOAhQ9zTHk9
tg9wGgs7h9uCw0WJ/RtLR/yXwukkUIffr8bzXOm1AeiOBEgB7nXs+QEPzpXT7vGkP6mmnI+6xjZf
FNX/o01TR7lDZ2TdohHEqT25JnArwq00EH3rT9SIs16ot/rrDiuSzZU4YgyPyBAC93xY26uYyTRx
VnoPrscSGAy9kBYpVzJj1LFTrK2pW0+56mQFFfzOvsMBgXkavPLJDYVS8xkV/onZgVi4g7sCUizs
RAwwPKadVTqR2swY7QfmaeMdGrQDezmkfU6FOD5Iy6uc/BqHZ/JQd+p1rXRWc+8ns8zEY8nyYaJK
Z50GbJN42Zxp5I/Krh61AWrlD1BEbL7nUGZlrzFNIq+aEVAU/r3IOBHBEiledi5NOoENwkYnAbug
wakRCngABIsGKB7wshPEt7GrjIr4gB2EktOAEFiInfDi5PC3uYKrOgcFQbkEUKT35gRpEYvWbQE/
QoTg1jchdDZzqFWZgMjEgfcZqVKtKinA9PA5LLO73k5vlppqt38teiegUJGcNJk5pWDmobTCA8wJ
B8bHfpLnjsrOPb/f5519m7MZli1U+Nww6xijZbgvOGE14kPU8I4P6wUpr3XefoScpcbspuU3aUWl
1aO05M3VeIpSdLqColX3vC7+HOdpVyFjz4Iiofoc4ycG6jO+pk8wu9Iu2CWBbrxGJTVQqK4oQLBx
6sLjsjkkcGGN4Misd+j3X6awKC72zFgx4+SyYDF//ihmlFKdp7T4M+vw9U4rwvSa4zkYOW+EbjLF
dCubdOtTdTXgOC/1Nb3jk59svt1p5Ii2b7nG+9ANecxy4iebk+SSEu41ORmz69qtA8AfAXDxW/iL
Ds95l1fTcNEw6WKcmcZ+UBfQlFnk0X4lw5j2LgGFusP1sNfn6W+z/haqA8pjCyzMnH2usfdK7qOS
RDOJiKLc0qalb1ID8FgLbk5jEvOhYvHgB1v2D22YlmYuiKoYM7SxSvQ3CKcBfe/cs7LxLpeVeT/a
97nZZA/U0ch7pRonW+PI9TMBl0oSctM6aot/WorDtUlVy/b/tW955mUpQ/5lNF6r6vSE8wGxMWYJ
6bUoD1HZf67PXLRhkJW62ghENCyGMdyjL4x0XJ/yCmoigpWleDiP4lRZH7/EbWl52+7l6nmrwUjH
C6++1ajzTdDGEwMDcNnRUkzi/ssfFHeGJa59N+1ORNuNSPvFOP4tAZOcKg6bJsR/4XkZIWJ3qMxD
PZNq0btcDHCOZyPEhxt/61wdoQYHXGWq1f1t52y54iqE+HKE8nM3PrZaOpdXZLvq/AGwqfzMHFKE
ZUFExeSIGwLHKDoXcBGqlPnys3cs7OGLDYKwwoIwQOAtSzmA3Fmwf73q19d+MV174pF+MP4Svu1A
kocJ9gDsElPmZtjCDzVP34adBITEc6kxthdmBNgyt9v8GvCKt2l2vX6NmZ+jdTYVNpXTM7+iDcJ4
3bKQv5NKWK+N3BR18Cqt2b8XMYiT/vAlB+5YXC7XILz2N2rmbBkW0CVVbjk1fHmzof+6uHiu8iBT
3bFLWrQ0axr2AapybSNleLf/HHOmUXO573lrKV8X5P9gQlyNVdDYLXqxubT9+qW4wA0fspUF38q/
YbdsA6d6LO2jOEen/jHLNP1MGPD417DFZmNWWeOzYmPSSWEwgEx7yhkL6ZygmbFSuZwuuHE723f3
ledUfeBZ7CfPiRDicdMwNAZIcAV5oYtgMr9iZmrgWKgjXBS6uW434Hh4Nplzr8RVQLSt4tL6/2qi
/HS7OFKtRbI7D01dOjk3KfSJ5x7fVoU+8nLfRaccx9u4mzv5eJI2Iewjz5xTklOBHqTcKUr7mgWO
FIKm3vhDnpeJvlYHp+Np/BhOTeJAhvidTfo3F/spTM9o5qzhPb9SmNGRdAXQLbbhdrvcmdE59vKW
YHj/MBghIUhF9L+5rdf40xqaIlkGmGZ4XGVeNbw2iSnvG1X/NSLmwsrcsoFCZ0zFMnCFd7IBA5ME
J8/zsU69CE+9zL+SLGA+1QSuU1bgDSZjlSdS6/M/wcWwzSjpYnwvcrTdkHoGW1c7A37/SdXO1/kh
WJ2/lFbklwL9g2NTK8YXlMpX9hyWyJmuzzk+2wKJaK0MKNRYIvC01lSFAAso66fsSfvSVMQVcYw5
kZYjHatKRC/tuxaFQguz+jGhM4s+Fa+DxcUMdhfxiYCOCMKKH/dFM+sOGGia55I+ObDwog2qm5mL
oz1GdO4sbD5shsxH3m2EHOMnOprauHOq7ChQwaIUr2z917xMyhon5fqlCmCEtTBX95FYpy/gS3uR
ZKSa7XOoqQ4wVok5+HI4l6lmsjaz3OhNH4ezLT9XsbrXXFicYDXNZun3TM3oofSy5+KgOM5g9dcP
F4ORdZfk23hlBN6U6cfvVxd+9XHsFrQN4djUQ/7TmQd6/molQZUyiWwPjr5VX69//y2C1l8niJEP
d/xjJd7gADXYCgIRXKOnIFYvy0Tc9P2v4EDWPVl7sWYnPDPrl6Pdr6WFnS+BNmZnWP9ZUgmXnGVS
SDSjrHSh0FZLqSvi88Q2XGYCihUKDoY4DjSWWtMf/V3w5LxMxU2VVevWEKC4sJY9DTy3D05mYHTV
PLUmeAl8m/snU5+OSKJxkqZ5QPXyMVH6LPD6s7edZfHffXp2R12rgygTLmx5Rnt5vU4aMfb5O8Yv
2Z2xkHUsZVUjDX2GkXU/O02rNYIx3i8xBVxkLP/Dr9+fMO7+OpyfxfIxhxms9Z9KDsmw7tBSKU3u
SQ5QpyA33KLozjbhJ6Bbv/m7dFzK7dAQw3QWNy/sptbbLXi7PkP/E/Z182CW+AtcEacuoTOb9pnt
I4H7CaEhM55YNIgQ8s2cplZGmfXR2329w4Y18ndU7hfc9p+9L3Z0qHREtc/LPpIxi6JUjV81sXSq
KAmmkB6zdlVE/gUOaH27Md0+DUtm+mk3oEA8u9xuDz64oAqGxfRk3CWGWQEhw2wKCyt5yEThocR2
VvxwkeHI43NI4Kt9iZpsI9E+a/OUWiXDv/nGdODFlzhLMAKO/NL/pd6Zj0rWxayLE3mL2xjdqdc+
hNx6bgrC6LXSPnLHiKPXZLfBRBeqF3F9mZygwCmvREH5WanUjE835lMNiEnKrSbpzY/arDJYNs1s
QvgyI/0qaK8oyKXL33Pn4VhbH3z3seJ0fQ5mIGzQNQiSoJfy3xxwjZh9uKSidqHtharqAoL2gRB8
GFWx5qXE7/gRSrhvQESJDGME7EOV86LOqvdBhVcvJhEj0IkW7Is/kF8OT5znm6Q3Up9GpDaIU7eF
+T07iCf7hwhTA6M3K1VbEjD3mAaz5RzCmPa93eutSBHXLBgRVpve5cQtdrs0QeIHn+vBVlSFDg+8
ZjwhhwH1bi284d7AxrAxUbbC64KQAOAnKPqt8Qx4qLwVyKnm6JTaU06rM/4FKogoRmSPeNK315uX
ApiRtrmtzz3w79z3n0DcSUEJBEO6g/wJ1TZqBFDI+vDxvmGDXtmM59+AkVcxQTAs26Ve5QYVMZ4x
qFDVW3IvkFuEQRJH01iZcLM1+IOnKkkI3NTiK9d14CfGcFSmG/ofsP7Y3EZpeAE7ZBy3kQJLgcEN
mHBx+yJfiwuf8VfCTS4LCiUrCnRX+oo7aLfMxl0woGfnpI4het0ziXJzrUTgHnIW9Ol1IxOK+ob5
fcv/W/cXWl4SQboC1hBqIuQ2tg4ZPfcbIBS5Om1i/mnaDEDRTNtUJt1EiVpQYqFSzHKCCw95xzeZ
uCwGtpJ+EkBaBgK/PFuRx13j8XX3AQOJ9R8Tt+kMZSZSe1IZ21YNoBriJ9ZCkxyHH9wy8V4p3PZZ
QJj+pdSTLBWyDl9oIOkog+OwLa23q8rWXi+jih66zoJvJaU1CxYdZmz2UkTI2oEyJjKCkq/Tu+8t
9HRJpn1vjbHpUhOzueose/P7a2I7gg0PxKmGYiyjWxeW+QQDuEm9F+BejjGoxPzM0rDtlJimKfpC
plrCDKhmFDMb9IZ2iwSD1gjB2TGPv2fCHFhhVCIZv/FAI2oR3MMa7fWe7SWKIdAL4D/IJil8sn0k
dhz1D8mJUZaWG9Mq+21LbyD9fJUVfxg4JhcVZ9lYFxbn4S2wV3HTmrpZTfveWbSpc3Tv6xiyoVQO
xoB6kR76sjYkvJtqF9BXVgJaOVW0Yq20GGvKVtS1rqAK6f4068DQyRTK6FFrz9rIB+mg6zr9U5oM
jS+/nFrqw1Eeec1yi/Bor3vVlEbNvWv1Qnlki/IY3XXSbS+2e5EA7C6agmtW50YlBpsqW7yPrGCJ
Kozmp5QS93DqcWUw+p7swDARthYYOBZE0ROaNkQF71FRUgZzBupaiWeEg9yjT39GW1c6Z5S+BupE
wHklK3YDH0wFmSsWp3BVrzLJeIQcr+26byBgyoPMDcJn9VjojnAcyO32gxLPuPs12H5ayv0nKVJ8
Bk0kaAqnbIM9jhVUWcJepGA3MmG3dykOEUpgvgnQ+uq7u2OtlCIZlSVqY6F74SNJYIOFBWurZrF+
f4aBIdWFuTIAhPgi9ND3uBSDjgyBBw3sAv04YBUR1RbpdUenQKrlEbmNvSwdulTeHmPE/LKyjQc3
2EieQKf7Fn/HgcKrIx5YsiUq9srKFv8T28kaYwA7KAz62B/gegvON+2IOErZ18Yv5UEE7VGsbDnZ
S3nv+lGFGbE2y/iauPJGrz4Vq87rZpyy/bEvqyx4KNFDdPU72MI2RyVg7mpt5w4QSygauvMT9tp9
jBle4yyzSU6P7eiNJ8txS5g8Vq6fMTJbKazlwPq23XOruirPZy7PtbJDs3rxnQVnK1BqhjJUqMEA
HtUBVcdc/zFSD2Pdcovz1t1BedR7aTyCFMoCtKzjQE8Pd7rDt26DtWDjUZci8SFlgVJOZ6OYEQ5z
AsaEAn8dwYHG80Mdq1m6Qv9LSaj6u1OL8bYk7Ck4cMnqFpDfsVN59Lw6rv/5KerFk5qgXPeKnhrR
vrlwbGEndZD0PTvi1UEeBir3tSrwDEozEdPLypdOOnlNi+lH/4luE+gK1rem57li5/lA2Qn1oZ1T
6l9Fe+8hQ0iRPjtDG1zc6238MBIjtOXooQkii9Jn0yaKWj+J+Y7+t7FT02Ni6r+uAtJ1nu0/OXKQ
Qw13ou8ZcGPBI7Gnm+ZsaVs20WSGYBcNMi2WUDkkibL6kZMfQKzxj28zhG1z8Ti8TNrKrfE9o6we
TpXaoJNv2RhCYfAl1jRa3O55N/WuSB6Jkmm+dIT2C5Ks7YAuS8CPADRyf6xSl9f1G7f9tDLl98Qc
vVi726Qdw+FW42b35BReYp5luNqfdyM3bDrSnBT6+PTu85yIIePrVlfpMx9eTUXmluD6Bsc9lcJO
HMNyiOR5Lm/NPzgexWg8b/gEYpk+swOUK6XeGyzFpKBZ6p6B5sKXsK9mLKn+24on76ahgKJvRGt5
UTwQnVkFIyeCu2/n3sP/F8dtchtkKXNqlamH3aX0l2P0aRc3M6hh0xdRYu9mrXDTDHwJOTDAwbuX
OcZrdWhRfURYQDxBjd/vI0ygtg9NHSkMGVrlLI8DfCbblSa/z9Gp8FheaNQjz4tovpOelt+SXTOk
oXa3ikxw+2o38wtyzq/GgWkIqh9PASTELUQhF5qcw5YfRMVDCqUBysF4ub16O9H7XAkEziOx1Yt5
TmARZxq2Lbw9ruMvlrZTaaLKFLxXQ/G5OBTKKj88EePdBjPz44i34kUbzYjTpVB5tAlbs7lSxzKP
bd8yokVW76Dkw12yl/1+5pT+ZDhbvYS5nvyaMdxO87lD87zscYnf3mKDwCwfBMn4B+8zGv/QQfYw
1WG5pf2CFS97M2n7PXrIoGcy1XSrVrM+MmTQQjNd7Fmdvopkfx7iWWZzQ+l54m4CnhYA6PqwHtYz
1iPMO/nULn0F74koOsQPj7oqmQjFFOmjieGwO9aYxeTQQhsNYxml3O6qhei/HMlXILCfC+zq1717
nDMH76A4IErMYSQti58GY6o1IwUCoeHyZOaIGXpzlzYQa/DDkmkJbHi5NYmUxaH3eij3g/o+CV0s
0DgFP+J9kCXE8LI1X+11i/oXt+H9p9dEVRCJfc7uM3AagohfH0RefMmx1+QF0J2gYsiVRZCjFt1I
XHwB8VZvnLrzdglISWa37SI6Hs6nmEgE0vFFljsBS4Ln4LmbK2AMyLlVx8u+k1oALSQEOO48X6CZ
dwJnIgs4mh1EGZEwib7r3znB8NonHfGgoqgVmhECQ/6HELuvVk6xL3S/+5XC48FLkj7hJBSref05
pmUCym3a9uKTlEWXVgtcnpWpL4OWVpEIsdRL/IKe069XQD4YwY9ZqAGzaViuGUPZREfnXS4lwlnh
8t5tZZAV+qFxY9dsdIqgAfB05EJDjHmTIzzHOmsj/h32pYwZ8e5T7yWPS5h/GqytfLNm3Iaw6xwV
eqqZUNdAcaHgH07uoVRcrgQJeam9sMGBvRbWUNF9llusPMb9BGUjES66hC9cMXGJ0vqaamvink0T
mCS+En4A1xLt+XE35zCAIfSh1HTVnKzpPL/Z9Ofcfc6xM+TlnLowECPRUEhIWWDk1CiegZGPYtjm
icZWzODW+0EjTHTMnOfU3PvQMxNT7oOjRRxSMGT3xDsbYkvJdDWtYYC1/lATihjv8qIwQaUjM4+4
/4vVM2VuAn8s5CjXVqpycyGPuhVSwaV5TA73WtRlNT5BKYg0qjR8qlvxJkCrtAlck3tsNvrClvx+
tWYQ3GI2tmwCOiiPywfxMRuA5qpgdL3jtBJ5A7jYduMa5oLFC/whJhRUrK4NoRiLYDiMoUyaXQ5g
SyK7og8/gRULzoYsiTrRZqfaCdk1LwC53ZV7T3oWGJ+EizXLbkf8N4bmhQM/AxOcVjQPxvj/cGBt
NyHy+Eyc6o2Zt8V4ZLuhTc24Qbq6jorchXAOC7P9NiBZbd0fgtIVTV/LlKYAGclo9QmmOiPxSLOo
DJcGCVKj1m+uPb9jjEjrIgJHUEwZ8AWSsa3WoSEBDpxdbsSsjJ3lWrqEJ940xggwGRmXyb59PfkO
jcXScvSfbTE4CtfRT9o/JYmTkQcps4Nmzp/fz0IFa4whJsKD21EkwrpHGM1T/IHhA03gdLdK3sih
XBmJD8FEZJm3r4msxNCps2rVC3VPrHhCqVAK376Mh37hpH2m+ZoCWxQ52Ze+eXWmUN10QZ7onI0k
xbdTX+4FrQqrylDlpA1h8stByDdnFWdyfoDX9BDuSbaFZAAbMa18soBsTI8jxa1sZQs5Pcs7w+5f
+zguTQoBgAWIXpJJoCow2zWe985O6vFp3bq6dXkVKQYOdHzb5+odbz1LhM8efnGRQM1qXVzcZCSE
2XylxjxqUgaGS14ogJFKlr8uLEDD5b+Eb+mDVqY8ZtTcAXg7heSOwDaQ0bYTFTkxITxjFBaRZybS
DQ4xZf0dRphBHr+McuHV6fCMvXTKuXa9TFeEppXt50H8xK/wKEAb0uQ5sPesRomE/4G2V+03bkMk
KOKEkcAuDTDuhuajehkITfvwXH1Q0pgaacotX0h6URkwMZX+CoiRUQx+y9+2Fo0NZCmL5Df1N0GX
I2SaeGkAxIUb4Z0J3zjM1GW90h7SgDTL3KYD4AKYH1WKb9JMEII8ykArPZGE4qZXUFejrXZD8l2j
LI6KgDaMm9TJjpDPmOnkgkttAHMiHz0SHrj/HxRZWOtEhXu7HCwTU8oOHXtJteqJDGkvLbBkLVRD
6y1gLnHMM+awxDDlS+bxZhbsYEz82etI6COJsj3wHFWBeAU5BozM2e0VqdTWZrEI1iaBgzQQuElQ
3RllKW3j39YmIo3Fcnb10Q+hvgVa2/xLIzwVqmf8CWjpqLdl6AmQWPU8t9vlkozckQAOX3TerD5I
+ZvOoGmkmKpkNkkkG7VqedFRMzPMSsJCNacE339+Mwh6QF7BgPWbg2O7Twxd1myxgTSAXvmQ4pqV
eivT90qtLL9JSpmP4t1UPQzkvTGIT1EfKTp6yLTbgws5+TTy/QAq+sRFpe0hb+9JcfsaeEdFBZ0Y
NQId6Gq9dlr+L84W2OoFWeux9Eu9LwsQe6wU18y6HgXrxZWE6clMc0Sy4iRXgrvsH2Ft5EZmioWH
qh5oVP8+Hnii+IAI+EkbhfRASNBChAb0yBPgavnDT9nMXhoNa5/QKKymTzTbTQ1U1wCFXST5xEHH
ZeGw/89Xu1D7vCFPTKh7Mqc1STez8+zcGT784KtgsgYwKHfmhtffL+hvH8rgL37oDRNR7RU+Rboi
FXChFgpSWU+bJGv1EtENxoJewedFyYfjNObP9b6lgQpGhUMpU65K2FhY0MeyJJj9UXNgrpIOBG0R
H45WPnMg+GzgimDzvf8yjKxtG2BJ7cZsWXmSlTfP/21yUvrBTwCPR7IlpqbexU0c/8Yi7cdCSoV0
EXUUxZdLl0SNu1Hg14Mn/ngx5WztO6O41plj9q88QGzS77TMMCetnTD6vEk2MzfN/jePRFTjgQQe
PtHNXEb1/6EstmyO/nCSRY35fP4RYuvXBWiiCWluDZSKW5NXrpELo1P4Nxhi6IbyV0kwhR92eVmW
DpJ1OCwtbWlkf1ZjHHAP6kyxC5dsV8RHDwBV/oVPUzGd6/TUuUVwE8Jcp4ceZ24uLzABV8zUFCwU
bYY1J652c0vewQes1gccD/Xk8zoxag8mlHxdr0osMR0kY+dDqUBb6PnI0Ot58XQVMhwXTpTf9d84
qjJsEFGiHyOLYEGsqrrhS7jgSzBxwVCaAfAh6Gs0koOfTAUP7VUZLGHQ9mIvIUai3JMnmo9RPCQA
aXRTvmvj5z9sWQxImfAvZR8uLHJy6jEsbhlVOEsHdERdVxF3wPVufZ3f0wTvUMcXNYiC2jDol1yb
3voqVDFGDzVSyggl29JNFdPU8rTUhXkdXlJLOp9NbpwzXwxrok2ggSedAWzB4/tGkUhIarTIS5W/
bA4Dz3DnF4PyreNEhYUm4RFNVhWcRwOvZEoVclDrcVB2ZD2Wlm7KMhQg8b+UOtcleFdKsB0cxs60
mAakUrxaRA31+EIEIVoK06TS0I6CM/nKEpBag/zfLRhqx4mZXjXGrdI8a9QlF9woqx7d9Jy8Ivpb
iLYhYYiZ8cX+g/sQDCtuelTSoGQk+B7PXQePTJ2c90IqgnIqqxMJCjx8o1sjhy8iFohe6OFjYxd3
Qf+lL7nPNBt1WDDglb2dfh6AEvnLwZe+wLwerrtMFfV1KN9reU/8zlhZrg8ywIHO8r1XpdqWz6kb
Rnh4Bqy/cwAohfyrGmGV0l8FpuuTv2kowfK0Ju416jNelfZR+MckRUbMGOEuQ3hNMdRKv9XoNlsM
xr5sG2ukphDKvubCwnlqt/prv74/flFn7MmyG53/VKmSepWl28KOH0rfYgau8vAZ4rNXJKf2vqWc
Uz83p5zPAalI1UBdh7McWVsooVnq/GVqjUtCPIWlwQMrUuOO04pC5O7Hxv5BB7//A9Vbip45PtfB
wgS55xuSFjXAUe3O2uFLkOS1BVUy/xjeMJnVM++wOZ+Mp/2pY8/E4cBiPWcEo/24fBP26I7MjepX
m1nHSek4GtGcKCNZFnuDoYQqjlEfqDmwq4+++dBgdZro0fpcdzIEqgo1MLam3dp8ApLcy+TWBXq7
/lqkPxJZWLmB+5pgAcA8bjBBbTNtJHvhR8I7BaTyJm8JOMKIJA1JEJoktjYNRHEWNgcEj6kQ2yiQ
0r3fIdA5nNYFHmCjUMxYAVXNawYbgjUmrr5FofyyCgUDkFAtTnSJusJIquhYSsOrlhN+q0SdX8zQ
C0YDleRS2uAOPCVWlT9X1pCpmUV+6eGW0+o8L/xf5AANA662mWMZyscrbb8VqAJGa1faR8cmPcwU
rMjc1H85apXlO6Ou0XmVycQqXqw9H2rW+g9a+b9mepHfk6j3Dl+52MnFaTUsDVuQWEq1xSCX1mkb
MVWAkVTafvJhPN65WvKIS3q/A3w+bmlDUCBsqVYot/na08c5ldRSomyuq+NyFMNhDAil+PixB4tK
l/9PqHsopvCm7vXrHufo566z1ZP48Iig8Y1yA/YIpLOf7wBdFrLuzV1pS1mJDdLHADXQGAT3Gy2M
UPbvzJvf4vlVO4SNYDTAaVJQOnIrtXGJD/Zr3pcaDV2G00OCpEizMXwnoxG6aJ6pG3HvjY/X+ZDK
A4VoebwnZjuCzmXLuuVkearYlHFqZCNjdATqfZKeg5owU/GKLCCrvfSm4Ym85YlDWCHbmlTFuXCL
sKHV/wJTAB9je6wx1nFJeukFi8oop+GqKHWHWAF6Xe72NwkeUL5fASw+1McSHVhPnT4X6iI35tU8
/wH/ZaM2I2AGoDs24hUOfAV8idXBqLFFalw+SJsP3rQJG71ItDcfnYncITxhZxcbXgvvwTA+z4ph
mm+lnzfxJJMovxKPCNMyzEL+04eTxk07vDWXSzp06FwG7seTy5L0Rihoi+Q2Ee45dV7jhuaodgYv
UAFysViykWNycBnsa9OTvZGoBlqcbYLFMOhP1nCcosdjX1lKcIzpnhOvhRl7hynN2JkJ6yQUquiX
zyZbpc3/6DxAZ7Gc9u877V2ePAy8hQ06M0O8KqFh7SjngftqOFQku7cI4A2JgovLTQ6cs3n0mGlQ
nCL0OtXzTVRDGxy7Ak6/7m+e88knNPgFAS2rIaNg4x318s20pvF4auJeR5l1ik5eLnwikHGuKl1L
zguiHsTyJ0WaZ2bKawp95aiwhZnZvbVwhGU8pA/Rg4HVOV9wCixrSuOJ2civdIGAa4mQx+gktiEW
5g0S4UMFzmgUQgLkUL/NhyluvnLzRUnneYSbDWbm83qoMO04SMwmdRwKQNMLlx5LIDWSNiBsKukS
pnZCYXOt2WBhHT5tLd9MhHXIYb3EXodi1Porl5+xnS/qob+RBQaSzHxCmdjznt7z4bdsjx9k4Adt
0ooYekMC8Q51q6C4vCWIZN62dcQlrbZkcvbIKE6NVC2u65Alu8Fq0riVODFwnAY9KGqbVw5gBS01
8Kcr0nop1ZRIxTv0W9ZTRAEMQGMmhFwaEYJpLB5nZNN4mzlm04FTuHQbRdGgtZDyr+GokQS0bokc
8vSVB90bZUtPFJcbfPumuZOmuX1lraQjRhhrZMltW0FKXwMS9mFYBuuNorpFcuzwEYXMxZIqXNPJ
cLvGDXPTUF27kEUGrJQtpuycIJMLGyp6CThQ3HnakrT8tymmIDHnQWf+Mf+5P3GRJTwHzQIU/cqN
XdsXAegh8d4+xl/EHgqcN3kWMMVO0PIn5EZEpaGn8TRVTbPlmA4dgufajA1lMT50XquuXn6BNKeb
TnDOxTUyJ2BME/l2FGa9WREhFpxq9Rjp/HpHkvqAnxLNmr4dY0Fx2q5UcLbYG5XyITW0/46l0mda
IG1lzbzJI40l6g3M1gIpDxsXGnLSKrEPAUX25+w85Dwan6AhMMCnz0K+OaYRgVzz0Kb52ukUd2Mn
aylBvA0AEfwn7+BwLeNRWTQtibv2+qkKuGwslKJlvk96+F3KyOns8V42F/tUdohlW+60SefUONIQ
ugwW8ZqwOkmvlFB7a9LazpR1WnhD3RKCb7Y1wX+G55s5XGLMIzEO9lcPqJBRd6w1i5iO4KupiAl0
gKArP5TjHPGSFQ2ZmOMwCg0OxgVBOjcHqDPfZ/AQHHtzrgTbuF++j938W9PxQFWH/cqB9YRimhF+
G72QXnGzv6PIfe0/c/SBaAk0fn6yZTgacMD1fjSoIBBdqquLR8cBL2fzSK0KkcYIHvgtBXtaec4E
oHgsZ55Y/LbQNsOuG5AeSWxHz4vBDioAz4lcrZ9dAuGysCkh7vDVxY3Qtz4WlOKiz4yAaUkrGPLx
hVM11ls5+THun/G89OSdSisxVSltrzgcz+tG8Sc5VejULOaJnxpLgXGUxx6hhori5MLjJCH/DltZ
sHY5PNpWeP3HMWJqc28MhvkZd+gnhig8T+onBOYDaXjBI4Zi1exsWzWPy6gkU70H0cYzYdBkB+a1
fVDgOLmY7/Kqr5GKmho45HNOD2fmsmhEWcV4TgVRc2nndziqfvK5i6nNKW5wBkmwKsMFpTfkFVEF
hW1eopCtRHmibfUALharoLRxy4xeTy6OylWtcvQxyF0TwyMyp1MbDxkRqb67Wo2QIpz3LyYEJuX7
pAtSTcujiOv3RneC4pVd2y6jTSY03fddT/OgIU79TLpw/eBQKlE2sVyZ50r8nOwLJMiQ3tLFGFjN
akJOtg69omDfn6ptfjO/guaneTDiupjKpqCpLdbpqIg7bE1bmzYGtk7U0ti7c7HoLs/+h7Ec5lbi
T250mDgVyx+yoUVZA+fs2Rfk18sRpt6cxrqOIlkzOTorRDwioMV33ANNKbt37YBqcNYRkb7sopxY
8LDwsYO5bn2m0oH3phrtdM1L6nQtzyKUSaxgmNVwqTJiYqUFziqDpSqitspc0Fvk4aAeKx6c86PF
EfpZmAqjvg4jLLd2cchCzGf9SKmGwjmmLxvSBWd13iYBQ6GfdAz0v4vMfv25BZc+NQmIrH7AXCfZ
Q0Zsy9hCGXLxj+bAOrovqp5NRLfYl+z5okJZMABE65p84eKpJsHw04Kv/F5EvfYtwe69SpccUdGG
KC+jpBSgwd3mnuNOkPX5dn2ZiLTPGBtPerUBD32MPcFZS1kO8RbYQp7LK5UNB8D6HUynd6Fm7zx1
KY6O6F4inHCdAXuT20If58H8THTOxm5kONOjPE2PGBqp2Qd7sqQ3SevZrNxzcjEtrRoL86DKnCsW
sRs87mi2+pcWuDHAHyHc+QK0WDxKlfWZfbJUE3Z+xGNjv5ZoOMww9ig27XB6pSy6WniPI8NiiIxZ
101/UKraVDdkAQDXdo0BxPUQ3iE1mpFtTW5yW1lvEegK/7SWPP6srwpsuv6VaunoBOaaoN4WCvx5
k9HCZEORcHfkJD5kphKgSTrY94/jI3LkaE6gb0vd0xjmVD+/bWFh8NVZS0jql0j5OJEG/8IrdTba
+6jZnJjEJLP/gigcH7JkXCQGBSHZ6FbZKQ2ehSojyveyLxnMy1C7JnNH07izkJ4lS86Uira2TYqq
sQUW5VRIFh1PkEkcMQI+otzj9K8YXTRIxI5Fbg7i+h0TN/tQPflsXWOi/gV+YL0ny8DlH/NqD4EE
dztLXIWmu4yr+U+8BbIghyZTya7y8vcJ1Hc43/4ChrvEtx6EXRYzdt0CjMuF7vlna/6Zbsvarfxi
E+OxGpIPZQgCpqCEIR31BYlWMLelPRYxvgkQMTHh9BOnwreoiIGuFlphI6XpND9KGvhSFscAIJiZ
iZUibLDbLEgnb31BJfOqOTAbtUNsQPTtCb7Hj8cKXrTpG1o+g17cQxvPJuqWwi+X2ysx0Mlxd8rF
mTE4El6klMwsa7O5HjDt72fhJewXATBnljabhUz0HwogZjFDPWczuA7at9PXUxEYH4F7xQpuyQ4z
hogV1pI0xVTThAJw00mZLxzbqEtMEa2Q2KRGrCRTW8poGRYD3z1yls+RgqSrRWDg6xVZcag96Mdg
z03K7XgNxa/W8Jpp71+LdousMfv/CaY6H+ibOMYib2oqbBwclTzeJ31breRPEAdaN7EqV9A4rIDD
3vTdI5RNifFnv2Oye4WmVR/QRyx//PFM5wnjff19xmdTY6SpkIJFLuZ2iZVFW9PzKFGtiPm1FLFs
q2ryKfG7MomvKgfc8aCKid0YIxi5b7gB0cBl3tjSD852w+EQBDlEFCbJr0BzQjhSXmnjunma3GBR
WrrXTBxzwZBZ0at/glnsQTFJa0iJV4SUXruSOJeWihj/WcYizcsfAoxr2ittGpxk1CeOuq5DBmY4
BZwjmlA71HGAwlE4nOvrA6RCefOsuM4zMUj74GR7COtE6KDlN7wA/hGd7FOWNr4lxIXk1E7/y0rC
Ftr1UO6q8qw1u9OoWhe988aJbbB1GOKCFEL1iQZxo5Fjd2UPLTBhPr8VYIuDt+SyGczi0RCiDSbj
QyAo/VeCGXTWdRhtBYKD4ONqFDlI9D0r74fHAQ3ForLc+XjkSSyVNEOGj3ckyK0gmrzeSFW/Q5ag
nBPZoEj+HOfhXXxBZnGkAZ+kKNxNSbgvHxG3gJGZ/aC8+UOYQNWgC47XWl4mj9MGK7SDpZfZ2i/D
JUo2bLEseWqqBiBWwb0BDbmbniIydHoLhakSIgkCH4+9KagLDj9ylF3JrxLfuk4jKNfXDebhAtMX
rDa7ffTfTHbuLlSeFHmXo96cebckTGJQ1pb18YLg8ACJMOx/4u2+w0UijWQ1xpeCon4wLLrzrCQa
pEdBaNuhkBsO7cTRVYLUWEFkNOjCAXFqFxT615PFqshPFL31ksi0Puj5RX3V+8ZN9kKR9wQt9weo
havYzlygQawXw8uzmaDEEEJHPddQ2GQUygVx2Yz7+np8eJfqV855k2BeupBPvE7aIdFks1o+tZAv
E/kdHUK9/abTCPnERh6vkCy8Wzg9/veTmIl4BTgclt5LSCjVkwD3x2FWXt0MsA/1UyrxK6xuL7Kj
fN0BmAnfO3Ky5WYydvoAubTQSWQWBFo2jphDY/aTMZ8/oS+vhOXsqrz8pUsfELxngQvQBdThaTa7
0lsrFZh2rm3X6AF6CdA3LN0PM4y+/y541a8R52kJDYOf3T5+DRQd4Pjq/t66/nbDyBSwwq176HtS
K/PCBaMMDIchLyLxiXM7GL92xkIBAwRvHQ2IpyK/TkU/Ktpd2NtzbQM4RiE4OS0vvXYc1dxPXZj2
jcciE2ev8TYvvr4PvBZD/WTgl9InMEdLyWntUFdxNFbtJVlBD5dK/1ctH0mbupwdLOkof2zxfsnn
x/fCYsicWNv9DyNrfdanJslMRzoMLXGkOB5eG7encRVNdVRqyGxNEpVF0ydZf3L/mO374BdZ6wOJ
K19wXpgX2p55NxicJQM/NHa9JEsjkjMM43mdAaZPwtmbYf6/3sqn9uqgLdTtzbHTZLnqsEHJ/jR+
atC3VQI6aTHLDKTWk3Y6yc6Es7OP9P/WW1GG5Ljr+/+6eobqaw/kr0N/bX4KQD5i6SQbuS1eswjU
X6u7dR4c7qW0nfElJbpjJpx4ytmzSataFZ0THJXFMLCPf5jVtMBJz6VBB6EzjxLq6auJqncweK+f
UYQAn/vRbRCYq1lhaJaaelpPacReoenu1vMi7he/0Ej/134V2azVSTkhKcIDb0Vk8Ae2kSXw100r
kv7CPEiIHRsxHczLXkxXqIb5/LvGI3xWEeabWYbZ0suZC5TwoXUd8Rfw0W2fxNAWOS8eh/EtBxsN
mxQymP75lRc8ZZYJubiGB4Z/GpRVXgnAt9MpTDdUi3fPTWPVw6EiWHcHZSfQBbARcavaONyyQC/x
K8mghZAEB1F0FqohtD04fXxMOCzOy1NoYLSy+/2oUYOnwobf5z0AZTPmYlY/g5rIMUkSS2cZVVRw
cc4EXbF7+/KgnDDUpI+QIVK2T5q44lWZF7QZM6Ge5f2kAaYAraT6hwL+hAx8xmnYs/ieMn1qgiij
b9a9BoeLMOkRO8Ir7gxaeH9gNyCdchDJ2kw9Oy4/ftDfAgMuuEW98zB7Rm/pqwo1kiAC5b8F8Y37
vb27khA5nvKQaUBK44GpQJhDP/YzIJShHGDCjBUc0uv+QAdm7PK883VYP+iIGAhY1jtkU0lUHIyS
yHJXUcYFDTa+nrULh4jnIVIiF1CMiNaGRKvF/aV42Rvy1qrupp0nlDbg2zWuPWutcGO1gFrD5LX2
OPaGVO2dnVLvRtUiKui/Lff1yAf8zeFI4aAufk3R+vXWnvjU54ELFsKaYLU9a5kEW+orun6yKDeA
9f4DwqsiOj9eWbus+xm/CirV3/yCdIJJrTu9kD4uu3qA6CLHVrieVEIyjKHDg0LFH5htisEjOlaS
d3IZYWpWKCE/oUnXvKzAbXXd5dfaubFcOCKx6e0pxpXG277UPSPhKSy6PtTRECviq+nuSWdKF3yQ
96KZufjq5f4BIa7SkPMCFHnBr4G+MJW1EJKSNGCpwB/ice32niSr1RGYB/FM2JRdrCL4A6OVpZPi
J9wPPesPvwb77FvAUFlYwvpbPBSH4qyDrZoKWGEpaZxMXCtDDEtxE6K3S5y4pqC4HA8hcY7cyBWY
Hfl8BG41wmqOMDtpTyuTRiRVvcdYoJuEunW1XQFFiAdllSE5+MQhabubmbqbUfA6NEzFM862YbMV
HErxbcZdbcjlM+IU/JbWYqKCd/+iVDkC6eWfkjUSZQ2LXd5mvtZbAzVXhdgpdvIckEepOOt/dqOK
VgKrqYwyaSfLOLR4BOj3+gbyjclOYmaQ2mfNHnZJ28tSqp9XQoOaccNXDPev79fBdXNgqeXQFHYZ
Kw6EH5sJQzJPMWRkPYfQMG9zbhQiEIO2RD1ArmmSBHtytWt8xf2CTVnOF8i13fvYRBG1hxA+mKVO
RWJz+8A0tmXSH3+zU6P5s/TQEUemCvmn7bBH58TAdYaorCFnVxXEZ4vysWJAvziq3zzJfXjj2/S0
HyRJh4Ownj1FmtCa2BGLUVG1tV+1fV5dZO9UhwDmEYlg88BTL7b/w0CFHdGL9ziEDIa4seyGRQHt
qAXAlNN9NKA8GSIcuE3kAvZfDQN29h8lffEOA4XiTNWYWXnzd4DsDWJfE8PBmI3mHb8GlGy/bxVC
2tqkhfw96mnFTMEGxeI8G7kjpK+koOf0x36Le5geVs2ZArDoTDHYW80CCW/JTd3EdukXWiHxRoof
MIjT27ebr0V0GYMauSqHlIaBBF9szfx/CIlyjh/Wprcy4gFQFLiLjBrWRjlK01Z4WwUFglYsHUpc
7eGJOvCmak6FEWQv5irM46WmBId5qKLphky5w9amOwFfII+hazd93OjEzqqvejXmqZcVRZ0sEoIE
q+iLHSp07GjKOKlC/OuQy3qmDDA0My6wD4boxqeTy+qy4PLUgpaqJOGFW40f/EgNoPfcBvqQaHKv
qUO6EFDOMAzxvsaWT8BTlEkGkOekHorq4u+cI3tbKKVbJYHMukFYrA8GkfDkb4+X8m03xHcRC0wF
FQfq0c/VW3twq+phnbcX2p4G6uMzpcsfntqF5+sYxjRvNFx4pKK/5+bCr+zWdbGZL5Bc1sZL2pEF
CskOxpfQ3oyaAHQlHTcIUsUfXSeoSl4oG9N/hPWCjzRe8hI1WxGSm5O4MA566tl4h0lzcDDfyW0N
ldGNkCnTb/W/iU89YwN7O4EP0rfyX5fVRQb4/+w7aJvWiEVYlbS/7AhNWmMJ5T/Ko/aHfive+AlI
UjbJC/x22tikjdmH6/IPPOMcEwUQm8ohH8vKfjGPSkOyPxXzyC1bzuPHjqY0DpQWjyH3MqyZtVpI
0RPX7ymCDjvGWGc5c3Z+KYPTFqRNawy7yCn77uNyH5pSE6UQuAIOtt8MitRF/u1LcVm2EDFAzP6O
4SID+H0+T6E3yP7XxycjpsPQOn7M0cdV1EmGwyITSsQyz/r2+7RRHxbU3aJXCa3xO1ku7cjBc4xg
oQx6KKzutO0ujjEZ8KpVmeKlvgNStjlrcLzwGJJgmdd73B3fD2YLiPoiedG9V6X2YLz525o9j8iA
AswyMOYHQVnW5OXjub1f0379bcx4y7sx8Sda0t4b+eq5zQzXe649qPUDQkA7/wa+z6HMP65OAab+
CoI2rSmCrvJEmfZmsuZg0GsL2I8Cs1VZdq7TA29Y5WYT2TLTsu8JhDtCGbevyRaBAxwcNoGQjJJl
3XrPlNsPp0I+UyCIDKdQy9GVleDOgKbZjNdPCvryT08nivlZYapllbZ/nPUJA5HqFajz1g172IiK
q+M3W39BpJK7bAcLg6IJGsA+SsyWI/oWVhixgLxM06wmJoctQ4dVE8Kx/p/+ZO7Ldn5wh88yj4wQ
7XFuJToVlc2vzuBrVRZoq4mRm5fIjBnXYrrVlO8Bmq47C8rMq2xZ1czxomQM5smqNd/lROljc5AR
lTxsK9fDaPVP5VAkih+85J4VUZTGqeI1hd/ECiTvojc9YeefgFoKLGsKgYNdiYJUpQwn+YUgdnI6
8+dnHZlo0Q2fb6XCpQ2+Z4e5Qhr/8D/mGtwH1U4O6V5sSrGw8H/CJQwNCcUaD/beFNnGg+wA7g8j
ssCk59Hd0KIvzMJ4DsJWBr1qm8udq9Y2dyKgN/TJGdWeDVZXsOv2amYe0dcTAWRaQ94ZHEnsQYFY
Ix17QtJ/PnuoRRixol/hoSGhQ+tqxZmAs9e+9rGDFIU6zjTbXzDpY49ZJh/iDdMB9G+oMYrPg7ms
AnFXrdfo/A9mHxF237W4RmLfmBI3k9ZKyYq414YCXy6RvER1OOnJLRf9BFzLOnkdz6IihUOKd9Et
2B4w4a/Oaidq/YeZRFkEyAJoWZdyDLAT0B6ZKcSrc6xGKjQqqIN/03pHGjREuTegPpLP4v0O/Psl
FO2XPulOf2wdl6wzuGn/IUk9iBoYoJz3y/H9y0mPvSl3ofw4Ff+LF4uygy2u8dxHECwLXdlmMOwF
ovGiN4i8htsZsoyPX3vqtSB/pbGcEHtHu0bxGlLJK3ujS7m2F7xtNbIHdnc+cmPJt3MGvuT2p+sr
rt3or/HsgJ8GyitAU5awhBRu+BosHGt0/ABAIWADTx/bG5wVBF2A+RGlSSpitd5BfpdlbawLbOCB
lHZWQtCXUWWkPS9IAMfBsh3AasCvljJ3XTMlnYSyL4O1K72cbb0Arq/T7I2k3fEodNZlwMbhCcXs
ozS8nE0P+e+IVUnzUXptOKiEpehTEpP8AMOpjGiL4UHUTlYp4Q69JJHH47zpQ+3kXgC+98BRHmAj
rAglF+LQMC0VlFABXoW/ZVJGkqoioSNjTjl+C3ly0xEC0u8gyhUgTjFfDCO+GpS9qBDvYXTL9NbJ
lr1mZuWrk4w88hCgTcsXHesIUyA1kuLu5ApVCml2PzUhFH708gAP4u2jJ+FZwMSMoxjz1QAEAbRg
Aq8GDHgq3TmiaI/NXml5l8Eng4oqLmXpVsj/24EUEO2Ps+fzbYSdsgJRVIqHSrholkvCo3rZpkcw
DZEu3QduyHrDrbS5OgQ1F0M59/ALg0JqFO3nWRr2NENI5/SUZcwgwZQ2tfDWc3dxER+h+7980LaK
DdZ1jJfNOzmq7S/sp5keDLrBjpDznfq7DlaYozTnG/SZpf5L6kLlrmre9qQxgFASQhoJSlaYxP88
LsABdnAXVEJbhHufw8y3beKBqhaWoe5lTRvvPKOK2JN+E+OP/o3NS27KC/zSlfy+W2Ob9PfijbLc
kOVg28QSGo2BklmF63ZklQk4kZgKO0dgtYZI572FczYpzEoEhyofBxSd6bYtloEloKTpujHfJ9MG
MqM9t6lK/q8KePM3tQ5rx0kdsyr6CtHXwDUomvb3vMVNVxmpaINBcFKtTo+9GkbGh1rX88YvX0GQ
nCtsKtv98O4tHIBsDbFBpunHE/cHPbdRICsP30cY3gfCcm04vsZSJsjRUMhFmn7Ljdu+cfH9CDEk
dGUWiBN7ItVWYQxtnJvkDcMcKW81x9HT0fxZH/Bp9t0Emi6p7j3ErksRW/Gl41bOVj5pv4Ad61yG
VpNW3EOBKQtt2+s/LHdo9fnaExxgxDNqIKlAtydlkf0fpKLqIAjy5vyFWyccIRlpMJ5fsqfLun56
lUfzyIglBVA4oo8XJiXXcwtB5hHQ+MROEWs/FEH74WXTlflnQqsSzIQ/7GJrBT5NnMtsESu0v6fg
n17ws70nEfQQbCIwVA7gzjoK/aMSKYRCUDh+j89h87JcMU3aFj8JQ9SeXFvfK9i9ZNw09hysFMyl
vp6MO2izbrSCY/MZqWa+xMaj6myWmQS4Ghztna1Y6T+fJTlDnjev1iQliC237rmmTdk41NE+hUPI
tfc7trw+jo8MduQhLNpe1A4+P8nEkOI56rlvE7eNbfEqq+ihHZKMygNPeozu9GnbPBq3Mq37A0Tx
XW2FruV6jLLSqDWWVJUmbDmWOuxwmhS4LRCaQhGkUQh36yYWC5pOZNPulwRO3w38dF2Xx3jKYwUA
TVUReiRplelLXXLLr5nzgeswkuveUJlRAHanqko9pnasZ9A23oSGmmsEdRsaZHa0owY1IaCc3Pct
j8ShB8C3A76THZfqWkQvXl88RR7Dd2zQAfgrxMi1jdbNnd0ZSAYST0+mgMFPaPLCA/YQpI+VsJH+
6ghuZngQrU/mRfK+a49lk3KKMwc8J/vXlAKYczRgQTFn0oqYmSiZgU+uumiLnacZUyywozf7/duW
jF1DqUI53gGAwOUw4+ySVvpkwglmDovrJcV2Hep0chWD3VUEBfphGzDKfVQLorFV+vU5h29RvibJ
tzPPtuFPuqj3ft50vxBOU9gDv7u2lbzaG6VNxnpp5xamGLBInCUDYMEIyC1zOnKvoeJUz/vAMnDs
YHD6FMel/IM5lq+jd4ZqZNWvTKgBg1gjN4S/yw2guiF2TGQmaVgRt/XcEMqaL5bcCYZi6DPAynMQ
vIqyoN/SFrWQVzI9knTpzhjcMVcFaWMG+26WjX6oXoNF2CO2VRCbQfa+e3/TyImPnVSlCuSsfzBp
2vQJDk1RT4mrV0Lq8T2sCOiS5cTW9mMtea53Pkzf8yjCoVubOFUMyuakEzC7Mh7kUTHpdvgFzhWO
WCZFxKFzkZu2AehuYH+jEUZPAdbStcGJjCx8I5XcSSMHobGcDgIsSQCS5NLRyPD+VL19RbdN73gc
pvi6J8lrgYNAdJYgraDmR3r8oDhUrC+SttPSHiVpnTvN2ZkQASW7R8C+OM2SrkrRC/O90zeV5m7u
Xi1i0O1k/+yYdKhmyxf9hg5ia8RSeV6fP7DGKKu0C4n6b50npPzPagKn5E3O1L3rcatFhOZq/SVh
s17Y7QOkQhihE7308+HMBD2sC01ZCXmfthrCzR48fc+38vep1FI5lwFfKrKVzEQIj6jWSvFa5o7A
cpHwFCRqQjyg4JGAex9fSvShxNMvF6Y+s9gjBbmfVWazVegzMxyAKG0FT/yVmnvau/MKi6BWRTDr
mTMkNyLyyzM9yCNWTu3yVWJxE7wdKtPyGRl8EGTdL6ueS1/e/W75Dxf+kzQAWljDHCRxgksvBk4G
4J+rt3+FI+aICacUnTn1K6GR9XyBTv3Z2+VN9dniHmHN2M5DMYhHqwEIVNFLKVVmxh6/cNETCTaq
THynSDOBFVG6RF7uBZxqaP9duxVg+X3bslO/gDbDipSIm13tdafCfgpcoTsbh2wXwwdgij7MOA1Y
8IsRYHUF1oYOhm+OoGMWa2Uhi7AvzWHbSNOUpyQdCVj05eSi+kqN6KFZi2pEMWaaSTLf61E7dQ9T
9hK5gzadEUC8lsHxecZ3tG9kK4po0UnBZgqXzyiz9X6onQYwzq45WDBLzUJ4em0qg8DpLIW3OGDR
HtIvjSaYPVZ2VUtFhaSI1fZdk/5auCwfutLVtHUZGLpOdz2w9FHQlQ/K3uiHLPm0siyQMT8lpUFD
6CAU9T0goV63xY0Xk/kZjIGYZte5I18zcjYF/VGnCXskK7p2WHGPITbHq7hlGRbTyE7VoQduieS1
w7UTZ/u+XQuiA7pZIGuXazTg/OBg2RD9Y3F4FTbF7ntgY70PtqZwkI3c4iAjC+T5X7kKOUV5CMf5
oLPoI9s0QN97YTztc4T8aHLYl1xLfk52OVeRorqQytR5eTns1uVXMjV97W39XcxXC4E3dvZz9X7N
kcrmzOFwHH6mMfayr6tdYatrl/IBrIpHN2gVA2UprHaOuxgrbIkrcv2UfFWAMOq5gQpRKHAO2ri0
4agdK3LeM8tEThlFdKKPzno8OJAU1/Rc9xskNGS5YrdLDB8uvojQPlxaF6rbBxfD7+kjfeAfsJPY
VlsFayY4IER9uWB3FAotVDoVJPKxQC9jZ/nT7D+sTsRjPA6Q/1QOgadJoxfPxvUy/88RkzzBTpJW
IDJOWKwsp2ocP7lCFeDqpbx3X76wXBDqNjPS5z832PgnHnB0EeuLRrgc2PFexlUp2s6vjokqaYm4
TyLfy72zkY2uJDbivw+yddPNJ1SIY95sNU7tqiUBeUEjgqLhN3ovjNN5/sKGE3aQXLIuhYq8gT50
tm6S44Fsr17ZzuY2ykM0Xzj/VmZLb7hVu48Tsc4GTUbXH0gln7EsGBdwl5x+fQufz1XVLBLjgrYh
PYLwttTWS09sL2Gbpv7WYxjwKe6eXR9rjWLVYmtlgms97zqsxQ4h0debx8PZ9Sv4FoK851HdUqBH
hJW3oL0TBZ47d34tihuJTmrUCx6m+JzxJ0h8hC+cYQX8feDRj6YeT6i10PfP/TxZzKZeWnujSRlX
a6YtPuE1c0IjC03lOvfH/VC1IP7UckY0jcup7nUGSJUeab+3h+ayY7dElUHQpXYkX5zKUL58581P
ZwgL8+0HfkSfROFAooWVEzVY0DZ52BMyAEhuothI/PquFkoxAtgQN7QyAqAn6kxWEd/TjkCEM3mC
w+P3LCK/4aFBOvj9OF4Zz1aKDFvBxGvBiC5INoEX1j6gAbj+eebr43begMCzpsuk3uvbn75Uymf4
vkHmaZw56ioaHSpfi90FzkUDcISWoMhk9R86N/4pXG68NAOG4Wdc7RfkjIFACuejaI9cURMS44Dl
RGWtj342G2U1ugCUqS1Q1QFwR6i7KyBNX/uraNw0UzANUvUQKtRP07vew0T9LlSmcnRYHt0tgBxI
2xo0tij05n9pF/enGWIRFnJdbXLEXcC1/Zv0j8KA3NaT9k7yLgGYtLBraU+x1VZ/nD9xDsa1ntln
gzlRiz8iJG9rSw2YU2Vt7VfM9DCdWPYGBbrBBljoh+TNwGcRxekuPJasnJYGtZunTFxmn5h8yzxW
CGxRPVcuTmAGh/AFmfeUYB3x5RkUeVBtNhXIZbE6jOj8rTsCFJLFBk4kSAxO6HzGrrgvtGP9mV8B
kRezLRT9YYES6cjlyuEnXU4IwpG1PKzKChuTGQxdr19cRrDHPNoPBeOAAWZkntaRg9gKsp00BNZI
3N6Pm8EzXFKRGstg1JG83mqBl1VxD/HBLnYX8KqJMXVHzwrSqDPVqg0WNzTIn2RUp8bjne0E4GEk
iSNHPE1D8clKVBbEBZlwa8eNTjywwILFZioCDAmiiOx0uSrR15dAnMwgCNyRDKtBVq3CMUy44VAv
2AteS7q59DGuJObDYFfjEb4e/ADtpgJd4Yx19fMCej6hv/0Ca7db5DFjnbw3OvrAtNvkMLxs05QM
GqTDswuAzUB+qHookQYGdyE6/nWj1SYPKzeK/3EsJ3L5llMPwg0bz/WgQ+XKkuzV69gGdcCV1P7J
6bQBuALbQeWSZZW4yiIPWKK53m9CkgtcNQNMQ1wveTXn8NukhCAGrD8T/Ev1Ap6OLsL4Apu4wFp5
Zcgjm1K3M4gBHDVURpyDLc4eiMMcRpyrKeBmv+CYECTvfCFDIMDQu3c5csXMhFYZH7KkMwL7IyaN
9r4/EjnCVbiXTWW3Z2aX4bVYNVpXL5fAef4IMxnxB//lUaSywKcflS6b7ARWcoOMepzDGNfutQhN
x5SnaFzILjihe091ybviv3ngSYoSNkkaBMQWY8eIAZ6t0TwGke9VGNhbw6MN1/oClm0MfLUP3oOi
iFRrTVb+ZNRiG2hc6CQ1Cds6RgRFWpeAouPx57g2i7IZfXYNNQ/buiwdkLxCBICRifI6vFHTsjDM
nXmwiCRwtCqbedzSRO1I2LYnIODDrP+m6WGbOlQRSUHWmo75mtjrS2Jn0/XJ8XHgyVwExFy0FY+h
zurswLaK+NHnrp1fBiMq10L8E82TtoMSFFnu27CtK4xFFBHT1kZh4Sls1a1zbHOtE0JXu0CgPg1d
04Mc6xCGJx8pbu6wULy+l2hdD6Qe8sDGu28o+QOUOcn4xzLfAjjjp/+Hi/vW1+e1YHhUBCkrt7Yt
1ZQvhmfJ/ajzvACj2JNNEJIswoOeDZP0wu3+p82ui4seQ/2j3XvMbX//1yCZYl8bTF/pF0+uV3Ap
1fsuKN/VPpZNvBrOLZoPVg8x1RnEeHEjG2lJ+yirFonqyzrzHpryFoUngJfBbitrm30iEwlDGWMV
VwoTRqILjJ4XPceNTv9Sb+GFlwb+/HLlkR/8X71/DbX02p8K1nPMZu9EWshqG808AotV7MAYLmnZ
ZBZXNXRYPoRJdkl78olIYfEr/CMYazwP0NuDOWzO/z88Xnt35+FH4yoHn8YH8FNHGeIKhQvO6oql
J08k+P20LzK4Wmwc74yrEiM93urFtogVQnHYw1+mWJ9DxBppUQB1LEh1omF7LIrbap1Slj3iantl
WjVi9yYgwajUjvrHEHM8VEmja+uRUN+fYPpLYX1ljJNnyGkqmYvSs0O1qfP3s57c0EPqnNp2HELv
BVK/IZrKngO+RbfCn8jvrEw2XWWSH5ZDFCH836DUMbo32g6DfhE2pE3HgFem7ZvENPVsH7CXvo95
Rj55jAoUQKTdh9HwWKt8SLMNsda2p97EYFG8qtKs6FQJ2EYQvggTslp13hM34coha9etU8PAnvw/
r17pi1MHH76lc2o3EmASvDvbK+GkTETpmhDzQ8sjMrzBiRasw2rdZxiau10RpXQW4F6a9Aw4IyvI
y4o44PgpO2EO8NfJKHi1eJUBOASLsQt6lCUJsLkDWlVV0WiFAfglKL/RmwIYzeVNJPib6+FeVsdE
cKP9ly9WS7rvHpCrrYLFGqYDLHYtq5+67Yc55nqjBAr8NlbP+R7lQ4hbH8yx1tMHm9JLUMV2Eg+T
ROgPjk8mMjkOb9uW5bJ64jf2mXNRIHGRf+/RZbMRdWBbp2Oqwv5K47xXL/NCZULL+9eU5PITJ3LK
5nRJl8bRkIoMwPcbdP54qQA0wXbCh+Jj/sdHbBtotTSA2PQhNxmnOY/zqyI3XkO+vlkg9aTK6FoC
AFXHD/BcjxxRpranWdlg3ht4KCWmedjJtOhSgaFbGoJbbOtjmM4Ikh7JNWeR5k1uHHSE9BpWcBXZ
WYewMGMytbIUHM+7roFON61lsRJgMJxh1ME8vlesnZS4IOiA7D732LueOf9BPEgYeaj0UFEvwOtx
tNS1ncxEK8dxOMnNhrL5xd0Ypa8ZhKeE3J3zLEUS42h20tkgoDkhUl115jthZ9SsnMrb4ZRnYjod
M6KGCpBvtKnwzNTkFLsZRQnWTBqFyE+teZrgvmc6EfMYgZ7Y4ZGzr4FiqKt3UhU2T1RDeOUWAcGt
28X9JQuwqJ4bpaS34Hl/ei3g6QL5AzoWFCjGBYOjuI3PD2gn10W0BU+lBI7Abv6MSJYteDq00NBC
IsYVPk7zLW72OQlilDEk8loqDLOV9DNxp7h470QGDOy56r3rXfP8pj/b7W0pICD7KnR6t1NyaJ0G
VFYpWxD7T6vsSPm2Czov12kiD1Z8tGtn2/QiPhGxLaItBzHO+tY0L+fQzH+tuo88Ah1eL+7HQtQo
NPgdx2FLS2Qnfchm7brJMbZgA7yxdMZVGQVlv2Sa9343WgtKSxnUlUu4QZEhqrBKqZclQyhj73y0
pmUwNYHBmm1BMkughkUbva1oQzzERGKE8h7CupNG18S0bmW6OGk6LAq+xitnm/AYAI8XIglKdnHX
JiZeRKH6vMYFJ1xaL/JosL/GZFR7dIgwUrIR1dpkOlfAfI3l/ldFYWGRnSkO7/N9uE/BDuI9uvn4
4qUCaeNToEuxNQnkAX2iVv1oWCuDDr5n/2NswzUN2ykSxnn7peHr0/v9zoX8PancONhAZbVfemyD
7bWfo2y5nlZ4kPLQz2H4r1A17LY1vkh5nDAr6cwlKvGD+UvW52UysCHUAq7VvJrbaxijuqFE/6zK
CLzBKIuKbKi1hX4PrzUkQbJIS1Al6ndFNIgUj7ik2MVEe1xJUu+ikK572P8P/9bb/gwTUSZ6q/cM
kNFXGv4unLz/Owjc60tBU6/tIMKGApFmN8mso/WoVxZo+EWQMiePUKgbM/oEood9y40gSYFJU1M/
wc7lG+3s2R76LB8djBdm0WwSvNcI0y6PJVGenAek43FZtuKAv3nesOmBSacovxlmZjxjVAeBs50I
4ov1rVzBLMj55NBXDrxvFKLs1v/7YhpdNzZa2OtPIIWekj+F8NbnqfKwukwyBGZW9eW1HBNmVc3P
/4bp8vePz8KegRmoezPm9YnPbRAcMBbS+xE3F1AiaDRdGddBfgzftI0enPi6JkWEdf7Qtnbb+NBO
N9wop1z/TwRwClRT7hOniQ9PckYFlm7OMgCaYesaqh+bxcrPaZv5EvAeK3FsHMm5IsjiLn2TGJqo
tVvDeL73M/t+YIUm3EDISGEeq4LC2j4qP64pg4BmXm32kdGd8VIDyFvJSxBsJDnwWuon6jc3dW8U
NVF/NV1WroGlrRBAgZWAgWKInICbhmTy5beL8fjojj1fPUVOkyfqDkk/IQFepUCnAvPQmA4JWLyk
pZJmTzQ5mhWMwHiqhK+lF9e6AoNf3vxdk5dtJS4hRw0Xj3MHBuouIu2ya1fgflxKIPbu2RvkcUx7
9YeHLDVPY7arApPlikhiejvLf1O/sVxams/kCajEu14qwmEox+mgTKYDMmjobUmN3fmjb3au6FYt
7iusGThDlmzrWobdKgijJs2sUiGkLq46mK5BErVaFlqCrJSYiCDG2F2JaX3mUmf8MJxw8lzWpPUi
b3Ti4o2jnwirWZjDYyv0VS0CHa9zBb1R08DcDyn4UX3AKaqWD5RBIG84E2BERtqve1+s3czQRLgy
DT+f2zz8yuqmClnWbQbJRfja+/Lgqllj7vfhlt2W+AWcqRy9+iheXvhWeiu7R6l11eNwWwHYHMKn
5triIrl9UnnS5DMBueFvKJyjaEkLB872r5QW1dRcm4/bILKi2dqALWG6a2866J4DYn1AWJqtwvt7
mK6POPSeIvLHs39o37ixuyqkVBkfpFu1lGjINNElmYVwtalbkcxgtrh7i1zZSGNeUrKc1Nk69S+j
2/tcyhUrNVqWdtEMO0RlMTr3hM9ImKljn87J6fu8EBmvNKdh6yBA0PoMCr1aALiqr7Mi5S8J6eb2
+d/7lLLwEsPTG679kd557ONDw7Vvyyu3HNExiHp5y+aUAJt9uK0+y00pZ1IXg9hDDP/g7GgPeuZm
XOpPC7oTb8ZtN+6nDT3CDYhuMZTcqfNWkRNDmVsgMLgyh9M8xMAucEWLHdwQOEgXjCDJj9d3/CXr
3BVskc08JJkrTT3747q51s9SQpg/Mr71mfyZL5Wjkegp8ZwO5Frl5oXDwQF/EAcDB1l0ZeOU8vvp
VJ/5uwnsixmCb8jkpAT4wAMMZ8hKr62/UhxcvOcv5fYSRoYWHSPN7Aej1JW/jn6I1p3lrzlWXvrf
xdJAQTVAaN79cD1FCKGJ4q9ozHlVuYmVhJ2j4TCyvJbWj/v6015bR4vfuv2l9Q2q6hlp7e3V8hvo
cYJgoBxGJVliIPjbhoqJWJz82BV5uWfvjBLWE05nGlxBGGpdT3qiWUvEt1skIPm4IBrKeSsRsyav
pTMWXKgBGvhHPevCa61f+XXo/27JERdrSukVjeN/tFPdLPDSrGzCQ0fl/jgMuzG96A1pXK437Nb0
PmSFumYIyl7ewcvrM1tyVgTSrPh5aXw2z1J7pg6PDV83+paaIkk5PJbphVgH46lnVrco/wENIVp5
sigcYhSLY4Ja5RVFtmQkSNrjtz4EJQJHJ3hFcttSsFLaGfE3mZi6AdHv5PJ6H2apaEQAQHmLpvSg
tgdyUq88eXbx+N+o9nFfSSnHOkxw1cm+jXNSUNYmkcUwnwZstWWl4Vjo/MbGr0/hYSqNtVuXkE7j
2xl/9u9E9GAc8hRRp7eznZijBLJT+7ybXEm31J7TGEz3cgaYnrKJArPPp8ESWCwldz4DbleGrxzm
zWpR3bqFr+NAH8qAm3nM4xEs0di4gkxgAMYJzux4JPP0p3DgweBZMuqyedMEJeEpsv5vg6iBCm64
eVOQXY7HWljYWSYS68zsNOOeyKc+mtKg4l5GonA2fr3pui4EoxTi9N4BkzYHiYGnSWueehK7JZ4K
t4WExB6f4WgigJbkxeMLXmKOGEVKl0Dk2avMwoEk1HjsY/9Ul/qBVql0niAjjn2WPzuIbWTALOqZ
D1XcrH1FmtWc2c9opWkauMPjBDjqtt0btuK9bDaapYGvPMJpqDJEFLYFa2IXVOO0rhh6TtxOKrC+
UTbUYTCYM8VbT72lHYnXS70sKzp0NHcFB7WODlHG13tnU4vDOE5AVfdl1O3CNFWJz2QtmD0Jr7Zh
oiOPtxCt+sITnyxsoQIOWU9c7CWAZ5lMIyieVg8+TnTuN8swzMDr0tYGLL6gLQUs2i6mt7l/zFDn
g7uqJ1XsRnt3nZTO1so5bC31SyIAhzVOUpFwrWak80DIKgmVSLHGbbuekRCihurZV/A1mA/kcYyW
LiBya2xSHDnTKntBt11Nn6kSSOjFG/gCV5WKRxGPQFAhaXSRZZAoXx63XGBtrmfsZlCG07vowkiG
GzdHeNHFX+a8xPYW1XmZVMisqj/lEQ8+AjTw5QG5134cbWiNSii2puGfxRYX2BwQkrRC/3l2oPug
Yo/ngnVJcxYiwjtveOFsZ4gYpi17WbeYQ/pEfo6t0HPTd0DQhBm1nrXuhPF7qv8s1bgyYRdzXKOS
7pIVXWBIHRZ8MuygqjaGbLJfeuwsmnYaMStKohYlqQCQLCiuOck3I2Kd/eCDdbtimUoct6F8HSCk
CS7a44mAEqJGZ7Hs7oxu1fO4EubHGpffsLMiqylp7hef3KNNndxNlARGgWxH2Se2LBRs/luD2/j3
T8Qbd8mf3DGP4I0IQI2h8+n71js5nc9r+y448PY469vcbDsqYAj8v/Us0ESoaDZq7yLpNLEMAd1v
KWqNr7gsFoEz3oQCM4sD8WPZd/IG+PC6EXu9JkpDBK2fE46F6tmCKho/WNuKxU7AdA2DP+y3JqkL
vsosxnAVeA1OIsgCxXjCMZsU8BcLZGChm/JdUMztnlcouwLbfUomkSF7N8NaG8XKFIusMJQewH6q
BNMDTKYWj+f1aysS0Bs23f9yFHR1f7mnsKV4xz42k73KXT8MoyrMMwm/H+chVBareOHnBZKKvihB
qu7qMDAFL4ai6+Wej8YZr/DJ7t57ytEq6ywp5rvOF1WGRm2kdOr5My1lEIFTkRtw7Erfrrtg7gWO
aMYnQ/aCUFTRtkcwBVvxLpSWQD2Xq3iVCDx2es5mHicA3rvOFe57qwDshP3UIV0EV/Bs5AgJeyII
MR6ItKtKSFEpMsMgorqE+Gg0ppIa1KUbd7ynO7YlrPGIzNeX2L04YR+R1HDV9flcdSwSkZjR5Ucr
1EmmbBs0ih09XSc1ouhvFt2QFQYK87lBiDUSlSe/Kr8CZgrp31HQOJt4mDJIzhDGvV2BTmh3x4wk
Q14LAuS9+xPNSzYrrQeaV0uM+UVezyPsQdGZOE69Xk1tPfPYUdHEmqLYXx3y3OASE/O/yig327QN
plIEffL9Pz0KycWAWufktniuAjO9OsWwKCFGNe0YEAWeB3kv/t6bsxtuap5q6XfRIazsTaHxuZWY
2BLtuZPforCaLR4eXy7GdUw93vA+NvwW5X2mD+dfeiskvs1aVcoiPGe9GV77H+9/yNy1uTtzxRUT
wutLaP+9ZhWJiTH5kEnCoL3kRvesvbJcoEIkf6A9wnxkuM+ssVy9w8rNi8bK6fN+jI9XltFnFfVB
KY6NgGtwaZMIHMNX2p9txA14yuU3SWQyfCv/Rgff4eejlwiLya9rVrMbb1pE1rQIp1SXLn82svOX
ihtR+IwdEg5TLldSeihycb52yCYOoK3Tgvu5wRSyu5VQTykD5nvHz9Z9MppUcCG0cNw7ot/VMeDe
GU+mwipxScneEYfarGXLgU17JM7FOXE0mUiyP7zAQiKItfpoedJfTqLE/aAtTW4vBTPQjPJtRKgM
zfhsvfLgxCn+bZ+xTykGT/0bLit13P+xP72BlKHh4zuCJ1YGJzbackX0DIfk297Jae7OBD52I52S
i0D3feFb3cvef3OaUitFsErkpQr4ybXCyE5mSU+PZiyS73wN1K6ZtZ+8EFFsYjI85mOygIrDVo9p
Y3kXEeC3tBGeuduHC/hXI5KLmm5FuBPCiZ2MSQ+btxUJ0mTz1tgKye+fo16Juq/i3576hX0eiFmG
c2HRYbqME+Fc8oWTVdi2kCsFpQZ0VSd5WHrm2tdx91uKjaO9r/HigHRAng56X4/ijLYpwE4pFmIK
6T09L8Tg/iyFLFK43xRXftSBQ3ymUQv0ajDaj/Cb8yQOSPuQKbyXobHb4mXjlDYPb03KUSmzItdx
m65xv8uwhmzuEFVKXsn00UT6ty8+EawXP2+TiTOykB2aKpTAfp2cKv+4lRMHiw7dWd0PzbMmPWBz
TMq5Uzc/WIXUwN8NTIWWsVTLKmesRpJYV6Q7uqeJUL/cQcVCFHINmgfs79Eqcps3vjU8+RNQCCsp
PybACpmgfhNeobHThXw7FbmdXZKv8mywiWSL0iTJJefjnH6XyvDeCMqF3n1zcjbz1V7ux9OVgZ1o
jHeXE/6zh1I70hn8xBkDVwxGxbO2+2E+L9tFB+P2qXgJ12je5CM44EuVy3/VFT0Pd29Lf+vNo4Sh
QfNCifVLDiQHjpPTbihBlOuJh+gO6tsJ21N99pQSfg7z2sjwTGFFUqBx7exKVvhVt9VJREO5OUMa
baskT2QdTnjUeLBBnGIXioEvwXMJstWi0G8bAf0L5cuS4carz1KC8WvJLP8uyq0YBwHgTws9BTCg
2uu24LFmLYIh2OcOTXSoc8gBZ4OANbgHnSXmTDvJ/G7zUYtUB+PnRbznC0CVH+/WrpJgv2M80zUc
3qeQNMvM83ezIIsYRiUgQz7TYz8O6Ssz/0kdOz6q1a5vSOJd4sKsGtziGVp967T0wplrcbadVVcl
wX6LpXa6uJSXvT4x244l2UHjL7W1m7O0ZcsiOpYNF/mjYXDhTbavo3IokPNuWgMaTuVrtTc+ABCO
4RaC37IyftWSOR4Vx2ga+2Qj00zH1sQ237ZpMZA1sXw+JgbDw3qvTZtjA77PP+bUXo9JHUXoQ5ko
rbsxvgfMDQGK36L2ZU5sbl6+W/hZnvrk3DfC39ifomkhhuiosndCvyAa49NynsegWYz5wC0OKkb7
3pMCGZg/AUNsBQWCVxMipJaGJLBCBBxopEYRd26z8enwWBULbIp5iwLSbg5O8CGZz5TDkZbsPPLY
AoSFCK7vOsR/cVNOtAA3zq0AoxYFqN/rHQs88XdS1HXlsnZ+b2sku90xj2ylhD0yyt+7jBThyTJl
uJzrzfgk8d797TgLjoIHgnmfpPLgiGj9eOpo8qNucJOzzqXe/20lGU3sHBeM08DVW1ASLE9T5G7n
tKdBAiJRlVX/62kWe3cEIMg6j70mdmuvrOIEd6WZ5+dAGysaIVK+kQLC+662wZqcNxS+lCRoNvwd
KeHcwQUlsyIwi2uQVYsDxWMcFTTloGBPAVfYZqhN7TAvsbf5c5pY8ddMpgG4SBFUzE9ZAnqNQ5rE
55wf5ufsRUj9eLexaTp3MHe9RgOJyKOj3hBnGQFjPcNmar9thaZErThakxOUE371FNstF1UGjVjw
WuguPo0VQz9YIve+65DNk4v++dzuKev4Z2BWimyOTRMNRaKu82OK9rxa+WYI4JZXKI/r+USDbTxT
fP2YATu/aczhyfNrpUqNVybh+q7CYYuZpI18kTVHMFd/HAwBBrK164sO7/a5k+DxCML4+UERLLo/
YXGWSM7UbnIN8QGaH2HYdENe3BOs9Rt5jWU+zN/Oy7rNC48BLwE/fYfK1c0TKMqnMNo4CZGKg/ky
R23Kip/Ug813xfjNEBTCt/KVu/xztr7y+4n1gGZbrZ1K5GJrQrWKEbgWDbZg2E2sFi6t5RO0xypV
nnbw+FHCz/eWXvkjGKiU4KkaC8zd7yokU65nohZvY0R/k7+IJf0bgqgjxWjtqGpAUi3RcnmoZPNm
9EZsCzTKQaW0Z2YctHxpPpFlycXqlGMKIo5CGhCSgeHPe4b6CbErn5WncBqBNAQYDoiZrT3zxRzA
knQC1moTkzSiFy8U48rxIHBboWJV+uu4UeGv5riKBT7XlknG47ktyWlgiD7NCfdv3XLqrnLpppZt
ohTbS/DeH/ME4wFIMBG0lnAmpojjEA+kQgCrCkx+/iD4/TleCj52Zic5GqcgfUrotkVh8WGWHMUm
vDgjF0x0d8CvHTv7Lf5NVwVcUcp8+K3muDBnAiXeyosWntVKjI+G0PZAtGPsRNTd3kOt1zczGbKY
6wiCGUs5J2k1sK3p8U9cxNl0Qafr9mO6l40xCqRS75HidVqVjPYfD79FjKZp5YVqN//RG6IKmAfA
PvaSfkmqnhJHr3KJpexdowwwhoQkqWEfTG0m84mWMdJkR5h3FCMCmus+Wcw6HlJUQsQGkRzKGUL0
O03NX+g+7NvtPE6rlEVYTjNmq1lHDRzdlM7h5FOSjbZ+zvxSCraZR2g3B4ilX8/uHnGVEJoZENer
wREWXYNfnmLkpQVH20qDqj7WhOuwIYmMS7MXU7qsNnHQBATd6Gs21H0OYHPAZXxeT0fqFL/+JMii
B6VmDlw1u+leg/w1IM4hPbXv4EDS4+lqXEvAfFHDf01kssFlLtYwghrc2iyOIH0c5GmCYGPlZZDy
wJnY+xQtkzjECysli4DVkw0VxZoTlZTKSCX5YqF5IRykNf4yGAoSWZQc6qwkIyJEjeN7EArIkP4M
HXOjeUAtosMnnV7Sh8BcW9fKrWJnufREA2yGevCuS+HQs22Bd7wbVF7u41lZaBRODpf6jO+VNGXB
Ls8KYYT9lv1QomXIae/UhyubhtG1/KuC8ZLgazRR2DSgNYDCcoJ2U755Mty7gpOB0IcqH8dA4eRN
cO8906Yzif9wX/Mn0bzTDkBM0TP8KgeNrhWVqYB5Lv3SvUMqXgLKVYE1JDF9JGmCoXXe4pqjASNp
HEEatOO8TGqMszXTQRTKZNXei0B2CBr5oD0MKBr6mM8KlIX2hAr+qEqcdme1587DoYU+hAaOB7a8
U4Waqri5DttzofpNbLdfnDJa/3VSIWJ0257GvLlVtZ4quBrNjogtyvSikNFQePVzlYEwMO8C2y2m
cWyUw/DlCE1t7XbG0aBYahiSDYUU5W87b03omYIlFucSrZ57O19WkL8m2o+ffzOGm8Wo/HoS9jZ5
1wTu1mpBt5tGfBjkoErHn4BHeRz9G4sM2Ui0wVgfTMEl9UkQCtf/pLZIjwb0Vl8Cgl7pJvYfzDM+
Qttl8wYRdKtxFVc0K2A6tjgP1tkxRRoMLP7n2FfBGTK0mPFlyOaQL2/RAq838K7SleCGzcGnsWB2
zK4DyFdSOePcRb6KRD1429TUqDzxmkbkGal+c+KP7pS9kmM8072zP3S1oY26Xfft2iOU3qjAzF7p
S1pZwz5n2lbzxS3SwCpMdGKvgR7agwWogFL8K/fCQblZtKl8Yw6jfedayGpXpTU79z/EEG+nWfSW
MM6Jnz9VWZ77qoVV1zVZTw6cXWi0hzIIMkU6tzDG3Jd0ZY0K8QGezDOxsI1F5qQvN3ZsT9/S1t9e
SrZN0TLUe3iQj9sO+COvFqM3dqcRwkBCkWgLDXXbByJrytYvBupRriUyoFHJhgukGG7fHg/TUzpG
Iph2jX8zL3BTnHEmcEP6GuVHfWFqNv9pvjslGOu0vcCLFD0BrjkVYd9kk4oNRRAPMzPJJZYqpLRv
mIGpwHUxfIwS4O49FOY6Tq1WXGM8yO7wccuozBL/II1JA3IzEo7XBNzw3YkV/Ws5wPP6pKnXHvOv
v7tpfHgAOJlzqrOEF0SHubFbXc9YNKePBmjAFrVPm/HkDR9fmagZQBFdopENu2hB583LU7Nwq2PI
b6bphOGQ2cBpur1GV3sjDBwnQWRF2Rqkry0xwZ7mPpHOXemY3rvmS89QKEhV0ljzvkH0HBIf/Ytp
Ez5MLT/MCT/LURidv+MzQixggW4xc8l9Oua95kT70i+OQu2c9i+Knmgh98shG7tSC0Dr6bZjSmKi
VvwQXE+4b7VcLe/BoQky87XvkKCGmHe7CAAzVX6QqC+Adaa1By3norIFZY3cAIkastPV7tomE6k3
b6VexZ9xn2sj/Cp71OGnRYa+PWWde8bZeRBTfYpoLiot6e7nD3Lp9TZVEozRJuP2wQWwPMsztdoa
7nme/C+bfqswivR2bGDccsCaehoubLxoIOkQP9sc4BNtuVvMOinno8Op0qdyQnROKkKtC1YddeBT
UPt27FWFriZUmdbnWAwS1B2RU8pR3dTDaDrwcRlnlUvktF0PS5BcfNMHx3IEtRgzBBy1zyWFG/8T
TR87OAjPy+noeI+Sifqp4Cn70rTN6QB4MQR47rytPZ7Q2KfRLhU2abDgS9zBpid+nqlhGvWC63CK
mKKD4/Lb1J7GXUtGmpxjq/Yg/kGE+bWPiwE2JG1+p7zzK7YNZSlUQSRSk6IiptpkuW3DSmWgrlvk
X91byvamKMCKhBj7rc3TzhKx5XSMwttWJq20TecG3N0UP1vng0NOigs9niidgxO27QUby1vKNNf7
klKaPT2HQH49mJgZvSZYGUSFKQDjPPNvHCjIX2WkE8iDTa5dVqdtvlwFOIWqsB0maZ1uLLgw1IfE
SLkNh9FCps4GA+R96YiaBcuIjXAYKxzK/c7hVZ5Vy/vQ4z/0jESV1ORXPlfQfuALy9l9r/GYjCw/
Kw6J2//jDHjWELBNMBr0vIqk44mn/V65+u2lHXJjCvnmMCHLQkiS1yTD11pWqcMAmBuVwO/NiXnw
fHVO40T6zdRggd65G9pxGadQls4sHdLJmvJyem9pC1qcY6F4ae7VzbedWJHbjMR+/LuGT3EpxkOM
ERohO1F6mEjgJbPBqGCIrGHEYu0CZpxVEcTGov1IlnwwgTd0+vp9pRdgm840RvsCiR98he93pSuY
QBEmbiOUhaodva3mAtnRyJJQmfLmNHP9CoKbz2EPHRaWKu2pxKjJRKQ6pjSAtfJqbbA3anK8C4zR
HkmXJgE1ZI9h7cYzwOEr/PCCT7q2oUN3CgSd7j26HdHX/QnlsPaxTmal4eaa+covdRR1sCME1Cjd
Z3RRz6elOMIpN84AMGEFqWaRQUaNAeAw5ywc3IZiXhiEVThnHg2QRiMNqKJmcgAjkUwuOyRTygFh
pQ2FV4odsQbExH4f1xrcME99apBfbZpC3sZ8qE8JhkseIYhlbme5ZHWxpPUQD1IdKipP2JIfF3ax
myCO0UqD4jSSirCGGrl5VuOJ+yuwrhubyoW8ZlMtqhlqBuCe0ZpdaHwnlcrCsfsOYrZ2005CwF8v
lfhQB9h2K2FyHFxtuiS0gjPBVECnp73C63vOFzj7v3AEPFlfiH/ntM2g92YXrq9ncBEzqGXy0S6Y
srbZdzJxa4jkyddkt1GhQ1As+Z3sxzUr/YO5KQE1Mek0NSH9K7X5Q7m8gZKGknUKui/c6JUBevw1
WIY8u1P/YW98iDiF0ufwwn9dKJzta3QunFFIvPhiU/cZ9v2DcEoqwoWpzz3MAqZD7xBt61wsAJ5e
mcKfb5QwRgWwjWt6pAXcEzvHoR2H4nkAwwQO1IVn1Khf2G0vXY8iWN8h5F7rbMCm6k0qj2GT/al8
jEgy3Bp52bA4ZJGVE6RKrCHJHOBNUYqEXj6aSefiswoyMkqViQ5iOWtROgQJFh8DSbLSIi5Y2XZ4
j8HQLqV+5n98aHgJCoW8RGz3x2hBCIGxmaSb2887lpZM6htWODklKjApZ4l8kIXFIzdDA4JNXfOa
F44wyA84UQJOCe3fwKJGwLrrpkPT1MN8MWJUbq1Qd7lGZYO7ywgsVz15DtzhpjOo/MTpp/To9VFX
64ekuIC+buAgJisKr1BsW+eT1l52e/op/VzapT9VUAKN+cAzLDROBdv9zUNox2vBETh+xzQ4ad/l
EjfP+ljCQwpFmGxAH9Sx0IpeHLueWLtnlVMUdmoCb/UrTAtqE0D4ehynJne/eie2yKtwa5haPtlT
s2LQ86DySvvsxzITMrAcXLCn0hAWPuO/Gck8JQspfzpSq2W/8AqKacvo7sf2kR0urAjmSegDtkAf
oxRMbbX6nhY+YcPBEsnflhoxjJ6NW4tfsTF08ODppeNWmQsXocZ9lCorr9QQs3MKpBbK7kzMOeji
idaJN8LzIrvRNwdPnHol69FggzejHRTZx7WGaNCoi/DaFOU5D5rpjpNjFrLyyXXpA046l4OHxo+g
UFDVts5EH4IFykoD26Bhx3QTnVQ/kKWcc0F7sAOkpOrPXL1ZkE4Qe1WRKPzJEmpa37Dyp5HU651E
z8PU/8S+ephCvHIDXgnImOAff6dg8z+JCteAta81e2cpCqHS4hpxU4UbIHubujLRUQFH8m0Jzpyj
pxGeSeVkUmp+IxRHtgFaqMHHMNIcoeRBlZvSA3z+lw/lzm6j1hPQGB7nFfAtWusgEF65GO9yCb+S
IktCNH3iuCHCPbLXuQ4hibvRv4WbUZi2MOYwHf7C1rKMFQ8C0mQ5Y9A6EXf6JZX4p3Mar7LbmfGo
c5uD7Zw3mNiQs2eZ2VxZchv4C52aQE0JMUR3uvLd/DmtfdXMJ8o88J+0p1RoRWkfM9d7yv3zQ0Uu
2HtPDgw/3IMqfAsXkiocSFdsihxz3uItzH3hip8ggkyid1iDcWl5HxclYPCP5Qo/reUIYzeQSS8M
W0TYX0QPXLxNoWZ1++F2kJ4hhnkOGPq7CdT8yzq9KlqXX19noUtMR+yKsMZBWJF+fUJyVAPcHdC+
tiQQXCu/0JDnP2bUuZSjPDBmMhxTOumahnScSijoyBatg993i1j09NdYzbMToRzYI4qHA/Ga1bPG
HzHyl18U9sQeMGafuKnSd4TO8rVQPL+nxuQK+nQs4mhWFVXue+v6c6EHPCqHDsIbDckATi660m9r
y9LlIKr+NgRN8DvAipcFaFDoyvoo7Q6tUShVFWk0VreRtwbtK1C9AnfijV/Y9sk0uXAa3HiwMxYg
0qoMy3n393MRke2ut16A1+qQlrtF4zcvkIBpVJZiXyrvrdbFKiVjeT+PI3dPIHZJG2rwCIvbUsF3
MDkE/0UXMIlHCiF1Rp+1/LZ6t1aG/89aXR1co2JroapaiXvrcSEuJ68D/T7XRcITx0EI0IImt2B3
2UYu0+Jqfm4O2PMLpeilKJj6TAng9vrcSoaWTR/Ny37hwjJzHp7ZlPD+Bdy4zrP7Nv1G7kDkCIpX
ccI7zXiEVyK6k7M6udow82YD9cTOJ4LOROy4LjvG780M/9vB1aPDJw3AGULXYMIFqTn/C7qS5Zxy
s3riwBW0oZZ2rt8AqULCvHFdE9zvh3Tj2vkjc27YyWKdCIPhQa5Ft8oKi2ISFyo3nyglyYmF7ilr
XFNvZl310WrbWM8TnJErtQ08aXpvx4Xjteme5FwHmf/NKZofu02NdgoyJlRG9lpTAD0LRTfIDxTa
4itbsfAjlbVhPakzclzeIQDepW80EXr9SdHr2qLsbn5ez8QQBu6DIXcX4ijk/xuMu1pZZApmxSoM
ryMXTiu7yN10VPDlM++AjeY5dxQjDomqpclhoydMwP6Ef9WCJM72vQjZsiQieaKVyJ1EgYXGMA58
gev698gaAcqsba7qQGLcxczNZw73eDyuJ5zIkfXdrK58elTYeKIZmAUJTCpgSKuMvYKb0U1PU/WX
4Pw3kolpXotOoB1arssRw5iq81TGtcmjGuDz7B6MY71Fk7gmnYwGjRvvS15P6Gse2SPwA9qg1RzV
7w9UMGy8eAY1zgwfZvvClI5XB4lXR6MhzjSrXrzN4VbQwxcMzHVms5YrgSZJw5BsWSZmdNELUwB5
Mx5DE7ncsetQ42e0sjm/A1bQ4qth4H1bNnyV9eTFk+fhBpUsVorf+BndKxoJNHUIeAOiiYwHxWdc
Fvjylltp8wx8Xh46oPWBjTcYmJOpczmQt9jqB+vtL5LYO1iymcAP6VTnFSqSEBksDTxxRJRsVxat
iIu+u4kQa/y5tSgBTXkOURghkrZfOq5J1mGZP7SJc2aCg08yLh5lyqKtnuCoPrTT25lpgCaDTJdC
1+hybc7OyJrJX6jTzMfytLiYGHpVFR6S8pC1/mMnzw6DD9ASad1e7VpL/fVxV3auYCi8o4jInwEw
0mo4NdqyMM6GWDmyWoae8E3bmw/AlyYvHzlUvbVn5Po0M4VP5M2T9RxmHf1TA6DJ/7wzMldXyLqP
4Em4GAqNPnqaRJjNDfVjO16jYtOfwBniWGrHupat+hqPvUMtuSkPr2/X1natVJFCjRmAZVa/WGX6
l5542qLkNJX1G77Y/TkLDieV9VgB6GcqtjYTwSmFqYySGBogN5TM/WNb4bH+In6NTvOZzQ1eH4qp
+APCzB2Z/lqws8TPCaP6pwgiy/kkQC02VqyR+ya7x/u87pKoYWHTgX44OmGU/s/FYgI5Io1vSWZS
Ztjww4RMRjrGfTY04alnRPunVNHCmBNeYfYsZVcMF0wIQB1HRfc6a4NnWoP90+fU3tffaAIFkUcg
i5eqBU28W24mU0D+Rv17plcIo3puCwX/3SaUgDI4MC6uSBzI09/ZZvtS2x1ujW5+P+VdIAiYZNgf
TYtoiG7EryuurhFvbAGrlao9pUQS3KvMa+jTNcqONuVN/2DBTeFSaPtPCbE4KyzNjZ93T6OzyBYt
oKP0kzUzhuNtzWrgek6RDh8ngjW4/QRzTr0B2izYdtZsu3xztCM2HrYDWnFvQMnaITQftGX65v0w
aE1AkYZx3DDg6rq44qJ3JDgIGMHWuZ2Vut9Lf4yjIF2JZeCwdI5ZHpiaRccxIHwfjJHNcWgkIvKq
JUFeiGsJfwGQjDFVEgETz1nGmh3xE3hyapu/UdKMbSdnoL181I3rxe+87vUyX/1HaFseDaInGWc3
rM5tTOPNQJf8ctgRtj9rr7GdshzzB0ZSK9yDB8SExNnVOKk3Swp0hCPlgqoVsb3XzySYJEJikT48
5QjmSJ3ZbIfLI5vWSc1YYyspOENJVItFxRSHSjEQaFHGSR7x7kvag9FYm1rM9p0yur6iPXoLtDug
y5sCb7BB4aKjs9Py8ueVfz9YUQKwIc8/TIoYJNAiid53bXjXcVBWUzuu31bACdJjrP6aaP70KIJk
ZZecuzk+F0NYkwaQqIavFN2QbGKz6mRMDmWf+cw1VxBJWiwDTawm08qt3LabCQUvOhvgmIrC0O6r
REjdxyaR5g120X438nrV5W7KMpEfOBmDs/mDDaixUMMP+FoNPRjWHsGnuDOg/U1RToYLS+n9b4OI
T/Wxcd01Ljkpiu1SW5Hys/vNEsElfWngYNUz9WfPs47dAXRAGtZB6pP/cqP8kKag5K1rYswdSNM/
RbjGds130P1QSZNvOL6ljFD2TTfGK0/NF9MiiZ2vu+KGr9vIGkK/U5kM6tJPXoQeUD7m66WP+sv9
HWdkF4aZp9rLSBZZybCBG9cDvgNOnLU5BWD63T32ecy+7GR3gAPP1xayLQ0IzHMAFNMJtHYV8A37
th+T3WWUdEQ6+zRUzvVrV4tTjUZuye6O11ZKyQHF4fzGP0Kcveylp6c5pFZZ6wOk/Y6SsDMfzrWW
k+5H5axr0q+nitc3LEw3wI8CtRXU72yTqRWtFAZiM2/pt+MWacyhm1dJGrvrk1dJhxN+S2QqYL+G
/TuGGfga4ByOPb6UvtYn46tye06VgZ6Ig4v5mftsOI4CD5PW41HlfqHDrDaltrosOyHaNhWxIoUD
YmBGzGkTO2nFF1RXFUw4tX+DzrKT6cUKsa5WVIwW12SB52L2G9r6xk+cEDKdKguGCqDJamDDyQwv
5zFG985e2kpdW+WG+X90etHsuTBDnm3X9z1Kb6RqEue9BIOgIsrBxyDbKnhRm7pPcIG1o6IGG/YO
7uKE/gXU3Nf7FhCNtvClP1mMaMfP4IO6QzAV4Kf2tu7UABncs844rRwCH8YdKCe5zW5m/6sjtEEv
+F25d1BwEhJXPZmuKLfjmRSoT2X9zcDcJABCpN3NwYCKnquT2VvuyD/t94FvkAr+WorZKOx5MhPq
5rvO6LmelXFbDrM0KkdrB7kbEj6JRVuBfsETCmxe/2sEQMVlrYWcmumMdsUIk1Cz5aYa0jiQcu7H
nrk0dmRjOsopbE8/u0otg+9iFwEGTtu4RB9DEOPK4VfQoAIk9skojvcz8gVD5GBEUjCAoaohBgXI
+hg9QX1hy7csmbeh7D31CWYBjjjWIsPviUVjF/GMU9XLvQHYkmcVhIJtw8ebyXiBPZ4YNhTcDZ/T
fq6qoRKNl52zBiauTSZ9fZUB7NsUOK0AyoS42EGYzkmFpx85Mf+PSYxpma4orEylEmL1g+B30WuP
GC3KJHV6UQiIaa2poYFrMc0RxR+R/dEaZ3KM4HNZicvWY/TGG3vql2SbwKinPd8qsmcLNgdex5kB
QnRGJdT5DOa8B2mELyxErf+DTvm7fgM4GtzTrDIf2dzaYaiAiiclYtSuhVP9Yvp/Nm3UmiMUht2B
GmVwJ43Bb/DUVvbc90sROghmv20aJzsol7+LyLOHgZKiI7pTSHxOaBQJDJ2dfTZaHGhINmH4vBA6
qrOTAlLrw9CH93MEjhdN5tGW+6O8ooEaxa+5VHKvbNA8HdJfr14M84dV7beM8kChMISQwPn7kixi
gpB55jZuEzauWcgWeMXuk10R6O3rtaaug2PS/xJH7Z/WQ85fyS4u0SBM0kbq+uSvVIqfIHTpFpjd
96j60QRICXmjOpZP0ujrKP+R+KrdWqG03R74UDJfjnZ4CjjbhWxb6P4fDW+W3b15wwRSLAGPgI3m
xNPzqkqTj4QZeQZU5AfIFP447mj3x4TXu5ItTEeHFbaXhkWBdGasxrK+JZnYFDjEHKSjfa9vsP5m
oO1edvixpc/2J0yjFmhTVbeXLNPwKNN1JZX7bdCqiNIlQ0d4gxOhyYq3Wbr/fZ/KoRkH66uXyhLd
6Anw681A1OEPpON+Q4OM3jWRPnpRaWcdxyzFK8K9FccsI45aaGxdSad1uVDllLy7wxPQ60QFhM5i
zXoDLn8e52h4QwtpZlcpIL2BCpIxQZj0V7/TJ/ED+8YsYG6Oy5C3XZ7n49+1grlR2mjuon3da+je
xY5M2WDw/CqDTUrJRSvw2BT+9DbG7A//HHTqaiKJM6Q+58TZXRj48IOv9L0DZRsPOnSXkEh5kW5t
mzddjDrVmzahv/vfwvhaMyIBDxU93XT/QBET33icQQ3fkTpM44/5N0fKi+sjKbgYLzMguubgAAbc
smEYvZrVPgUz8JJzU1uS1qlQ32LwzwLlyHKu/vQ5miWTe2nLJWUwcfNJFhMxFFU3Yf3Gb4v1YBFj
9rDr98sQdyo7RM1Po+df+X3c9cbmdW79E7VRLpJajrnStOb7K8GPMBgQJ6av5/qpedVY81cWy46g
vaCwiKyr0eMBbzm4SvWUgyn+00/SfIvie1GPkRwX7O1TZaGmrIqCsOGlKcfXdB1CCk5RfzlJOCye
Pchhp9GTfclKL1mWGFmNIS/ibg7KDchytE+VbWFFXRcSSkthJz9z4QRCxXA1BsskJgaqLufw052l
YULk1NSLBTdQCqvSMteCD7OlCeErwjPFSTQlmz3cheaBHPEM5bu0Y3OppwvasBbWZNGNpibpoVfh
yFwAUZD+NSqTDljCr7js/Dwz5D2TXd8uq0/b6odmHi++a+TaSbiTSEUDU3+u4/4pJMMvMWulHaty
LyC9S4rExICAAulb8lS7+SXPMqeP1DZGv0AWUrMpWsjder4zcTDa3EaV92BU4zJDthIWN+NEkrK+
O88+NZR2HZDalHM2l0POrqTQrgSW211gJfzKvPv6AucX4Xa3ie5sY46o4/qdxK0ZQLyuKsybveGN
8Uanlq9l9S65tsOwfyIVco/AqFo4XLljVXIom3Z/rY3qiUhdm1/YwODd5taKK+xHycqgjU02aMnO
aG9xY+v4aWNejsSzDR753rAV1rhC6WCreBmONum3X80llJDVjUuViBY4M7/OiA8lZgSVsJb791fT
/CDFzAMD8iFdMHkLiHNCzFmkjdQfEg2nCv6mK2/oEnNGtBeasG9lDrbs4y/VrmkhwWUfIEp2Mm41
LK/5H0TYOSD3u9dma9bVjP9gikJ6jt4+gscHuA8mVmj68asCwG56hAT+FYyvHZ9chUWbEAKBOuFB
b+ZBl4Op7tc2FrxeaNU8QiKM1fWC1i+HMKwLtUCBYuqb9r3rU8ojzHMj6aliX0RYqPWfO76KJJ07
CNAdMfy0WlXXA5lpa30e7ajLy1eY4DETax456dthYws0X3ULg3+dOHmnodTgjtZd7CnhlthFzQ+5
ZJ3UbpHjOfpRkT/X9GP1oszcERLX4cIeKHKUIbUmJa49tIwjb5pnwvWh6EGYQLxR54EeR1Xnwbwb
Dcy3wdhJZZpC9cc56cZSuL02JFeLcVGas1NWZluiLe9tyAdnmPgHmWr6E0ckYev3W3chE041JFak
tTToGbiV9CqhfEY/0GaIUVWb+gr4ARnq4z6n5i4fISVdyU3E8ROhXvJ0dtQJe5ttd5f5PLEQSp0i
XXLbPqDj0xeyHEDGPHmqVWQfn/m+A8VGX7KnBWRJeWiW6y88KzYzotdyUJokvlVqOdclZrarDNLB
8G1oaNYRkPL6Y9t/y0qmSN1AimAu6qFahE6cqwv64cq1Rrux0sL0ERQKHjO4sCsvJSBH0TjIZzuT
RNwOeNAs0joGtCVxd8YPstPNl7SW9FhooXpG1U3f22VJJ8hPnO9FjeoYqiuADRZ20nCkjtj113eu
o7zTrUii7xASFB85DTjEZX/iOEBRopgnknPbKId8Kx10gO2Hs/aPcU72nIliaydCxOBpAgR505W4
8KRXrAJTMjsx4v+UEgf05073o8QTckQN56wvk/jneRTdLYg85D86TW1VYKCUbTg3gd69S7IifD8P
vQErhGeT9KfS3K4pZmfMxmkNRMV5LrmGhdnKc6G/KOs4dmINzCGyvWSyf8KScB5ihNJcGj7CYddl
3314cHvPJgMEBws1u6qfJnKyTkhkwjvP1LLsqdjNgiPCEU1YiwQBuvep2Vm3pVnZIH0nTA2LTNbP
suoiA5NGdXqF+J5D7x3RxKyLOYCERLkYgZLADttNUBaULnpQ+I3nfgSqFmJqdVgvlFg7bj9eS9wR
zGRK9k6wHLxFV0oAmc1Mc+I/z1XZM+LzHxCHsrYPa6cDT3jrYwB6cqxiY3JWY5jM7ANErTqXDxor
DGWeNqYGWDPerakN1aJ0LHrPsXTR77uDukQPIg7BoFwLULr0VmEhSANnckCz4VltVgL6fMTRQkfA
ml/liPtul40r9GzDUrMrkknDSE68nB4ktuCyZXMdLuWRH9ukERrHmuGSkfM2w2A2tQPO5wRKndz3
0kZDE0I/fwk5NNOFos1UcFpG39fP7rc4b0lzxXz8OBW86EQ4QeuE68fBI4eUdP8yqXy+5+RReTm/
cLQ31837h/vVCl5N7CAwoxGl03e5hidAlTUsnb1eUOO6LwgBitPkQSL02VyqwuZzJDw22Pxs2zRC
HWYOtpy/AAsDxe6BS1Ydto3rSn/Sny3u1GeHTgtwxM8wftvJcYhV0Ibb11oKHCodSf95aHVDvthC
nI9Xd+JRxVInkYpLlixByMatmXMVQQYlxpBj0g47BIqAOoengwqaOvZm0IsXJuvWCCDZOI9w+oFT
F2b+yqV3CCnAgOJ9BUWnxfUdhi6Vmm49coSU4ICPBixqfH3Ozeq7Nyd+y10g0qvDaWXzVezVv5OO
ANLvTud3hPxgL4SjMlCBcbmF+Yl/gSZDZSO2EJd1ze376xNkrVG6NN67oyd3+6oKISXS1rHbhToC
ZOrbb0cPP6C3GR4CSTA8gOf9ZT0FDqZgE1GEjrAaej4n3W4QEPt1gNYruXadb0kZVIAKyu8DXrN7
LtqeZIjxmW55krNnvxM0jDA0U3rZug7gRmltIb8Mu8UdQMak6a6OIv/u2+1Mlx61XUFo6XzDVg4W
OUvvBWxcIjH6XG1CRPt41KEbGeQJSBWTo0XY9mfp01JwZvlxNuebLIP7LdH7ck9CjUGEx7yU8NGS
N/PwMXEkyXjQf4kC0Fr+722foSkWZjJvTDxFIbgmezhOIQHFiMJPCVKVtsSUH00DEwqt6cEGswYh
c3vg85d0aEMJVr23MwtLHJoSx/DSmk1zaPpN87jUhTBjZxEotBjPBSF5wjwIjq40XAb9GkNF3evi
cSbh/zbWlyDhpopkqQPdX4W6iH/Ti+xDA3ABO0MKYPnv1uN+WhiQmT8uFpRF4+DVSJ3BK4JT7j3E
dJ6J3Mphladzvks+MOwqDJemJEEN8OrDHAPm30pt4ngvHIPUhPpgPHfJqHE3f6JfI28Lip3Z74jr
rx8avjXDQsDaExgAAWnJe1w3Fy9/TK2Hfo3crmosbVEl2pYoJLDAAxrNAJCd006+OYGHWIDbPtOP
CfOForKE71igvkVrV5GhYeGGoYCivaWqPhgK5uMJd3SmQj3ISPYgEI1XTQXBD/BYepZzdqgb/U8T
pS+L3fLIJUoTgthsrBfPTP52tWKN0qgpr3QjNZnKN0mSeMO+SU+7rKkQGh2iOu2cN5o1S6dvvehy
4yUfZ4bbZC/kAmhfrB+/qfbp2o7L6+1OSQrL/nfkYEPvZCx06tCagHOFuT0uyZcSTuJ+GmHZiD5i
0dAAWX9CjKlZZY2u7lofbk8rdUpQt6fe9pa9qbRcg8NJ1S0k9hpyk3Mt+86kyCUPhXdJ2HBkJGzy
1rpEz0duLFEcMkQtQH0PlTKx6XmrNPcUQ2fqNSR4cpSTHLGGWyYqPmjS41DGfh4pQsGAncaQEhM7
isZvO8bmhSWcT8pOjEaJ0R0snb+y9jFwije9rcXEt9ay1qgGb+XZ/LiYleZs5uoltQ/ci4TVAH/Y
uU8F3aYPUKFcDJDZ0pnNNnbQCkvfScVGbXeFrqPSRts/BtRemBgHepqh4FgD34ZcVZRjOMkVyxJW
vC94TEc/spykW+RLXgLFHMNUTcWbXbTkYngErUgtKV28Pbi71SQ4qIdw8OrQC6lEcDNuIglTZb1o
4LE8OPGPuLgEGuATI+zpZ4wiGFq9HG5QosISBMuklMv2QSGuwHmKVLaY8tlgFgzudS3S6AVh6OJz
zInus0vqKoJrZ1awSTRY2nuwE5SwolZ+k7X37D1S24PMFB1PlfbU0VT+UXpNzWXPVuUTSfck9SeA
2FKUiZjfqPZdEKnnlIzpG/Cjj4qlVdf2fRrUm8DUVo2cUVPLd6QyGPtx8nyUsNIVS7K9sABVT+0J
ZENPo3A5UBWUa6ZZzsfEdMyuKIPRASETlhMh5/72qf5RkCUaki66IDN3X4rjrclIhoGddw8kFwqg
spAssJBAz5UVBeCzwMGKECuV+VVilHctCtnFq6Gv35G37iN6xK6M1xMUavp/1loKFUDz119cJgVn
kzGvnxRtGEFh3QuZnl/MQOHiQc//Fr6h3Eou//mJ+yFi1Zf/r5iXGbcEwDzZ7JPwLbEOlgjOTXHA
T2fcqVIVwzguW+ASrySygDU1Vguw5/jSid/MCwRu4eOey4gPifzYysTZbPlfmXmfkbtWUThdNFDA
xA+qYU33WhIBAaQntHyKSefHHhYnww0U7MvGdzse6hICK0G051gaU0fx3FapnowgrDS9nwn+UDSy
fZGD3tfGm2m4jbZzkCGvxDaR7b5DbpT7SToryqjZcEu4a196zeFBLeA9RVOOfcuI/2SRTWrn4S9v
177aLPody2SKg02IlMFnnZHfoniqI2/8T0OTITYHHrTS8d1H+mhXXkL+loOdFJ2+pfulrIOmYdpE
QV1PovW0vl6z6d9YC5XcG4a+qWRW3x2Oa8eXYG4UZj7zSM92RUexKqLmJZodwMcWD/jM1j5a1vv8
6Fyj4kr4mSJe1S3RZ4BeLIWsDrcfCKfxOzqkEuFVw0iGWRd9pkQNZksQjmg4cP31W3imYTD6uMCb
ypFOfSsX64JB39J4HKlCKDi5UM8u5HrBDn87P8TCDu0G+8sWVhlavJcUW+/qxYGh717LsbnuIMEe
73WKIFHh5m/piSg42HfR9fL8EuNZJ5fDxMQE6cicoKYI/XIMzFw/NbjXsiuqkhncT8GLeJ8zVcUP
SF1en+A+cowkKEtf7GPmzCwnsMSJI4KXv6R7KNgZpjUNhcWH7OsVQqK+WA31VBaO9VH+CawHQ/hM
5ME/vNO2lCXo19fiT4f1XSSkX9OSrMWu1GXbts2FMH+YEmzd0lA4SYrLE62OV5nX2QivgDixCekN
rdOij+mYLW/2V76v9a5a7HHJyiKTHSNoi8SvPIqcPU3Iblvs3zwkH3BnywuNQmWvwUNrBFgi9Jqj
axj3+ru12W7cRz68zj59vmD3RHxRtFDuyBgujlFMXB0zGsICZKMBfpQaiWQuH4UkLUL0g4rC27D3
envDzu0YBfCw5kdqjjPhS/grqNnT/Co7FApSajtaxaqdnU2G81CvbBrKvlvzBU2QRAHeyrqkFpYN
alm5vNrUEd6gs1cGTGAFPIYS0D5XytNuzE7Nx0ru4c8uaiv0mUvN7zgUWuDRBwVnnU08CVflJuQ8
Oq4I7AHWwFcypGhyUjH2ayEQsI/NOfgcIUmMKGbgK4UIleEQy/BbC3tHbImJlEZu5A1qIEks3r+3
HHFsXDtMWvNoGaOcmstL2J3KQYgOxk0Mm462jivWWsB3iu7wnFj8gnmeQ45QRKX3UBAKB6oNB5UQ
4VI9JBRsoAqrJvbB+HeLLA/O2m0i2+T8cVy1kwRmTxvGd9c+N4hNBt0HlZBzkWDaBslCKAO5kiOZ
7ai7A7wUUHFhBEGE0P4o7GH9v/Z/L6DUAzluvs9favVW/0TBWi9E0Zcv7rkGe+0y7ZKBdJ4BdOiH
LqCTwghvexHK0eIUvrLl2uyNSfmu9l1n+E+bD+YSyVSaO+zoEJ+55nYTRHa8Nx5E9WsmcVD3srGZ
O8HGEmtH/1fDY2l7emDtUvSVJP4llmxmbG5GWBRZJUhJD/gzXkoeGnDTvnzBEppOPW4hhWkkyDuS
Bg92niJznN+NWB9LF63BxRWyFLo/KDj/uecwwVbbQKeTlsFbAzNGT6FCfcDs4XPJRIp6a+9DPG0J
vQzYubWuYB4fZhRqQE3xQv6vo9pirLKY9jlOGD7dVFDDb0gT4baleTW+HrDa+gCQypUGhzXxxdvE
CU3/t1ReO0dZnjK4gKHoSwvyBOMqvde6V50NVJIybhg7QlOzZhpV80+1/GjtpcD7Z8ddrNMHqNnu
HjaYPQ8kPsL3a7vM2Nj+TrATnWiUHmY2uTzkuliNeFwHZwFEKiD/F2V2qC5+ccabT3HDncqXGwCW
nyPwMhYVa7AsNGiE4HCPjtbrgpHGBrtlsTfGsOWsOAQTzRgOJi+6Px9gtTqHH2tl3+y8dbVAuaNA
81HpVltRVfz3K7YXCUnOCCAJxDsnf72fj6qi8hLImuZC2n8KZAkIcLYqdQWsSdb1KaD3SL2i2Hoj
ZOepnu0QwX0kym0NU85EVhQfEzndmeuOoxyuD409HTnZxO2O2+ekwCKx7JeCjtGOokG9aBF7xegQ
3mN2O1MdVP6aJ0dDB2Aw/axoxjEbpYuWGjvsOc4rROfCpmKQuLfHOGkd58tQPa7Hcd2Nzro60dmJ
1xq8vLKkH3vxYde6NwS5bKXhLOJgls7GMggrame9t5xt5sCGfDGRPlnZkwBTwZCBGerA9fDoiqtX
7Vb9OOTzBFmfdrnfCiH2mVHbZFbA9D0hjHtsfHRAgR9FVQ6lp68dvOZprCggG5HPlPf1LLEJBgrT
7jsxBNF88kGKENlzD3KAHwNHCu/atLJscixW5e6s3Nj/apAPP5KAdxC8rHYnDkX6s02JiiWrwTvn
qqnNUvxnK9X5AAMdK1w+stdLy7g/DqLAJeTJTPBKW3Xw1ocWNbkrx5wK6w8f3aHuIIWmzLufgJYV
YjyT8qfBYSi6d8ndtE6QWivTGTI3gWTOWtCPD9fJIdDc1q3VkgjcdRefQQkEcEjxSHDnW9oGwcHR
Ra/OJVx9rWLb7ewGi3QGCsqgj2UmvBLWGeSAq/xeKU16OpO5oqWdO7oioMVgR43GWZOvDBCnjXpO
jsCE5dtl32of7d/3h/V4k+28M4D9Ojk0RlVxFTL/YnSVdZ6XYAJdkao8ll1DecoJBt65ZF2Bdwpw
B3KLQvLrgwbMvgU+bs5BfiS3QcWkaT1259lCv0heDh5os2CbR3eJncI8nQZ6V9pnX2SGtnakQRwj
86aNxgVfpZMCCtJP/8MxTySlIIQ1XozhbplTnR08DvPr0ehzyYp0gGP97pGrRUa51C9urKJtl4cg
erUo4UUUYiACiQrjyDoOjx4teaNj9LR94YDv5R66DGZSK/oLvyjcay5+rrW9NwDvKQ1xVABQR8yL
bRGIwE1IRI1k9hIjigqdaSmlfPG8WE1KzNbyn88kPKAV3AanCizRD/KKBpr3jzLyqD2nTk6cmgeA
6bm4Jy9Kpp/BveWORSdze+fsLki+NA2ymsxThkzmdwU0bCY0zFhj/1AGlpcOE1N2EpQHvsWfQrxN
zexC2UtCNrXMwgBkxHemSEROYROzP8Mk349+gM/4H/6RXU3uVfU/WWFCG2J5ipz+zLjTVWGj0CnI
VRXLZkz1gvnkSZyw6eMYv0q01iG5Kzg1wlLzyMtYxGF4HHrAHw84NMxhgXHi2todQfAhCgMPxSRY
K3FhUkK/zQKtSEt34BtprMsNYkcqnJ66ICj9/TqQGzUx6PZsWR1bfiMIa/LWr19cnagewrLg5CkC
hx0p9RThfk/6dU6LjnZ8er7yAhdpbP/khFUq8rSZSs/ndbN8WosXbVt3NU+cxtjy/BW0dAjAWH3n
yocLoFNWf/UXuJ+OI5bUHRBF/qgU5F99LtBVBWy5TLCHVSVS0JJplYrGCGHvIH+bRGNyyjxtAseN
jzWumT8FGEf3QMRIFqNkjg2pPXi0/XoV0Jmx8y8GOPBqCvKkPsg+5rSTEGAbJe0B47xQRnf26g/+
REXCX45EBr+hPAIQdRTtRMTBMP3H9MX+OLffjDNYj9YFRjXX3+zEtK3mcbByXOWOvO1kD3lQOOYR
uAYk4nw66UDSARZGMJPjKkO5BijBhXP0k5/TDOcUWL7O+mo4uptv2Jl7wYtT9tYsuCeutJe41iI7
6GiEnZ16PmTObJtotMI4m4xdl3FPLDqfi50x/YlyfmxBfAAAsMBSySmPscGSSjPmFB/03vuKuSEY
TFlDKjg7vFbwDTW3KtKOScRAi51amq5nfmQCoy8TjXNtlhDXTEMDN4KjYa311D9jcxXydhqQ8rnm
GG/mFjYRWdlH37mY6aXo4oyWX4Fe9zE51c9iLc36VVXuwJXb5Y2eQ9d1JFOJjvIhumWFUX8VrscF
w46Sm04OoPuogBBjJio+czDHHPSrTGDpTvvWjoB4i8oKApEG/9rmIaPc6UDjiq2Dw3bSqS+fis8l
QnCdjbl1p1yhM+PREfBKKrWmZJGEF7O9WLqDk96GdE1D7Cs9mVGovtRPwqFIU4109XF5nUK0YO0M
b40oijgi2bbNtTcHGDZWJ6I7sGlEIS2oHxrX/wr+3mm6gLLp0JAaLwFIdVzecB+4SVe4sI1epPl4
ITQKWb5u6Q+QfYlW6UpSVVpT/MJ3L7t0yNp1P8A+qjZ7v/HNhiHtoj2JQPF+vkWEvXaw+DBA0lVR
UnE1YeSjdCfxh/kDEMsO+o6qqfHcVjnY82do0stF5ycvI3G5mA0X4frw+2ldnDmNc6N8JuFUn9xa
iH6Au2IJkRrcZKgDM68NTzayEPTJLGWJGj5F1rXcHaWgJfPTehVkrx7I31GpDe5ASRrHTNfBkjDm
JwNimRkk/Zuk9KJMRdv9Lc6UxBCE1DMILLKgg2wYqYCqwsxmBVuKKEJzKIgVitviHcXBZN/fjqx3
Jg3o7/1UopQLspz4iAIiqLO174H0IPCS0gpMdLHc4iSmh5oNRj64YqQpvDsaHz/uibchQcV9w7mE
EfqwPhXU8bpEzrFBISUAYUF2FgO3+iQyMx3zX4QkciSD8b6gcSS7zq18pkCPCYDTF9Yn+wJDYCc4
n0QCel4u5Pj+1tPHSJLx80oJZyQUIxj30Cwdrew28HGycb1I4MfS1iUo9otw8NgFoxQgwu74Ydyi
J/fd5Nq04hH5fB2zOd+KP+8mP/bLWMSaaN14x+/QGkyFK7misFoVxbjOaD7EiTQRpuhx04VJXlKQ
lVtds6Av+EMkcgLFENLh0VhyMlpDCerV+2Gj7DTq9K9/sqz+v9Kpe27MJXe99SGnlJ1O/5pp5sUe
EFh5w+oOj7Y+cIjnCRQXb9xAbS36cMsgdAT/7IIa9A8lm84pq3KwqH2W2KeP/5exziN9FZdxspWf
5D/HTahIF8Fy4rDMCyzf3jlXV9ETsXsd1ydtoYB9to6xzLtbWGQMRgUVlykEhGnF24R4yOwbOlvk
5jb3S80MUSoS+16GIBQTs6s7LKxGivg6riIdwnVWYJDPs0eNJEP+fX/Ynm5uxNKRHNGh2AISZsO8
15VTYZu1YsSkkkkhEF77gdTMyMqPuIjd/eXJI8uTslwWYrk3N33iar+xUiR5NpnJhDPxdpu0VTzI
bizpYfQS/82qNjXWCw4wIjHy3GPLH8PFOeycvcEFxiak70Ugjc0ZUXt1NUYns5VTxnlcdvoe/XuF
JyUTBwlYcL9o5xHFjeXbwHoJbaq1CHqGL04PiEVobGyhkSHqzwSXAbkzydDjccl1kH3w6CbWw9Py
fZyhVHcflBr4AYhLvrZ3EjnJDCYb3CSRrkr8oMijHG7c1DC6mXcRVvOD+LLGseli6r+eMH4IzR2i
wfiq6gB/2KZBEsJerzm+4kex2KgXzwyeiCPhTQqhRC1x5pmeawq31DxGurKWjG9a5oA8/SL922aV
wnJOioP7OM0sleQXdcEjXl6U2rwcliyfGzwpiIjvkntWAz7c8yMRHflpmWOYbEqYuk2uf+w0MogX
lZuA6G8ffu5A4IqjXa9LDDe+Y09XF2iLyiXxF97aksmDyL8+Lu3o5M1WFUNJJLWpFbx1L0lpLJtc
31gFxHkJKbywQ/8sBnuq/IkEcyv8l8DYIwgvW9z0Q+LqTMNGrDgYlXCKzYWnS/PQz2g9X/JQLrJD
HxjZzvNY6VWfV32Q4toVmUGKgpczF+nEHcABiHXyRBvb4+hkLo5piC/HFoRuIj+yoQYcQt+aaujQ
Vbx7+oxujyY+b+4ZQUzDE4an4N1NTWj6kktdmpNxHpu1qpGqxHlcKhpXkNSfkr1Gx2GCOFiq3qgs
asMCWTp4BB+uThutSjXh6PZ5YZmkfU+HL2LTU4sZlWdPHAgtYxHAx4yGzlbZp4XH5GoXiJUyEOPg
92vsBJ6dohad+rwn4jvY5SxWIDKDFL9jRObHwd8PhpfC1P8D2NTdPHs7XXd2S8gLJDVWEpyqa0p7
rzDfQajjireySLOUuxRIQNZs5czBedtusUpWR+kNjKKNY3hmIt3F9QMIOijN02qLoT1wrPKbf5cY
ZdkA8A+QWGAnwVk9N7cM21mnYPSdkhpZz71589OO9lg0kRfvhpfEWkdza6umnzMnk+FhPif5JBMk
arKi3rGpH8njrhdIjGTiCoHNjxQX2NHZtjVni0cMo47pmPTr4wGWmgvUle5mv6YRO/cXx+RtJy4L
ifu7ZKhiMrqMrVObO8JrcRDsgfMp2rZTsjim95J4sRG/LmndBI0EcjCIZ7Q6OhzdNP4+SujJjurL
KNu1u0QprDC+Lh2mjjV3yT4hxu/cSQPGuq1zFpC2lkHsDeP71Ml9noxuyJF/Q/mO8Ae6GUK7Suux
8iBBXoILKAVpvX4mhnqdijznyHcgXHxNUrYKh1mmjGedJ146T1963AmhodlwFwcH/wT9EOdD1XMm
Ja2/XlOhHdDoSGgzAFgbwOJ7hwPU0p+3bO4USipQCR+cw4Jmdsh3JKSevDJZg5Z9TC0pmj6zjOrc
0QsdHTDaoITVjiZXhHAqVC3JEAZardV5Z076LOj5MU63zJany5xKZhzJRW+TQL7jfpmzGFHi3Y2G
sEGVV0KQmVHUBL27RusgXJmIuIHQyu0PDmKkZ6b/fusFeGjlaPC+As/C5PkAqaimsa3dvOP0Cp0D
PbZCVuGOHyFVw0u9v6KchI8cIWT7XK/uBVpqdQkyi7/7IuwQIIBgYczzE3qdwq942q9DLvpafxGO
kQ+H97aY4nAqGFSp67+B1mwZcc1r+CyxfQOs6eYh9d7Jc3vrA6exJ4pvUJFbjdidjCakz+YZuehB
oiZPQ/EiQhxpbBGNM9bNX+hfnbpjzhkVb3lZQwslCxVPV5yhOopMDOSz2nZv1WCYp2peqxVMhlZb
Ar6cNjWT5Ze4muVl91+iX/IT56CGqZIge7ijBSZR7G+NQKOkyHJuPlmZlIfV6BVQd3ikzD1BHSN6
4yXTCPt7JtfIj0utUbCkw60Ft47FWBmT1lnfRQVAbb8BK+4Q2plvoLF9i4UWYSp3Sr3X1nqFLxIE
ZuMmPdUWfLrFOAyQq+2nQefgUNyECKjx0N1wndjot8WGNqFYWdGX+FN7qdTCwRfTsYRQajyZK0B0
Iox2j80hsAjFgDXvlu9JlEPJPvFrATZpy6KU2Dbp4ESAD5aIouKco5/r9B9cnFnQPALT9JoYIL58
odUMx5UETtOE3r0e+WMd8DZcYa35ikkN1lF+zFhu5y26OoYq2rshZRqEnt1t7qk0oMZsrSJKObSd
Lgak0xLvpmuI8WCrPTKFarCacpV0IaPHRcEHmHT+RrL4kSxiVdjgu4P5yJ1oNq5FdRBuO0jG68v8
eXc+GYSKBwTPE5rChTulj6Mgr70Ytvo9WVUC00Xk/3CpSowHql9cO6QKvhui714aD+nge1ZgMG9O
JMj3Lf8JXGCHBUIkb3Zwv/ICir7bbUgiGMlInED8oX1/6DOhENuzYvlsVZkigmgUBbBmAh3REVVG
udqtview+EvBSLQK0vUp1H8svqbaAh34IeiqAznXVemPwrPCWSThtGyZ4z0/cn/uBovQho3LOT+3
XZlaPD0s6IGLeqVLVmmXq0VDNbJ47YTWFtqs+FYhAxecGxECmcxDosp5Ob7qdNOUxGjQ3Q2p58uA
Ppbre3rpmEL7fukpKrU1YDvhnE85x+rHMc8uIgyk3wDEHarvDwen3ncvTP64o2ZGfq15j+ZrdaPP
NFuIkqLVq+rXSJgBzTPVaVQ1xrlDzmyA+5F9hfASEjtO+niYeVWKDJdpR4bSS5Z73GO76hr/F9qO
H9AmU6wDmUDFViPvgVqZ8+yeAA7lOg/DZEYb5eg6tsMvSAzqMCMZASrRCE+dBQ3GdIn1i2qd7/NU
crVdfEIKfSDUmjeaguAFhpNFS0KlwMSQsc6srDxCXddrwfLo7D9iQAQMgNFHlrrp8KZhYq9QCm4T
rNL3wYEbzQ6+TCRTjR5893yjLXIUhxlFKUTqYrr/2B46D8KSkd25eXPePLordoj6KY2r+ruAffC+
Tb+MwCEa/WfcY7g7py7FFZw6c2hTUrMOc6nkU4OshWETl7y8gtJr6G2Ut67W5Y+nvN0Z8G5r9gUg
Qf3TOM7y2HwenAj5D1q6ZfSETiPxVk/ixnJJyWbnF7wGt2G2J5FMJdVbqNNEJ3QrVbRx5LYONNCe
tOw9FcRO2N5Ed/a2QcE+wkAyNA1osW+E2GBoR78KKDYHp2AV56r8RyuAocS8pk583xRuYRm+1lJU
h2CDM5OP4hEL3/hqqNTB8mthvTRIZJ7Va0ngIFLYKki86g0avIFlRSRC/cF8FbmRYMC4xXiAZE6v
sqnkGukNLc+neky/8jah2+TQwMTeAKTt70v7AsPMyEhLCeqhFHWQ3A8RRAMTXbCcXv4/GFhC39rG
YcT3Mr4La1Iia8BMLjOXKr24mkLFbUuPVf9pCB3bKzVN7REnLWWL4qHy78CI3y5qs2Kg1s7Iv6yk
qsVoPjAMW0DnFdbCsE6w1SkwEn7DEyxDgSjRsVZ4ke2FA+BCbHHDacUrTwDvK8rZzKSvb7iWUVSA
bZGRQVOGFreUoucs1bFmIKyuErnjM6rbcgieyXkuSw7ZrvUO4gvo2do0QIn2wmOlu8yXZmj3c+ei
wN7RpNXOLhQDlEICPjK+Wnxfj+C9DtH1ufk8Oyhpkeun4XNCspp0ANcf6TM1Z4U5wEHivfdGeUuS
A137SnTpfWLaP/xsTur/eMX/r6zvuW/eMFH9Aw2XDWwDpp105ChkhSiqkEEE6Y+MxHDmyhFZLQAp
G5rKsrtvim2VStpczWY65lhnrgKPCnJy8NTXqaHBrQfFw8pjOADbEcN+uLf37dSeuAr6Xzm7zHXr
VijPTo5IWcdbvfPeyFDmWI32PDchk2yvaI757heAkaiIPQRQBWp71wFvtE8cMX8hOfHKTxvZRmty
lXxN/lglA4aR0LEBAVisVcnZ4U1G50Tk/67/7FTW5/hHFLnAMdJmsuEF2/vdKgpQMDe6IB1Nt+q0
T7I+kIdPnaYK6kWBN/Hmq+Jol9kWM42LSHF9Zrscmt0o4JV8IBYwXcVZJpxwqie1LRUKTt6dAxIA
3KMPSz74Lvt4gU4Km/33ydpNOzgPm21y2qPIvVy/QgozsXxUxB3pJ71Lwp852waEUj+VD85YJcBH
JXTcD2sX7c43KpcKojQQTYSxCcjnoVKHDt6bFijHwolW6Aptt4bGt8Xk16mF+0InzU78A5wPsuL+
9OxJWZNGBEoiL82hCSzGiCnkyFI/SewZsINpYKztKwnIM3CQVmQhbMXWDh5dUTX5/xwrFljzYRnm
tI4/dokvittSF932ImbOyTOW55FBZygFwJtFzfNT9RRQKO72Hu9IXP6/0UTo1KTG09/uJRT6tR0n
siuhMDeleCOkkvuzzEwqy43ykONqCM8kcnKCnTYGDNm/XILhSHj1+5QvZeLGOwsUO7fdKmiAt3ZF
SjFdGp0yHjQQXOj9AWYeAcLlx1hI8jzO0sXZNeYY0jobvv7NfMMIyymrw6sUdrR07EN1lDHJR3Gm
vqY93+PL23HR8fuaUYKNPM6OJlPnZhNWGsmG9H1c0zcqj8TSdQprZiYMQV7LgYvX3HxLxODTUjfK
1Hr0Gele1An3U/Z6dJ2fiXezO9RgyLRIqW3qGgz6C9S0GIZh7HGgAPHbCG/KGo+/dGzSWQaZSVrv
OMKSawlzo5JytLnSayeKGYHAg22COEGR0uWeaDCCU3hB58vX+jWL3Chx7ke9gEFEq2QNbVmyxvYX
He4xroDWzW9YgY6WsftN7qvlZkSgR7NcGZZ6APKZjQpKm5EVlog0shduXi2ED7pMYSbc4AXOKpra
rKxyKHZ6lBmB1k4lCdaPOSMxXuwKRtO7em31tlJ9LDThSL61/GcQPolIOtgYsqtOlTcRZFKkxH+j
B0hh86XQunbL9S1DB/z6EcqoQdAlnzoL1td8DoVa+4u7/Tob3xcLsbc7WGkCm+cezVG0vP1cZc1x
cIkfNoC2ykwc2dkjvh88rxC3IgO7SgNrnDcrL8NQ6AHDLV4Z4rhQKBzaStIGZJ2/0Uni9pU9jPoj
uDm0uYmeNTHzuxwkkN71TIC4xpc4UoctwtGBK5bkDEgRF99tLO7Cox83ZbJXnegP/Hh+4dNw8ial
se3siWmcRkxi1Ic+vGC6bTbY1tBQ2J6pwwd4y5yERumUWbncnyAqWI9N+s38BnwyS63XaPemFh0i
+3FGpDXcU8uE/mHHpAs1SHCcoBGxcYRRTrpTWqq4/HV8s5Bd3ShPkccCjN5kFn1ceLNQVz9r7uTv
teR72tx59SP6hUKeLhy0BYSHXqJM79Wl/uYK5lGuHMbktj23Jlc60BP8BNx0/zkN9Y6a1Tr5mskD
QfeI+Elkm6fhnc0fqfO1eNygO0IX7h3u8J0oj3+RF2tWqa+s5Cc2r4Fi96jUwzwUBX0cFa74TKvL
7ry3cBokSevFuOGHUsq06d7YppErNUZBF7eFBCZOIYh55dhgwnDakQQXNGUw/vOJ5R1feFTP8t4w
cR4D+KiMg09WUltaGQQAMYWBT1cojZsci+Eku41wQb1k3zMqm82GcTYbvIwN53klU9Gy0UlMrVdH
qS2YD6pfHGGpJhKYmulLwHiO5oUoWV2iXtN7Tgv5Jf12IUOX33ZBh2kN2MiQPdge/R9EHSVqmbmb
0z7zOBo2ihT3xPa0GavkX30xtRKIjR4GezRhjthDoXhD+YKRMzFeJtWMby04yzS6l4HVdMJ0cn7I
1BQL91Fs5wcBCFxl2UR4V4CM2nOThLjFPLesiHC39SkZB6B20dfSXGRM+YLvvFs0oXo6YfkQDsFX
uirWD73eFS00J5ktstoJ7QZERyoYfVIyEsEwKi3CJmqH7Vd3oKZmvt+NQLLEOcGfEjvjrvqh9uux
qJ+hBOvmZe0blXWAFkoZ9u9PrnNTSfV9sY7AuFoMXZxyVEzZaKD6KpSD07/cQPSJMj9CxzhxagVr
/uBBVpkGNQob6yff1JIbNP52UYFGmkzRLuQdkxPY4fhixNoa7lp2F9r8/hBq2mQ8OIbMeFMcEKaR
kWWOCy1sQHl6ErsTOnWJA9/ie2PStuHgLHtBUm6wkUm9VRtwS6yd+9RPBqgQUGX3D6YYFLD4y5R7
wMBs2RTzjTgPIkgfIdZDvehu44Z5HSgcRFXFSOH4GUPCy/T7aRA7BaKthxJaylROQW6AZAY5nejV
SZ2yq/nCrGYPNU05AQ8JB2j6wIEwrb0g6r6Tc52ASva+u4Xk265jUOmm+gTi/8lPUiywDOgWyE5Y
nm9036gmuOK4tm8frjKfMzfCl+CpWh+rQZnGdsXJ0vzWaXFbO9d5AlDlAd/kzJBkauRBlNlRLHmy
++0Gh/k6Z+HDeDLrwuhcJEIlNNgQYdG5KkIMM3NDX8Hd7vTrGV+oBj9RnaKamNTGLF0ojjaFYpzk
v64VqKv6I73gAPkvqKDUQ0KFlB801FCafiTRv4boF9Q3DXzx6yYK+DWtEwCuTnbrO7PDoNLMNeI2
hXTuaRijz9ptdQMLpObeUB1HvG5PUrgyOmbCyZ5egBdndowDoKOYo5Fc/GjOv0lfT/C3Hh4MpK0d
uI8eMwX9PXykq+z14Zu9OYX6ykTbq5CApIJsHXPnlO/NHSC9k+FTBwAUHXOS+mHPQrCyKDd44qCA
eBZH8Tz0Jq1yJ7I/tlqvlPbmR1TN1cDOeX0xMISoRrU0RkdxKAXf8TqFIaePgqCRbPkVJCjohdJe
qFQ/gQAiXPbRuJtfxUDn0VT0EDAwoAeZG4RWijIQJE0kqLEdG5jFOuPoG8EFyRyoOLw14LEXy4Zu
jCteXOLC1ecc5Bh9ZUKX0hmNT36E5ZJc1AdMHBE8wQhCN/VM1tTzQKxor6KlyUNg8Au9DMdT0eHu
twMwvONn7caevwnJjrNG4FN7G9a3qlec/oV1lE8vqV4LRb4d8GG52zu8LludSILfqGMayqIBAeSJ
IagS40AXfQGt0G6mhZ0YrcYMBtS0/h7jw50wTQigeld1hRHs5pMwodjCaYlKvXESN5eykBVHOZQV
J/sTn3Phlzmx+POE1is6SFNKl5QBcoQX8jNVs9dxh8kWMRMJu4PcV5BB65sk0XvksUnZfQ894EK9
8QfddktIh7OKRXFRM1F/hW9GijTiHjE6buXv6Xxsy/Ut6d++PeqWnRUC6lGSbdFsy1rmoDVP49Vp
HvsTEd7WbRWUkTwf1zy5A0B6YhWOe7Y8/K3vvrz+L946e/yccE41m94JbH+6BvfoYL3U7Kdf9Rn7
XsH/m4ogx9ke+cMkJIH/iFSTEVKCe12vOLfprwkKGqcqsgMjKOgR2+wYfdNqp7OE497ZsvaMhgYN
hUyvybRGOhHqFTT1O+XCtFmkMs0dG+sgGMYmVl8RsUMFP6twc6K9dZrgAg1bMxKKAk9Qm8iQKSOv
0/TJUo49mEvDJKbtzFHnPhdFb4BYDFrzWZI5mnTt3QGZ+p27awKSGY+5qUYuGlvTJpgBYRybdT7X
NecUL2koon8g+vHiyZADh1KNIvtS4YOYcRPa07fOH2GW7ZHS2wlo9LtOIzK7ISE3Y0Brd4fe7NXs
NqaTpwX7f62BSNDSzao4aQE0TELOSI6dRKueFlO6tED+f4tNoISyO9et4hnn6obuot4DegkF+vUQ
mqoSPdaSuKqWNHAmAY9XRjJZQDk1z5rT4AMp0f/U/O5zSmbSKaaI0pVruaHPgphU+bUQq/DU1E0B
vGPV/clS7Uc+akSRV/WDKAI8eDsT/SS0Tkole3ggEeqhUtNxWwNLYsvT73u9aEoUTcU9yzz1Pbnp
byEopWNKG28rjilyk3M+Uf2PoIak/c2uZHkzTqvQlyE9zRT0KJQnAXtGZmvNLICAnbGW6bBZVmiN
UEGsZOh1VK1q7+y72qlwZVZ7sRxJNRKK/lke34R/3xq7FmMB4Pad6m6zmvaWDTyWvkvG9YH+Cq0v
d1jyLN9djcbgvziO7tAa3F31qyy01hZTMDwGnZoS/8CvOTH7fWrbZSh1lsJVHVB0z9tGsxWYsvTa
NoquFoCtiW54ulqQgF9mwUWhtVvU9/VI9VpxjkNaWu2SQctnuDAE0CZtC8XMSTYdgQSKniWq7dh1
26VG4NXw/etOSZugvlgg7cX9gNOTAuPr1XJOjBugl7fRVGNygnRk3e4h0Ur6QQ7GYYQR2q36Y8/F
wf5MT+QKlPUjspxMOJ8EHHBAPdp9aYYM6jiiONWB8DdI6SiZ+dNR4ZUGpBHLNiM8hQI93ObMP3gP
I9hYjI0BeHZ5riV2BRt2EhuhW8LZGD6UugIKvQY/AacehNejtw1atzPORxpKZNmIRfxVD6dfoDMr
oOlKyG0GyLsIyemFXd4Os3xQcFtTk5jfrJaod+CmkX+zmMol6jAHhtHc4bF/174RkfhxSLHNNwIr
wboXM/yPWdlAXGxPz1m7ZHNCpr3TMHTSv7oei3uyFiWDmdwlz7O9esTYNzw6HXMkeGxS8rlRBHot
RAa7WSHmmkCZG/iJsm9p1zs1WGMMsjhPq+VbBD9xbpY713CCUZ96ULCxDnjJ/97WIBCqqD62e5C3
ayEQfA3rjHWQscRTa0pMKfYZo15PlRfS1TyVRdhixlF0OJlMBoZzVujQkMn4X2440Sjxug0DTu6g
tzj7dI2ucrcE917HDHbeNOKf+GsUHyCJ+VGV/0z8lTwI/FutkFoaCec8snm2MNbT0j7tNtQWkpfs
kvbeQHTPBQxWG4iRuU3BUdGmHN3ZJSSYi8jhvA8SPmZ+No+N20n8/Il+wHGMl+tDYRVbJ6U7QjaM
AFMAA5ktbh2nX0ri5hqlBUdN0V5PZmIQzfLaOGcIBE+JXplA7BffC3WoHmTjwvi21eFpl0PCvjUJ
APsbDdFKvi3vWVr3PIeStNa1Zi5ySddGFh2l4cE2w8TSi7d+NDaoQGYJZMFffD4tR5wD0xyaTkUD
6LCBtK/xwLX1y4p37eTASPw9sroH4k2M9GcVfcrXl/Qy9jB70t/FygOgyJ3vwKG51STPVCEJiE3s
JDF+kz66N/fEW2PsuRfktBxfAwtdhSmnRbobNtiDJyECDcSSd+rBCGy4zeO0vVLG4A50hQ+/ZFts
Lk3sq+cmYrM5VoW0Ql/Ca8U5MjslN1OtdS2j8ris+mLW5c1w1OirNocvliyCO3WWO8wxFTRYOp7T
JfWq8obS+2u1eYUQz6WuUtRdZr9nj8JWs9JUVQv5BN1xY41+DoNq1IHpa2VUNpnZcVnANlHx30BB
Xngepq3A62V1CvdciND0A+IKkK6xSoDswD9FGDRfNMgLx9N4VwUNrhkO/al4ZbtQwz4Y6RU4iTZA
qN/p5m8715PZTh5JCdNQwf9K0EBb5b5Sec71duIOd82el2HR/SGUUT7GE6qkncJFPRCEksJAwxQ8
OldQwvQW0DmqUE2dZPDX3DKrE18z0lqgKMRQ74rnNID8bGJG7Li4C3zuOPmd8rAmfbwyUH6WtJ7U
BxWvsHQ73Co96EO8VZ0hRLUlQymqVx9Klvx7tbAx94KLlOnT7BKR3Qj9GSEMX10ODKTd+6kFJ398
oRVcVljYp1wqo2M5fLhn2lHl7/blRQfwCugw6LknBUN59BWCAGq8hB1rZiSTF5Uc8QrAHzAWkCbV
3fTBg5rrrmzYjvcTEJ2vAPcTkYyX2/j/YAAMW5fRcTOtcZ86MWdrW9MpxeYXrC+Hr41F8CamvR+Q
UvmBtJwJiAcCCkXBf5eJIGXQGRmsdeJw5anrZbR4OwCI8lVd3oAGv2y+hdh1CVpzxAMZwLcfPTsf
6eABWci7OTVYeS5RuG4O4Ngj1ka++nHswaEh2mTsnbHZ1HvQ/oBUS7Wjoj5+uQoghafI4JCMgYdt
vpZjl8MDrAL4rvdk5bg96wcmzQ13Sbkmn0CWFNzt+CwndC37EKA4InhKnUyrizSIevG8MmSRRYSU
ygX08wt4qDqFoBISkIxKd/1Yvfz/gpvuULqGu9K3/KE2lppigDy9677q6SWBbAHgMW/XHYHLBdMR
yEhS7mtoM5k0CQhs4RbhWjJoJYSjU+gfIdNktaDCL9r1b8cpsDtrgpVqStUeKv566/DxeTPYih88
SjY0aF7ofb7fShnbEwn20QlIOiuMOMQttvNnNI33waSUlo99d1kL85zGyCVUV0Kd5eFBDxe1XjhM
hNDeO2pyLVCpWo+RK2ApVq+H9++B8/yovTLeZ1e5QySc6loq3HrjAOZL92yOOg2f3xB+YIkCmqSc
Qf/RdNAVedr2HRq4TiAuuayiS8hTLN3Htw9xz7YTnH0MCVckOnrTj0AsvSj7bkVgbK6z8bKNfhz0
l0Z0yJUV9Jh1f0ld+Hu8U+wba4GEix/p7QrdriU98yeMQJf9ZJRUGXmt216ZAXNsqRHebLZWbjCM
sOxK1S5+mebtCAqlHYfA+M7QQRMbudHX8CVEQzlMM2GpwRDz+owPOoqbrQV+NWh0X9jEgb6ndyu7
X7DFOu8qe+C+Zy2HHQpuz7e1szBSjghJBK4t55GenYbJJBvxqL6lhv3OSJPAiX74KDW0m0t3abd6
6U4XA5ousU/1HtHprNRFweG1qAu6422o6Bg/bUtnLqAxn1+yg8rnfrIM0PFYyM4gXPy31kbtXhpg
iKcrp9Jp3sX8+5QNcZoRkZxSgMbjnJ5n+6qHZALKKcvuHqQfOTGuYuPZ+yp+cyRS0BAf1Y13olzL
wzh2HQAGYAJ5tsuOcm74kf1k6OckLtlikr2ada3rGZNH/eiKINfh9vOour1UTvDeAkRFyQYWnir2
5RRl0wJFwOUOhRh7buGU+WQZsWotqzWttSJKm5JG1aExusKNTMUy7h2j4XZnnV0cuhwMh6q4fyWH
ct7k/gbZgpe4SAuZGMLYgrXcBtKJf0f0Vo6s7DwDmDcIUun+8qt3mdQ6iajx6bTVFu9o2GkOcbdk
2KAuTkzruzzpN8vpaDQXcAjn9jYjbMiP2NLP0qZY8xfUx3X9mGQalQy0DVDjkL4BuYYFygyB48QB
PboNhNcHnrX5VR71ol0JjVnzle8jUsKdBp7kan/Gx+Zze7Nm4hENZDt9gV7qWeeUxRXkOt4d1C+b
VuS7T2g51PZC/+UySENH4WYgXYcaNwoTg0uyL4LvI2CURuD74G9jikv9/ZY7SUjqMDIhoYKAx4rX
LaRhEoqcn1rh+RpQ4LKsku0QosOHSbgBUfqptGI5VjR9JgJnNJrmfzLS4buFj4TS8ZGrnxXzsaws
l/4ehyJYUPKbcsNSzFnqmJSDOl4XFl7PBsRUuGEPilBlxXZyC8XtZOsHtOARxCkajigKHwoNm0HY
8s/YUaZrKnjsMD5fbJRZckvq3TsU7t4YFxX4OSRuBZXF9Wc4F6Laz6WMSH8vf8bEdyZgjBxshj50
UFyQCR5yuuVhQYFEpjkrsloVs0zxWedcrdX1U+FKDe1p5suBJcux7sBZQoghs6VE+ei7Ya14O0qH
30JA9ezISqRINizNFlU5PJ6SHiNheALSBN4Z/qu9Yiwn0xfeUemuDShUOq39NBQmHc4AF71FhuV7
tsPwH0ELUGIUHq13cpGJIU4EzkyqB/CqFYC9BH5LuQaKH3Zgg3k97oPtFNwFwbRDNrqTxt3/pkTF
t5atxl0RLl4+ULm67xLI5MOiuQtqpWRbIf5Ra6nt5Wf91nuKpM6MbkWPHLakKlsH6CppTL8A8hn4
BSRbL/Eaq667H2yyBC7y0jIogiJu4fo3LI4ctlCn2zT/a0cJ77v8lwQ+rqdF69GzLT1CStGAI0La
UgfXMP/8gp4dmYVjZsa0+WIB/YnDVFoQY9KP3chju9mwpFvA00WiU1iOwxLNW41ExOE1aYp5CDAX
udWISbwQX61ZiNbNNg5y3sb8rjcuB/bkTe6KlmzEHqIEPZA2TseKr8YyS+pC81l2AjMMqaSMoxM1
9RWLdI3XmhtZl6bvHVqoX8D1avHRkKy+4I9XxYC/c3lBYkkd6HvsQpQ7YbWROvdCAd9POGiM0XAy
lwvAht0JZ8yq7rL6ogvSNIi4X0TpK/LGmzuBwf3BKxsTaaygP9IoT5JWD/COiV643YT1aBFXY462
5a961+pWBrb9ZlknPsrFQjhMJiH4n0ibdCTvYltHd0X+fSYQxa7BF1wgYLq45bmsyE+1fFtkA7gA
WTnehJKiZdx/Ch1ttvwjr8Y64PPePPz/pQ+D8N65dG1bmI1kYjPtz80/+ymEdLSuAsCTAdOWakMC
I08OOnTltHFqa+MdwlJMblPKH11utZN5+qbDy3SON/9vdEVdFNTeZmB/Gi+C38mAfL6fBNi59Pwq
frJ+wPJlDvOGvaDa4m4rBkzVTpcn8aPaZx7cl0ql0iltXzt7PXP+xQ5Q0bmageO4322I+X8AQqrp
x1q/PPH/OFHC1mvnEA5ZMaSXMJFX0lTqOPISg8uJwrp/hw1+5CNTztag4imu0jp3De53VR884RaG
IoOmQEdOeo93+0tS5OQ19p9p3W4FOwug0LA/7TRvsrGYu0P+l2bDcFZHbwIb7OdA+wvGcDJIWYVd
UDBP+xAOGALTi7PBRlBvFkIY27Kiq5NykEPm5h06uo9Kd/DSEwtBd39QBxJElEOI9BAVf1m6Sf8r
D7krfLs+vv0Aagv9ELHggubjqAqDBjJp6/JwR+FhmkcXtCOF53c6E05w5f13pvEXeRZnp8j4nhfx
4I6YFHhYovNJklMrUF3b5VeSWFBWhhPDYq8TQ+qo2LBWY01oGj+8rvcxF7qkmLray3g+UaOoRK8d
r2wXdomKVB+cnnqy0N0o+bo5oxN1EgOKuCQe59dEHHLp14iTsLrhDEybJx8I2Dky/nGNYK9xr6/C
T4QucxgHPK5H+TqRP3zmggWJFDng3nLWyDk+ivIOc3wzKr1gjk8JNQ+WHl2l9NNeTieYLZYDyFrG
hWW5NNUuDuzr+mCos082tUxhpNTKfcEQqbVa4SwxnetOEDkb0U83WZ0HYMsTS9lmgaBhBnmhf50S
MN15/p/eTQkBg25fUAdP56ysS5z4PS3eFgD4Wyixn+xZcZos+LXAcIWxamPOJfna9wm3wUMy6SGo
cdNE5qpmfiF+H+BwEYFmAhXtjN4/PkY7K+7LIxK5oWTJ1QMOvqfL31ty7uRPEiD37eps7dh7alEW
JHWUhYqcN4PUoCGqMfIPs8i9jpD88gshHQkuzSY2gO/lzV6c8NbQqJRB6Q85Lrhdzm0pUH/B2X8m
NgFypd2HfvhgnJL11XZ7XWr0/rH8o30+QMQ0PAoYs7ANKJjSmH/IiX5tJ7A1507rmWDF/NJg3LZt
ev5/lDi7OeC8d18hwev7glM6NBSL0SM1+DZ/XX60/iOGXCjNZXG4bJE/n6MhRYcHh8UcEHmEmqau
t8fVTQ7G36ItuhQazOuf0T7foW2t5eYcJo+vZl9y9W5kujKlrAxMQO6WIdvXM0AMfbo9S7hE+AzH
y4Vsr4Lb2T9/NaOnfUwjchYjfjJvETWk2Wy+TeMx+m2PNy81oOUfH2bW/7UMVsl5pZGvwLHcxmot
AuA11cReVdBL6R0WSlYPFlNGrcEVMzkhPgtcZXPuPoHF+TvLmo0AJeN0tqRnmkDEgb0LrtgTOt88
dqOVoyHduIJa10Wn0nlOONYQUthrLputRq+bQgWETVXCp6DhX70ZPFmFrlxHsJhFIk/rSOoviA10
e4StWSeUzwm5rV1EQKsjqR9ExFECgkQ0fdBBrt/UsV8Wi2WQW2R+g/Dvbn8GMbzUQB6odIqjAiFh
Maa5DYQLSAWFK5VWvt7JLGAc1uIq6wWY+vkDhqvmu/dx3exiBKrQjy67MMeLMOQsziIsklmAb4k3
Y1Ao/RS/+vNfaqpHBCD6XFoRg7gds1dnBcGV/v76sEYiL8C9r+i90KcrvvANK3WTzgqC531hkwZj
wd8I73Tb96XIw1jaUYexLDd+8u4p7YRmrCxgAQRqpJa99obAZ3tpm+Y4Pperq+TyVszbFtsfrvLW
WiwiaXBq0wl7IArrYKzYOyPC8LeHnddjVvdQpbo1MLQxpEzvtRrW70aHmOMufv9nSE6pcJvv9OLf
oNxDo7kGXUt+Qr5RqT9FHtZjopLMrKm3e/RokG1ZE33DOGXNkUG/Ol5fyrsAMkbKqT+iBEFL059J
6BzBzjPbByg6cP8uZ/u3ebfMakFceEqngTCztA51bKvEJl8xFC6yjr5+RP/Ztsn6Pcz1j63Ef0a8
HjUux1qPrzxuyqx8/C4H6EOBExSG/FLutoPw2x34Y0LWhOhhMyYzM8UXaBXMKCswhsfoydkJCkNV
TNv9qk8lifnVTnckoHbuV1Eo04fPpsTtR6MpXtWxxq/b0SY8wmWKwsl7ZBcM1rTexxXzxG4OeefU
1ILaYs/EQeZR3c0awBtAfDkFHfpY96aTPV5v3uzfEloAC+RdOOVS1WHY1+irzV8Ghaj691Vw5dTn
WObA6HF+Nw4mhJbK4Aev6b+7g290OAK6YeSz3F4EQGSScaWEvAofAKaCI7XhdhBTEMTlxXya0T2n
3cm1JersNxr64E1CEpYPORKjQEoCUoIRnUEnV3JZkR/3yT7smv0rTyJ4ft1kYyWR68XMlCrmAPqx
3IK3RldASmu/qMopK1hKxn4f4Eqz5ZIcZ7J8tiWPa3kAFInPaZGzv/0N0XRHuRTrvYtpgmGYf5Er
zMESjvTUlP6bLgiLRfNv8a9Z1t/yv9I2l7ak/ToqA3D0LG/xkXxjmbWyAbacvejR9fPiXZrwytg1
0AwiWf6sRDDkOIZ5FMkM1HOKsfynbpA8sURZkfrQWGA79bCNZZ/2ZG3XbVMcZSh+kEsdbwI4An+h
gLFC0zQBmSul+F9jhrd5Hq0MmD8GckfbslqqKgT9hFUsJH0R3SwWkPElC7Yo7fI4XKhgiDRZvCy9
yWFgnGmEB4eGUd5pSUFqtod0nyEe9yB0eK/M/wijKru2anf0j36lPZU3xy3zHCMLk4o+P5KEZqIZ
Dk47zhPO+pDDntSYWcfaLkftgUHjhX9vO8wG1xk4PTLrJhqXAgWBdI70/HHezVOlA3lc/NXc6Ty4
lZnRqR+IaM4tyxat3XIR505XwBIoRtJtkn2sw/iyZWpPHmLhThgic4C/izVcAN3I5HR99/QEysej
fYFJ/hd8YptAhYQ+gFaWsy0x8Sq/Hkb2FHruIVPi02gWlJHZ5KkhQat1YWrM1rKoBDlexIz+x9bU
8oWp8AAnh5MVfV0LfMgRYDLw6krKiOB5B7I3GcAUtXDOW8PMICvHGKkXIo+It0kqwb2ntDz54gfq
enzEjylu/18NqM/dbbKTjuBBtWwJk1fEgu8wfjsqkkXmEQHgYQzsX6eSMoLeaeEGE1fabxcnGrj0
4sTYi4LESgoEYZXLU573+JluCSrvlBEQxJShZkG/mUnrjqL5EDLW/oRLJTGyFS9pDUj1OqisI0Df
zZVOT/LhMXh9LpKDQ05wvLlJ4/WVISrwAzmEd5m8DvTe3L+oF0MeF8uK2j9fRlXW4Rv3Q2MUOHj8
7Ifg3DSXIlW5RTtPA5HfTeJGpT3vP8hJ/HiGvCxhuiD5diKLZEvpl0U2xMwfVH6+qVpTPJyHjAbS
+u3u8FJzskTxDQqW86CAwWJkgIjvZU6o53nQDODEeB0RdjtKFyAkl7bq1jJyOTtbcvAdlf2qfKZd
lnJASgXKHsjKKEcSOUhgWbPbqRABRbvoKPqpfjbLmMYLtzZf1QA5T8Li8QdWdydiWqPqBA7beFPi
iuImIqO9Kox/YXyXKtcYsAwKX66smJM87DiUG00KEqdje4/MoVNtrB+PeajEOA5T0UcM5SVsZXfN
V1q3IXPvpSDw0pNfpJiT1XcjK1gk+NdJV1lcspz+MsenazrpalJ6wjLbt2oOr0aVEOQHF1GmlomA
o6VqQ50BbPlOX9cPr5nWm27YpzCI9nCW4GJChPQi+je/9X8E3Cqwejwa2YIbGQKQlEeo/Wunc+Lj
109+pNVefWz1cUZYSFIpv7P9WRkOx1EcuKsGkppSXMC9ueXi0bAHFNlR4+PI7TCsFHrcRRrXBlzN
VI0Si4/ooLmMDP6lW2hFo/FpKSHV0ypLShE9XGYJYwUQ/+nJfg0ImG5ERvMQcWz/o865X0nu/d4m
UGGfRkOo4LmG0Csbljp1XeRF3+BwKYQzZWwHR8zVV+IT7zqIIV2a5+NX1iT7LGEZNIFE7qbaABBI
YsWgMeLs39NTKYzbM/WHsGONXj6s3vOjjS2xjlBTouPxeLYlU3oFl7DIEuYeUR1IXAnNGtO1BMs+
rfJorzuP45oUXMSU9RZwfMwnpH2InUVD/yRtkEYKrrbLNDXUJMb2q+y6ZaqDUA263hLIKKgKVJbH
6mxbQvfeiTkoWnXpjDlL2tujI6jD+weEmnXzdsMqL+zFs5mEAMID9q7x9O/U5hpBfw+57aPT4v02
xP/H0we+WSlyhVI5N1RMP5vbsmpjAkbtyUvkFtMTBssqM3xy0LMBuoQU1NfVGsp9KIZd6vNxtrCF
tUoQfR34rV3PI++GR691lPO7QqCGJy1lVXrSpWUSuknAAnsKgxssK/s1vNklR7fWo7YmrINbq519
BHVDVSB0SDjmb9vXOnYVIrc7eCS/uDovszaABi9NKUQXh5bfqv9HsF7AHXyhv2N9CtvhtPGQ7bbJ
FIYWasOv8Zjl8PungrkvlRjm65hA4pe105rpIVbA2R+qDoFR0LhbAv8BNziW4UrP2Ym9LUs7l/Dc
xKWbCYzbQUNF+Y4FvLkGvifh8UtiiDYjsFkuGFa3v+ufNe5P4TW/+Bn9whl3B9jJq+z+ZHvlvc6w
bU+Q2c1fiIg59YJBPg/C4zhQxkCqgjDBnv3oqnx0d2Y5rll+8VCZjS9Ve20nJtGC2plNnve5GpK6
wMLmai8hxv96RTllARCKY0GFj/h/+GDqDbw26HX3zq/hJ9PGa2/jBEituWpP1ewm6f9sfZXyLXcb
lUTa7mccIItqacpDLicgdc/Y7EQOBNfLsFieri2zxmsDF3D3lOswVGkr541QitJsuIIoZOz7l3Em
/iABA7hTreGVl9WY5kFQ1hNesWC2TfGOPrybRg22HMmiAWhFV2PwV6VfzbfGsuL0/f990/JOeLJO
ahW4WGN5wxc0ExP8Mb+RBAWPAEB02QAJfDFjpu5yws4cCuSKVx4e1GWYgsx0bvnXE6nA73WK5fyN
mQ0KCNRONVT2KD4t1GCcDVGsVe080NeEbEhZVQZze4/EQUhEjbh/IciOOTK0ecU2d4r/OHIjiiT8
0/YRyky5xKRe1n273bxhQhBb3wWCFFlVPTC0cBB+zfv5xdhrxb61FxftZi3TQ0Ei/dyezug6O3l+
owZoyAngpRE+TykoTzxL19qxlrlJEsabSf1FEH8ID8PP4NO3Ve06BzXDyS1Y8qpkg8XBZAWnS3zp
sLYaOA6LX0Dm53bZtYPWnH+2D5W1xxdgYs2nlD6Mqf9h3alVLbQef7lBxQJFz7YaV0hL7+LNuo/f
P2PkTCSYJBJJffL/V3IlWC2xahTiL11ZVNBakf63btMXjAoiltwn4T0mD1VeVm1Y5ZFR2ioKqCIP
ktC0MwvLq+N5m8zvI3yLYHNEujPuoopsdB62AySJd0MixncdwXwNfoXt9BByvxdCHx2zLWuvfqKo
o3oPYT/SCBTRtfKR0z+XloW2UbsX6RQB1cJhjFBF5dwNGNS6nf9QTSvReNCnivK+J63/PXoH9ZqN
Y6mrLVGIASniPmMlsmGsxbqPedwTWknHGP4JpvaYX9A1ZVfmpymoT0oNJz1VSGMY0XucE3Z97hTC
yMUQs3PTGyuPk2VdQB6RjNo3A9IPQVXMT6gPT5ue2uY/wWjQbBMdhpudIPLLS+y0devqE43HNKT7
Rda+eS8NS9yeev+SkLr2ANu9ovWwvB66gyyATZIQ/U83SYGcypqqhrHB4rPdXzCXXoKSXMk+6EYU
Apk0LjuR0yFaitCe7LqTnI5TpFhfq+y4Sv+cVcFqZMNiQWq52TUEPtheKWe+sisR3LQ+Y6kvusWa
OJFLGa5XR5QYjyXQbVNvv4HuYltEb1ozAl8azC45cAu0qecbhh/Mz8W2T1mKgn0dBWEUn9OQqJFY
fO4+p83E9P0FzP7u2g9spSxMiADwbHlgkpv5KJ0fk0TGdlLIHOcxEiK5dkDn5UB8mjhHE1CkUtWW
bKx7PW2cF2xbJKN2KL0EmKW4eG1Ei+xRNKUqr3tX/sN/ytCbxcvZ9tXvmZbaNxFs/mwlmY+WCOUG
DeAgmcZobH6uvbn9xrU9z4gNbPnm1a0e91vd2ZM0n7pDoSG8U1M9AFuVBuMSofOEotK6Ng+sPXN4
Gcgu29NFI2+WaYmHzBIpb3gEJHIyQR+zg3K6xI5bNaNtGnDrDCuFZLfxkWvp/JNx4J526r4LIMe0
y3seNTX4WGQgTu7wEdO7GR9CIf9Fn9wpzgEXbd4kl2MwfOjlzHatxDYIf3z/c/uDNEKDSNLdr1GR
AK5V5WWsvrDeL4r0uBcYOuHOVftmDt1zppuLTJE81ufXVyFOd5TWkxnU1boFADUTxO3bEf7TN/X+
Nc4f8h2bF1GG4t5EYzmHy07F1wBEb1rMWa5Vlg1f9KaWhUIuR1k52sYoa6FmJCRRgGUKtURhK23G
2JVmdPnaJB1vK06Mf6U+di1IK1nyb7A5MTG2QEIRSKcZ2I7QbuqbUrXxJCG0MqFFzdofa4znrIj6
X3UwxtbDApKcNnvNuAOims1UjRzqOkDkRvLwZr5OdF1ttBX743oGgyVBKHO787Gjn3+dLKp7k4oN
aKeCxoKmWEuxJi0fho0n+ZQlIO0xTlOb5DG9qlGMYmwzP3X7N62oTDR/gCM2R8IqbzK6K9wyaK70
7Yt201UqYrS02fZN0ySgs6MtffnEcW7ziLoDSw7F/n9s54ZE6V1sRzXI5Zw7XkHWgNc7Izde/r4X
WCPHg2NtZRUSmCPAA2SM/82kRSR7uikwk5qZMDqIKuqQs79MDqiTuSfdQDXxHEeqieiU21tOL5h8
FNiIjI8LWy3WmA3SKTT28mGWHCUV1IVkSHmzjvIH7JoTEvO7Tq3DaO1OUBIubMBQIiOJwb7J1BYr
ekPR/y0siWgJpKGrseBqRrL5cgSXDoPvP94l+7gwBhslbe7/Dm+BQm2ZY6UF/e+wGwoWVPatdex1
Bf7MgkcSN4KEhuNaVHQYlP2Q1nJO2KxwiwmNUR70HvGsIR18C6fDf3af1AaVHBdWcqiTkzMPWMmz
85hJo4a72zh2wHR7uu5i70BqMsMWlZpT9cLMA5McKTTXd/5mGjRM59knGTEQEwiu4zuA9IXGHQUP
13XnBNCbp9e0GQE7N7XqJGKs5ln7dHId8Ifv7G4uYSwzIFyd9ehF12lNq1+vQ2OmcKes1C0K5Lku
eB8AWmzKqfTlae5MmTjKFs/jpl4hvBW80QVzUq3pmoTpML4jg0FLNkFU+9E23kLR9jvvJiCqdKxz
LB63NaQdh6/6em/v57iBXTdKfZvpY9n9k1MjIj83Faw4SN3SuMeg4+zw6YypSwQsSgpQPXR3X3gk
avR3//IdLt8LhCkdfLXCqsKmm0bEyQwPTyLXS7R4Jq8j9HJgJEccl8+YxzNr+2EeI+JPuL4v6/7e
4LqzgMG09D0goMMqTHyNCzzimPQE+5dI5VHQJ597a1CZB8HfPUluU07j3PlcyMs0PY1d0YeB/gZH
pyOwDae359JUoEXrIm/H14ymRUInHZZscGylvCf88kg1Hmu/TD87rc+1pKsVbJ5X9IhRrqxjeb7U
CS+0cmdJKZqukg2M2GxUF4+mpaFy8m9AFpn7HHl0LNYij0flPhGgaM3Spq8Kd4+cJUZaLinckbYa
2VttjOcRSWxGYY0+4mLTK165bI8eWVyHsJInIDnzrWNgT5Ypd9c91xeLlk4zHk02AmQQ+SJeqoH1
l4+HPVTbNHMFF7RQPHKM/V80/1YPJgfkqx2munoHBtvVuZYx8b3fGMe3CeRa7gVbtjmE1Eo17yKG
7RIPQes5/urPHW7EmYs6xTB5lzfUAWt8lfvuMlXOnznn/tIn70JnP+XvIYfd7y/SM6XpVywky4Fn
avvjCnzbyOL7+qjIkrxQKSOCe/v056Lf0AjhxcVdQaSKOjPQeYRoFWT475ICEBSbKCq8X7vfORaQ
Kra1ILkAY4XMJU1RhLiYha9oV9SsvNdZ9sbfnsARsardv205AIvQjz63zARt1BAr0TlHkjHVDcg8
C5gWOareIjdKq3jNKBCvI1hZKhbovhI8zw2KJTevfXkRpyfbsk8Gj63slo0R11NdeCegMAX7pGHw
E+oLzDGzyZgr4t+FtXygTkNR34/XY2pfYLTMDRYNdBsSJeDAHFY8lqY83MkO2pEg8g+15KjMqwSk
HZQrZpN3khTcJmNAk0Go2D+8LeDtJFblaPzb6vvH58kpvh/19ST4NOk6ThYgmey/u96mu3/09i4H
AW1gYNH7H0WplqTiG3KhUU8+teaTpvLmeIY+ZhVvaCmgmop7iTPMXyVqQLeV6gypbeu/wLSBaG8d
0mLnxquG+JTnkgVHXdc4xWuaA22x6tyzIYrS5ZfM9NTEopFYPXjaKzXRCHXxqE6d6+KYxze7bU17
jdPsSuI7P46vU6L4a+vEd6773gFpNn4yXYoe3Uju4R8AhE/Xv/xHg7xtnnJnJ7Er/KOzwxl86EJ4
PvcnTu7+DNki0YEs9uocAgJ0YehHHmm1hsPEyKJtt8vKKRFl2mPxSz4Nf34miRIq7V5xGqAtcvuZ
zGkxTDMCFhrQ8BXL+tTXkZ1qCO/TuQj5oD3NzQwUtjJj/3uXQk5hOmPd5QhOcAVIF/FD/dqajWuF
lAdlWMs8YqPoVM8J6QORsTBBAou8hcB8QieyxEkxJYGTTwjmyekIfdYIsoWEyfgCFePABcJCH6X/
1tfRx00xYgIyQdUG3UF2TH7y7ZXIZMBHCyDN5x5oUZ4nf7aEqq4pgVotx4G18UVx0EPsGMShPD87
tCAQC0/jV8qq8xhgl2yogdZB+/IWEShu2LBkxDXvYgJKYDe0J5EfoHpC0pO0nJBAcwqnhZ1XW69t
wNzcLmtZ5Otq8obmpcGB81QZzTpBlRfZMfjiz+Pzt2h6rJTfCJgGFSoT07Vnsq5dTT7kE6nbwAOB
yc6+SGzZ4nrL5kfUaHS/cM3wytljHogeC0jZwZZzJZFVog1LSy9mOAlDbrYkqCX8QNAek7IEa8xS
pxcHnLQfd/wcdUlw66UrpFFbjsqyhicM6NrZF6/VrpCZNUjpa0s9/TB/EImx3b4qgluGf4zAah9F
laAR7v/F24fBdAUjmFPb/A5/Nx7yMI/LfhqXQy/T9nW09GglzbKg5t9ZCjAvQpRMXcvWPNZK/sQj
fie+DXnOR/cuW80QfRyE4PrU4LBuvt55Xmwek4lw90uf/ufBL4aNtUGVKHz5NKpEfoxK7wEZl6Yk
XIy3ajAGAitRIpE8oUAVTIdO+Q0uskJvak/os+LWtWZSrEnReICPhZV03iO+TTbUdEvJbnXMrbUE
lXifIVcw0tXVWYZPExD9pfaz0vplU3PNugGoHkAkhQ9SnWFDpNpq6WpVxL9Cox0sbbOqHr297+ZP
fZDxbEkFzqOc6978JIxx9d+eruSCb69i+Pw5Q9o3di/VbkuNigq08kSUQwrJNyRBgfRWIYGLjfWZ
/2M0dGL1yY7pCnuDFCd3xEzXPfbLCRx/dRJY1Uu3+mPN8r8fgY+8d6e9PRl/YuOBS1p+l4fPu65T
F5hCYPdWEj+UFZEEtU+cdiSRruktY4mE7gMEJls4aNFMCyWsQZ0n38JH9IfkUTqQd8EuvRF2qa9y
bChKL02D206fwmOAbMlVnoQnGOA4R3RXrVzwEZy2UvhkHNxuyIY1VkhkO4xGgaHUPQVIatNMv3VG
kYo3dOdWRfo8Qsz+83HCzSyJTMGS/YY4cQpimmD8QdcgZaPiz7+ITR4ms92faHm8CaaUZr9JF8u1
rTEz6xuca3LSizQKOXVwUHyfZkWRaBTVXDiUmVIevy3K6iUS1w5QUX5CgcPeKu71MlmB//2Th5eO
6Y3a6AQ9Rgjx1MnuE9WdVWNJwnn3gDXa+5YvscjLTHirrCPlUk+YAxHQKxvQfrmym9bVzc2DXhZB
bxiurRUnq7/j/YF0iSrJfCnjjUyfKkmw9bmL3LSYu9JClaYN92Wdi1CftsHoAECqIWSLnunUSwmr
CI8rRIWwl0+k+BfHA5mfU0Q9BwfdQPgr4BR+osHVMCjXz1Rg9LDaOUpIkZUTsBLvfXxTnW4vGrh+
5FUenhLZF+Cr9FonxH9/Ob6+8GllLeEDt1JCnSAUpHDqLWwiQsYucw0EOIzdu/wO41rnJX8CCE59
/CmZr8LD6u1N1XQjyuP6ASMqfby8xkOYGjKP4op/AHteabIMmRwN7GULyCThZcFnp7INRx6BAbZK
3e1tbZ5j5GsO9LdkBKswtdUbkAP2JHQwKHD5AUwTyxN5N3OH45zcCeAV2+a/12CAnhzWeXBtow2g
avsX0sUwAG+97QU9eaBkjs7A8sSWxSef7v2J7OVTPnxUWrp9tsUM9LELpJ39URTtlQo3+hml4O6Y
Ce54VTiqPwJA3Xn4swIdBqm8rtkQrn9bvbN4RXoBtV+Wbpbg8Z6L7FJcu0P60MFOJE99gy4xcZGn
3CwWubf9mf1fyY6X4jycoVJnkkDtNQNOrD135y/TISPRYTT3tZ4NaN5vDvg7b7aiS+6AtZcuhUaU
7jss5qcAaI9lOx0pHbfmcx0McZVkWUiRrrAgAs4zSO2Xb5aTuhN+SfNi+fz6qdNlcVnptYxYLxqe
viI8AyIANB2UY4//IOc11fW0dm/B337VRUq/fcahP+ctza8grdIVz8gejSHAk1KeTUg2AwKJLr3V
wmGFG3GLEuxZePb8ewwEjMv5DpXemYiOJQPlDWD8emVE0W0nfvcZ3klDo5f+dmcYgoo6VhODrg+Y
izmhXnSzRo0SIeq1a4QbVuedr+Kmq213DUJQ9J6lI9dNwC/MmYJ+xCtZ5oGf8hz6lRS0Pt1MpXxf
dvSVSSksKSlqZmiVXxI3UWFr09zJS/mdZ/lrARmZs+6JOmWBZvG5koswWd+sPs6N9BqqpSdf8f8F
1s1DPMXvEDh8B+WlDvIkuMkqgTyvuC2j+m9vqLW0d2e75Ln7iUIkWKRMsI5dwsJkVcAWn7A3kfP5
41n1xm9/idNzZ0wWfvNE/3YlRfp98G0hi5ugzKXpI+vC/1A9iqjbqntLmmuOX0vBAsglfGbOiq2U
mWYaxOkMYOFP+v8aTjetXbPn2sku8bT/Tch/W3MPLqfwscLr0BcNlJiGDp6+zf/y19I3LpVEhyNt
qCSryNeBko+o3BUs+HBVgkEFTwr4zHiiGqt4PHTHZ1AmZZ15a4pdkQhqbQFtjLAtT5b3q/igaekR
y3H4eKMNQCLfTy+GZX0BJTVl+C2jEPAxVaHAr4Sc8kzFCsf5Wx1BTmFnEH9vqUGLk5SM8TQ9gC0+
/y2ByVcJQZ1u6uHokcsgMbeQ5UolkZF4M4fSwN6zr2PJp5ahs90UDVzCiTBuOfsqULr3WAzL0bKr
l626Q3iiPWbjrXXbSjRY4znuPQUrWmJIwmwk7Qtf/+H/HJgV+njdD43L24RhlxEos3nwHILFjSg3
zHGZF8uDBzKx+YlBPF/5IjwKKBcdq9PNofZAJoisfE+3LfWcp5fM0v1kc/aNvzmK+i0yAK04XvTg
oicKKt8mQOekXN2OtDwZ/F4lrtxdu7xUhcOzM30e2M8klPFQGBKB3iAuTVkXosuefUOT/AoXbaq3
OJXU0EFBFAOuuR+dHBUhvSGVrGdtKclA9koc7QdT8trsSH2oDe9Fez+aWT1Um3KQ9u3CtH5lCP+3
0zs4eS/owFX7OmbVR7GqcpmbKQjdMiV8A3Siftq+684JNRrhCXGLe2V9ZouADg3bMIxyEA4SmzbC
FosDXfDnJ0SMsXxUnEHmWijGPffTSdMoim8PBV4KLdWJo9CBuXcqdKy8ChEpxfTdoGvTkcth2gtY
7KwpIAhB27vGmOQWau7w0CwH7WyLtydYtYtVb8RGPoJm0QErgRKrVLKJJvphWCgzbTeILyFUFUoL
oG1zBAxYNhvGmWqWnkYJ/vMQD/Kn2h4iuDd6Wjc2WODmHFSuL2JnE2+cQdQ7y6ld4UerqLcfzxZK
MZMyFaMfZM4NYd88pzMjLghdMjpOh8Llq/Zh7SR3o11nXnJ6pw4S/FfTmzOLyiMnxkkm/r39A6wJ
d7nMWwlSZNv7or+HSSM75zydG6OR2O5SmAUn6/ENi6QegqYycmikr29poY4l1o33TUPVI6kbKg3G
Y3jDD7/RTVn6WO1z/kUl1vdUs/UGNN5ddC0kJMC0n6EFfuCHKhUxk2Dxe7zkIa0G3f/S3PMXVayl
jjqVSAJz87Fqpf4j29qVpsy6IoBSQl4yL2Vy8rHFUEG9yzjFz7VpsO8Uu2YzU/MYGewfJ/UkoZVb
KpW2PHrO3BaderOetrHABXZ4RZCVopBQXNdpux+fAh7bhcDoD8CAB/qWM20Qr/lDqhcxdWOtCADd
XVYFgL86fGdv+Y3enR6h4q5P8kfVWvrrUVnBralKGUbOMyg5DzQ+Gh6wnCHDIEsauItqITomBgP5
gdi64FQb3O3Iq5D1diHI7uoRvMPVwBIC8YeYHmFKCpqLb9migkdSmYzl4CWwONnluRfWdLgXRp/e
Znor8iPZQOANW7cABJuzwOjvvkbDbPnMAv9KVbaJvmu929KOClvBK9V8pCISUIEZe8zklbF2OCi7
qeNano3lLKiqoxV5G44aTGZCygudRe/DrFUH+biu8lLBj11rylt7rWYyMToefB8satcuXTGD2bF7
Le8F75SwYZauaxSA7PSJ/ss80N1A6oVY4Ts4PdpvsXTWt8lJ0Mfg77NZKotRQxO+cudX8HMM1/rF
qpKUeWlB0fx3xH4GLhAN9bK3adCjoi2ycGgMtCo3O32QQsLdqPtq9UvvQ0o6PffULUKeasy38qp1
Ji7j/d0oAIz1SPqrDKu5/QP4GMOl7BXlS/ga0b2MBA6VaERNRyB7fr60pkoqLGtVDC6rUnflQjP6
kQUIeCK4o79KGwqE2zZwSinz1RlRZMj4FWiS5oVZ5Zl50OG6MFYgFspIuIXQmQSkhXwSjeWpju3m
aGWqARpj814j3rO9zSKQb95P0OImcEc4VY7F0RsM/QGSHgCn/Wx+JWhh1vDGSubpZwFN2JLiXw9r
QzuA0nMhy+hP3xkeBjKtqxXSD3/RMbkrxW3W8dVRoYrIhxwedDKxiMjD6BgtkkByNkQwrkTO7DZK
1bbNZAZQejcvoBHlbSlwluQsr6Wf0yrMe/sT2J8paSnlsMoMuH4G/TkYKGhLnry8RMAkohS5MYTH
7yvnyUwO8OqFd/5/w134VNrtRKR12y4+dQhd2EWy0wOs0K8a0/Mpa8Ni/ul/ex2vmH2ItgEdk3mX
eMcbTgQ4gaxK+WPWtPs4EOKlerW7FWOCEnv9OP7zTKG7GDH80Yy4lJ4k/F+Axw+oDYHvkqWxKEGX
/p5d1OsQ22kIBFIKwpMjaxBZJMg1p1oRcvLuwNo/JSijaeab8PqejSkiwA2JeqVLX3WgzkvU5n0B
fTdVsvuOL0BHVGhREDqOZ82KnJyfyDhtdC5Yggpt4+sA1KMyG1riAcrQP3zpclq3279PKnIH/KBR
eGJxJYPNPWIl5OrFgqV5540HCWE6oEhdYQVNZxXXQjH3MicmDTQyr0ruhp7T3Mb2dheJQnmGlU6F
1zZ4FHzy4VY8IGfdPId5R+Jli1MG4q5GBJIfJUiiE1aamh54PhtgPiTcp6OKaQuhoUyqjQSkWYsQ
0NuEkpY4TyqUUDdSRJK7AFbffr6CiUdM3SaJN6G41XdG9ay6IpnruC9iIL7R/Et+ZPrn8jdqqRKh
A3Mv8CgQyhfCe+v15PgkGfOWg1DG+0mr6qfDDquTOOSSfqLcdSWdoP9i3nFnDgFMNS3Rcf/adnyF
VR1BjeDQwYxBRY//D1jfy9q3He0TaO0VP2+4vvLLLqRzvhpVEvGQZbQiCZ9kwWO9dbMpWB7KBR0y
m3UGBofcith4646m4XMjjsvVzdchiTjMys+O/5U+5LGSj4m80i7tP9CpPzEvjj6wgoHHmpE+vXhr
+DC+4zB6yd47peP/oHKomIn8wVNMYjq7eCINCUUWj0u15eR+nMbDQWP/mb/dwrjHe+OBTAApV0F5
afnOKsQXN2AZsdQhmVXMM6FGWYCd6Fxjl5tJUVCRPIOMAiYZ9O2vzmNmXT1lwKP4b5ni7RbLeTC/
7+nX6he9fY1zDyN6rt4qRgRx/g8sJtCARiFkpA092/KSZUgDlnhVxegn3uHlpUDF36ijfhsE6400
XpgtlpyKo+eJ83PYCNOP3dgqzjWOz/suy2/CqdRQusDuKyaIM0c3Q2/kPQ5PNvNcyNLFhmrEOdXo
wj9ZD4ePi5X+5pHqFsajYa3l7X8Gu9S6YJenoWfkCyEJqxzbeHcK9Rh9RvHep8IazPwmcSnOV2hX
PYtezZzV38YR0E2ztIZW/8xUPTlDsYwsTSkxCm0gzcZTztjvJgadYwmUENvKWHmY/XQLBMASWwga
Q1GanA3cJVaXMFu8xk5WlavHsQH2Rz3lpsF1a2dObv0wxePanlq9TNDMs9MWUCuvWKLRoiA6K57B
areVePLj1pVi6fm1X2e2vVGLbgEKaLgmbKkwzU44KoU/6ix+y+4vNmgKCPI7EUhvTtaOelpFHwFr
O0iyySC4jWdk1TtAksmgyvIuIU6Z41ythlrxqdu8xSvxFhaRpo1nSOJlBjgdh9HyuUk0z0euaU5+
qoC/hnElI83bo0i9kyDlLDbVXfw6ij1Y7L4LV/miTcqxcACxTbbe940Xkfwmgctf3p/I2qtx6UTX
ExXM9+zIh3zhJISjji6iDtXyJnkaqrL8drT6a9bY9ooVSXD+5+hwrA3o0QEadP/BWdBiLeWm6icJ
/zLqnNqmXGilPPyX7xImuqalQqsjWSJGT0Q1iX2FN3Tt6pDTbHcdevY+t0rzicL4rnh2qXa6aBZl
Aa7g2gVbNS87LdJtUQMvSW6gTIAHL8DBK011QUsjrBLQHrama/Igl1ktx3Un9gHex8SiT1XqzVPw
Ik7oD1tw2AVb2wTtf+RItsOl9MCvh8Q6acoZX4F7LGfVq1BiV9CedyqgC4gNqNbuE+SUXueqEjrz
CFADFJRZIly9kqcjNXv8kAxF9LB6+IUdK9lZpxvG/uuiWGAcISuaWdSzJNPQLWCzY8BC/N0hKr6l
Tkslja1kdTdLqDpStttF441ZkjtoJI3QxjgLWLNWKJoiSxjMEPEqAAWrgvq7ZS4vYVFj378Rzbid
V5t+N4Jjhp5xHBpoTiRxvvL8x+apjSp613uym2iVoVd0FBRHeM9kngctxJ8Zl1iFnlt4K96Xtyt+
3q+UFps4lYiwoxag5BRWkmAophvJUGBIAhcHklzbSXH7gM3KtqSX/Ttc9sadfVUU4I9DXpmn09G4
ZQ/IGnRq9Y2XrrZpwgMsyEaUpSbH+0oJ2ZUqj/uv7pLC5chUuGkmT08NMBlWvBreyU52jFhwuU3F
NiIN+WD9xZRZy4ErUXvHUJxAgKXIBFOv95oeqVG9Jr9efp889/BXhlVgr07MjzbqLFBA8Inq/OOI
Iv3ZrxOTZaMBot7OtBvJRlcbZDioThJZnjGOFbhQZfZVATUvrgixOEE2U52oa+g38mB06RO5gpae
oO3mx29mTr9KYH85cEenXQd9AK2/OI/mXRsybu+9P4P5AteDXVCfId5F5A+fLKAZUvSPzH3KGuAa
VOjpTIGo3sMZLHpdxqyMUNn2kktOYB3n7vPrFAeRY4e/mmJmmTNaaqfFF8ST4Vh3ZAYf8s6gnhpr
DQlmc+KamrL/xRUw2ZUFCLFwdXiwljFiOzG406t7rMO4Fd8zZIsZTd0Y18/uOlP9iId6/WpbAEsR
UJJKPC5EYzgpSAh+vjHeHIh80NzLuKtd6iN20J+XZtfGQDGoPTeqzAqo4ZDKHJn300ZdRX/EuxoI
lfxqPnbAkWtrlOcxpqimqnGnh7CrixXZom/1x3u0eTAnBIETUrBqVcdfjLQh94flhnxDxyfjfkzL
Zm0boMMQYaO6czsy825k9iU8rGoTgdiwNvI/VpQ95b9DxwqA3YPe/NMaMvxwDk1hZNbM3uVFrP2N
UK46Eur3VnRkwfSKQCUjXm11rhfWWFBdOOdOLgAWf4QL8tuxkeoSi59frZc2F6PvNv0YcPpHInA/
Ys38ukNZFbGXjZbSEFCtP9g2pS2LYRLurZBnbP+eNhCUXvcPA3SDRid4d0mLcJ3RnbyTs71d1YPz
5G+IoWO2Y3ulD2QA9FZbVkW4Zb8iCvRA9969w4JvSpLb8udpHWEK4ah0hYkDcNQ9G9UR/m+ATQgI
fFctSWmUoXAVMyx3BPC7NS2Qe3MryLSTsLvdwKtCbtjm6dHFV+u7+DPgFZD/IELSOa6TEIvrrpbc
nNDQsELogwQdZ8dZx8m86UmM/mK5IaZvaruIdQCZUQlidX+g3ZVA9DoiKrMr1QSVLN750a7JhLK0
vQjus/KXSSUPBNiYLjSLddThYC/yv2bLU/T120wA23NuRA8HIgcbncEVI9ygZ+sBlt33AMSRF9x2
9LEnqTNttiJEc+4L6fcZSghL5pqLOJTddDiIIlki3JOJ183FxbGDud32Ab5M/iOXz+st++3CziR8
wlGx3jfsc+CAoYW5DAZ1GdfUGyMyndZqr+nUkL4MqGrDgES9ENEFCj6+QcL8+DedeJdSGCKkNtC8
sK+TamkSieTrCAWazkSfr71GA9434z8Fl0GzYcRDQJHLdP78DbSBddk4o2HUvUCCCFl4sJ9Dr615
Ts9oNMtzWMQKVPxa1wrESzGr8LatHrDA1PuLMIdy+pI3OtGwPBj0R+JsQDh7QXNCHN2Sn+ufC1V6
f8wzFe8cx4vY0+XrWQifjb+tcKacQMKFssUhQ1vaCZaZeUIivKBV3vaby1xsQ3hc4dRNeQMsJgWG
EZHpu3ySapUDAUL4MPko0e1NhZBKHvpMp1fF54rXgKHe3RsxaIFoI0xoblwHDsl3eyfdETBffKgC
CmWC/UkV7SGmndBODfXkAUnEKwlFs2NNoL55juXTpfq4+Nj6ukX62T7w11dJ4yy41ssIKw/N9ukc
eDfnifpzfopxeYGcqE+Sqv/eamaH8Yxy6QYpVRzTbj5x1m+owpBk+ExqwT9Arg48P2tFplDfALRp
6z4YR3d6W5o7yzotgX+eUu6hZZa0OlHHXomKEQAgpWG60QeInuXFW7FFsZxxjDGtknrUI6k6E5Zy
0H6/6eOtIMAG5QC+rXOYkLFbg+aQAKwSVvXTSdvFdBok7KdOIqoMCXmr1glgVuWPkdf60cfmZM1a
skhDNGzuaEkk0R+pGvc1KDXMfusUdHeXt7keFOpTcuZAfh7fX6bCa634AB+sf8432bHBpcEi898R
PBLmCWvvybAfjoXLG56h6G6wddYxaTzHx/5ccFmqevfdtaQ6C2H/Kb7Gqg7dJZz7uVAxykj6rEdB
FbOjGboRTsR4rvONs4zlpZYwjvXYCpWswUWCPFY5zx6wbr8ta5t5qGkkvhh9I9ClLmkYFBbl1Te6
2pEha/3GjO+0T7xQROhM7RtukXOlSpASsBNXKKHr/YcBqviyz8eV+9hCoLyF1nayTu0RBbb71/2f
l/L4kBw+S4WuRZTvdZ+aRMdUrxSjnnJllyWOrI6+tLd4641qfMVUn63GrBJGRt6H7MgbqOcRTWEj
EoVIH2IG8zsLWFSS6NG5R/7BFU32kmA2PWA2e03XMMhsBUT16g/xmI4jLUpM+1SzCLdOaaeDd5Ff
JZE5zEWwVbLNN3iVkJT7YyQ2DLBwMjV9clctxcE/xzspo5/PLyqGnpbK4Y5RS1kq+5JxdEjo0FdY
lKgpBHBBvME03HQStaNCFCwl4CS0aU+c42wDBLHXWei6R0xq0h2//NIogu9VhAyKKWxf6X8VnRwn
H9DcK0JpTeQJvPRrOnvNMgyI+/CX69Om5cvysVjOWcOch/jrm0P1S3hq8fLYSK7OMW91NcHqPmTT
D2XJMkgfEQl5Q7yeHBo95TyU22BuOjesfXU18f3JpNV5KxpHwFRTIj9QAZNv7IdDqr/X5TtszYTq
wc3Y+GCVJDrDRlk6sLDkGDJyKkuTMWyloM8YsKWTnT1+L9BgK4rN5EOIH6iGHm3vuWJed0SKDS4V
oq64kirxJ6Bi1v9+Xlp5DeyT8qViGvRWnvRc7we2/nffeRF4IBjjEW1n4zQFNKobNp0VbCJO+vo+
XEUS2TKljwLDHhIUKEWk3Vi5mONV/OH6qoVmbFinPXG20g3csR3Cbrv2EUIhf3Erf8tgyBqObs3f
tkJCvaidlZeZMYj04s/NuhKbP5YEbxglE/LVELBTAOlR2A749z+e4itj2TfKwrIZRMYYWzQMlhw4
08oyuOIIqTA/uLfijNetLSofhINAdlimqKOYzuhwA56Qt6L23A/aoldX865RwJAWd2ivx3B50lq9
NxitN/kgOqYWAODYFCsiW4nLW1VeQI7P5uUrL6yDMbdS+jJOVRxBtY0ql9G2fBS2vnDM1GMid4TA
68qpQvFr1Zn3e9X/TFnjd2/RJf3gMrZ6vF4V9ajy7iwiP2slHy4k5//bxU0rFDX2k5WQTKQ4fmXn
kOLy8FvLq+QoyTdVxk5jPqfvcVv79p3aw8ApVi0E7Hh89deA33+1tLUi6i55d03f1h2vDjyH3oIc
M5knQqV+LIbKJJLqxi4dzQsYJbMp1tagYmBf9UfVVakv8ie6RxL3HdYTK2pHi61dxmbH1FU8Px85
RXMLcouOUn627nH+DagwbrrY660HYJMX2PcueII7eAx2mWsRIVMi+CWjeBcpCztI2h8mJtpdXqtg
OCPvTtFtV1ED0h94/okArF/+ZxmcNdMSnaRRSM9uQqgZsSR2MbRNJjL6EqJvDM0XYEWg1tOAhqHM
K9JewwHx/ekkH1KImuD9OVFnJfpqCrLtF0A0DDBM1FcyqbIeyPR8W9s+QRWQRZjXXWg64bONVYdr
OxHp2lHGA0Dp8cWI+Jr6a06XZ/kxjgCNGg/tGFnxLz6WRQjZpQoeW3l3DbKXkj5nsLfSYy9kGRS2
RltwYV0/XpdyAh8gxU7PbovwDMcj58S7MDX9vhNFVEO1cpO4FsykFhGxvqkD3qp8aG5hiX+o5UXP
E37hPSVce4XJtSKTUvfcwGSRswSrSfs4o5vvb2VzNI8fQGC+sjdXdrGad3xJnPGLjD9nu2vWnxIl
FGRB1dEcFCkyxeOEzk2fMJ41yIzdlX93q5AqKBsFmB1RnuhnNuZGWMt/jjKrWcMza7iptHfeJmuy
P8YQJppGRI1hUxZUaPjrhVdb4gD+VtbzFZlrIy5sHrrEl4P3xA18OwosW3FdaDJawb6c6NGpRcsC
rPJOPLv9JXUaRo2zqeNEIUxtO0Sc3/OMd5Hq1ypHcTnZ/WYzn7RrQZ2abTDRVaKkiBAck29dJy16
9K4PlKXQnPkqAssvr1cJmD3P4wYwBSscoTKFEm38hz49GwoIwb0ptsbUQgoG4FIICmY9cqSaXsnC
9O3amvDZwrM2c6gw7WYV5i0OaR42rRZ75C50FTzVDsmiz3tOiaLo8hMq0HMNVFchylcP0c3HAHpF
aZOKVGxDI+U5ADgWh/7+PLmYIMRxvZ9Z4eNxVH/OXPNMLqbMW5BUp7eo3rQyUsP7bA1+OkXgmJgk
KskUd27dH56/P3lsiWQSW65bm7CkxVC98xv8cUbxi23pqaiGLjbYHmcBqqsuReKL5dPvbBDy2wLz
qPB2VVg/XwTa6yWekW6WdtQ4p18dptOmqlfxQVYSdy//Ij0XwjqlcugGK+g3hO1QOVeCB2Rv7c28
XmaaHPDSaDJsZLUrJfh6gZND9CGernySt3mo4wEpYRGczynZSqkYMceNRjPGiJK3PYP6zakF9X+n
bguwaZqIlwvT4v82Ib/DMEBW7W9IyedeN2VF4qam3XD3RMf9zcWKbBxtPr9nrktDR2zOPwaAScCV
KpmLN9SzX1yFKJsP2R7M5WnF424BshehdBk248nyu/eZsWhCZPhW24Edq+OWzZLcI3iV0OsSEq8V
h0kvwGqYklzsXJ7DRmWrWft8wS9TFrJKRiP6PimR458Hlb1P7t/El6dQAhMWsRkLGa5xlYUhmPLZ
mOeMSM1VvM3EOUM2c3jqfwU0BsrxEXlSt28w4EfTxqiPh4GaLvhAMcawW07JXZWm+WEWU0NEO0u+
ZEayQcQI6UQZSvVywfzbB8LX3ljRjfxz4cp3JdGfkWd+NiYNmCRkAGoraHMe63FysrhqXSY8+avT
SRsQQm6e8HCW86070uD+kKulyuJD0wW8Pwodw09UMrAxJKKHODRx/reBAo3i0tSFSglC1tDcQhzv
I/OFcKhDCCTcleAP+QHsczS6e8EjzbRtFLVLUfDFZoDny/nUZflfPjmKmrjMwEMoSUfZfin0rGxB
xPDyTgtPZM2WetV2N5j/u46GG0GJgECeKm+xn5Bybieqjlnz0/fiTCdBDDsf4/aVBJ6xGSb/NqUu
L3aEIIwDJU9lGXkSe5TZnUEKCS5vpXPCGtM9MDWvJzFWcM+MlirGrbWjdJPeZSiA1em62GvTx5Yd
DE9ZT/rZrsKn5GYFEX56UQ284D+i6RibGj0XW0ly62g6LnxS8JZ8eiNdARuWOMMKSZ6OFV7M8cQL
c5L0CD43xdQKRlQQkXj0jcaUr2V5HBGQfcBqRNCWNCxZVFwM+xtD1GErir+xjLJFXTXaRFxA5zbd
PVH+LBl3cbe6oRujjqfszEFgqMdWSF/li0vP8R8JXId1X7fv6Ius1HyfIk0njY/7XEVbRm2KAfJt
TWtypS41qSZpeq1vOTE3cqqorXPxLXmkMuS7H3aT1ll6K0UfJ2n4AWvXYumhhtyDCNMR9ZjU7ck9
xA5f3OP9IzWiW27eVC4/6O2qt39T6bT4n2opmb7Qd0RYUmUV89/XiA+IqHkOmhyAJxa+oKJV++Ct
LnrPeZQ2Ber8hXcVyFPsnYS6FRVy73Zy2+uxcFZBOFhvqKANaf18ssvDSgiiHrGmBa2Z8hRXR1rz
Fsw5vE/5Bz3h2Pdglw61pknJ+zISmZX34gqlYnEdkX4DCtNvTvXgPL/ssfijtlXtGudgUUbbsAPI
UUW9XenP0nniViWeJDLdN8pJeFrFb8Kb8H6UU5+mCBNgoaUtwNLDLt3KSA8ayd/isylLmok9Ol1k
AmB57X1G5+2YZV/JSZmwjjpYWXlo8Epx3ER66rJ2VSFf6oFFRqpTbpLeA+zs4pfPt48eTcNSxYK2
JFoAK81G9GImQC92QRRgCG0TJUfWGg7TYw27lF4kwxESgLmf+2Mujp6E0ZPIkzy1PpQJeNnWTNNg
8p1DM2aCDSCkJjUCLyYa24odE5TimaIrSmRGDKzfZj+yCJa1GMTg5/SK/IdPRdwDlccMq3FKXEKT
InNJfH7x0qAPWTLTWtGIjAPkU6kOeQzPUwQbubq02ZykubIDJs1uSOTZbNf/XeHj/Nqo4NK7PNTs
EFY0gMah4z/Qm3LBI3DUU2HkVEBST3BgnvVAMWOpEBLVW74dLQr27SBGrpsvNKPR1/iBpvqTk/Cj
XRTG2GJdWFwFtY8jQQlL5SjBMeJNsHWHvpm3wiBIxHamwF6Eue99sBOVBcc4nvIXfmPO79axxax7
Z2Jy6+GcHGWQXyCpcTaohxiow4gimItK89ojYaAg+FqaUeGX8zbm8ojYVqEBJJP2rRfz6pg+2YVd
SHsdKGj8NfWFo+KL04nKFqCxrl7ZxmB1M351qZdukIi9v4I0jmlzLMQB8B3CHRunfONeIeeyheWh
h+kHsQYgUqOZEU+WOYGRrj+uYoS99k9XmcesSg2wTgY27OXX4EwtzojK6Irqft0Q0wfjxceegbGT
cFpGCAxb2KtoIIcXJNs8wfniciiPi1CrJCXjy3KVObaJKZ8SEOkr2AH4w0cVELomgqeCeHEiy7Lq
Rt1D6D7gy+s7yR4GtSrI13iYNKhZDXrCvMW4rEcBOEjPhjSNlsai/WbIAsoY2X2ZRhCoU2Nni6JW
5PenawLhajAPn+VVVwthNWwDfHVBjYFU3P6QIjUNeL6AWSMEI08H+5lZKVUVpJps+po7vpLUZBUh
x8E/Y6G0tnTbog50Cxpj2EdiCdZlvvnrytjygo+29kA9bG4pRTnJGUIhc+Lcf79m+bcHSvECl6Xv
bHo3MhfvCYaijL1xSjSkg2Og/ngbx9ctlL3AZsSOSNtTrKCNZjRaKctP2cY/5cfXnih0ZsFYvy7Z
zdQDddFgn/fJb9IBXDJklB7Qs4O7eWzC5feBykCmqox6x4mYAJ5YFi1U4+hKzokbPIQrgZLDgArw
/wA9lgvOVb3aE6eTqLRhULOeWRbm39vgjutKQh+lA2pjo6swtgw9Rby2UqYXCKaP9qJMr3KdNTQ6
Tqpyj8M8ibvstsVzVozfmtajbYJUmr+CBqWqe8ADX4NVvJT7KOVzyTWApfqllV3FcALpqOmCRqP0
35ICfj3f01h4Pa+mwl+xyhM2WoN6q+2VLFlF4R4z+pgT19Tgjx2OWjJownwCIx0eCKeJa2ki9jJp
0FJLjwfqj2zhFnTofIjxWqGfbgVwHvMFSWJ3Am/7mahViI3Bs06fA3xAS6Ogh67/WbmvD/qXfWoN
f0VCnPVJXgTDefmYePouttVO+k+77LuHJCH63109byKuPih/OU7oF13CAkYFUONhgNY+KEiWf7xw
QCCQQHzLbhKXUpcXz2P8WRVwf+mzHSZzrLQ7ANlo2Wm2fWzG3fz6DA7zFglCo9g7Gou4oNP6SQ6R
6v4pAO6k+zq9y8gDhJPI37jOLtJoDLrgoR9S+Z1K1KDsATUT6fUOrV9FQXUdZI5bzKTPicwJ89WX
dGtC+uR0QAu+IzTljj+bbThNr+gJEDMuR49VLZxw556Krfz5DBctcc6Lhmox98Vn2jVrqecHheyv
TpmYDQeA0lQHPydY2x7sUTTiGNHc2z8O9jzCTXbkuGwlHu7Q7Sf2gPoZI5Mss2u+JtSHLqBM8Pqk
qW39aK14zFQzNQ7tST4SnVPjNJ7y7GtWdiRrhRnhCG/EkEbfKvaN071E8VLnY7BMILagZJuLdPrW
DPCVuZdk4IqhYkkcNImAcY2W8cZeMX7nlk3tA1dWF1lX1UziGMXFmI5Urt48PEL4/OFiQi5BVhFH
k0uoEBT9Y1jSqo5uN2FyNr+OIK17F7XhLeEXC9tyfqv0QZug/O1VG2yaGwdh2TDCFlSg0rT6kisV
A/jGvAbStuhWMVeWucglZ2qnOgVHnPCV0tVhOZfXzELXRUyzJHXG/H8F6D2KoeBSWzdOmEnH/pUS
jDEX52/lLBYVbV8NVZDYMugH7q4o63F9l1KftQ0WmInPHB64Wxemn3RYrAJDVzOqKzclWt9Vw8o7
p9N251CmI9XLQXJ3tN9EAvX4VuTwnNtl3cnK0vl//f/7QZHy8VGoy32l3JyIsky2au8M0if2LqFS
5E38ZBY4YGkUcmZ+s0lSu9Lu3ZilLzsuBpXrVxCQ4j+mPeWkgp2x9a46796BZXe6UR6/k8e1W/G0
DNhy0NLBUUcQZjM4uXZzuAP7lo1+v+E4A9gZvz6oY3OB3/nSiELYVXMARQVrDrb9NOZi0WnNuN2Q
5q6sob4tIleG4aqIiy6EW1rOKSvjsU393ZlX74t2IYUDi9T47e6ScDJu1HJhrTAfRbkdTaHBZjJI
6q3IQ1PZCJ69V3bpFuIe1XgYKkG8jiN9sEqxlwUujVpyNW/zt2mIxcacr+fox3JyW/SBAKtDpnU4
Rhxh1os20Y05V+4IfBEuABDFJgM7apE75ss7m8/xMYNhniDV6wPpBpXmNtdDrupEdKP5h1Mvzl5B
KMRwOrFK0aU03sJ+nBafkuR3gPXGGFIRFqfrPDJ1Y3RTVcA2WBR0WdCbg0naQ6UXLXQp2lcX+T5/
ekSzj70bnbWIe0stBt5Z5lGZfWKcqI4KfWE96X6N8BJeIiCnIXBpOG5vSplHsW9U/N6P5gdJLBlA
i69FFzi01W57PJSFZov3/XVKRCvdaIdwxFjNmOEq+fKeHVWEGDACtjpdzObsdbIt+Gpe7FaNXzz2
msK2MTBIigKk7yxfs/YdfAtEhPU3pHzxKWsdk88ipqIaziUSdbBHeb5V6JjmtXmzPyTtnd3INeiE
mvz6gocU0z7pA9fIv0F15u5EWWn3JJXcc7UNt6I24Ia49r8eYQxnrk53AYOAqqopJghJcihJopci
8OIk+Yvrrsw7uj1WdMTaqwCERGacPl/8nSSU3Tc8xuSVBIVEfKhYGeYU0ROQ647whiqeMOBHLJMT
cx7Ooxka/TePp0eCse+g0BqqGyFX0pGESgKhTFuqTT7cVDMGAbrJ7zJ+rN0Alk4qVi81b1h3cx9D
EcGMWdOQoQZYOOf/2u/vXlBhKCLtc4/90fP072IBW6c3ROcaWN2W93kqAM/6w/GbWGdJuUZLkyMI
RruYfTG+qExy5zgafg3VSbaWbMPozG8UPoOoy9obB/A/+MmiGwDzD0k1kS82W6pnTolB0cUCb6ZH
wcJ74Q3tK89Cm42FFk93PNuTqawpvkys83izKq9H02YLC/SSUi8Nybdg6EX/6jX+mgfAvB/qHnr8
2z+Vb5UxPUH5ZjNPtXSKTNTFxkINusa7DU2gl5TLIDcLbn60SNVbP8xec7G+QH0dINZYfjWShL8y
NCphf3OQQuucygCBs1Yl0wvXwFHdZLiWcv5VS48b7YYoKS2MRc2QJPOalmaTt5RuwAXghavCiJjz
fyDcM7xYbleiwiEo6nt35kX9iFHckF089F0o+M+lQD0PDQY8OxXcdaTfyeQTjOO0cVPVOdD5zOYF
yqsRCHM/TWlxDqKgKzaUuVYHpLvT3gPJhyrUJ9+v94fAuOHDtbO8Q9eheW0kOPQ0I5f5qM8LibB8
IQ5U3GzZCUmUVPFMDnw0mJ7k5TDtBhPraO0VE9JnhpMDj1PeYPz4Mu/p9f4uVIuB6Huol/Ka5G/R
V6yL2d1Ol20ONl14nXE1nk2LJRdklnmqP5uD2sIKIRnIDZuU3ZNKfwgldeN44DdN9iUpuobvVOVb
YziQm3svVBDrWRQcCJ0YptUCtvhNdJw/kk5DD/dlet0zNCRAR8gR+1O2TY1PGBX5huGOOvGbZ+Ps
XguM/HqzXSYqJ/yblyZxJ8qbYVZUra3j935x5A5VyXeewZLqCxGgzGseTMggGn0o+aUqK4CGJVeA
BGJaJYw00RqbwxN5M0Zbkb4zJP1s2zDC9LwZ0LcCRnVSEyj9xI8kuxl8rnjSv9OGxhhakokRj3FC
rSlN82nZwUj4UyC66CaWVojFdmThdI38wGoqk6a+Lbku1UoF4E3aOnAxpLqm/e/syT/TG+qNYVI1
/YLEbox4zwt7RCslP/L+ujRksGJdKJ+Os44D2PHks+LT6Ip1iPkauw7ZhDroCHulfBGny1mkua+Y
xFYh3IpISjvYPn9aaXXBt2ttEcgGfs+YODkHFytAuOUJgsFZhdywfi+wyrUXffpoSwfYP6zZ1aWj
SK6oAPtXlrRmQbRGPhNPydndWilJ7SUmADBb7z69xZf790pq0uXvTzG9spPtABl5fgIHDoQH2LUX
2bo/HHsLjDv/PCra+hnFRJOU7DaX9w2QR22k82FHZoeItVsj2o/ebFuq67VlT90Ym7p9TkVX811T
tGyesh6Y65zv24MQPffjxzNdHOYSBSaOEL8cpjokTVzSPNbOMCBWBzWqXV+8VkbdUb1WXtIi/+kW
9P04ApO6JpbhaBbvt0i15iSrVg9wMty+N0CWcwkoox0F/zgKkwSESLaCn/iQuTPkY4M4jaHf5E7Z
0vJMunQBBwhxDqgVC+/PkO8mOEWDbEoFeg/CDx8QJzxmOd7A3NmSU+xryyhLSOORYPO/PJne/jjq
4MRrd9rpAjzQ08kAJ/gHeOu+nRt3gzjRDrLfdVIqK9gCrTNQM/Mug9rJACq8z92EcddxBtSevWb0
QqEUhB2Bkf4S84IbEb0qYQPOUh2orOni7yAxV3ccU04NDAOAntM5hGtCLK068wLS5YJON8XdeOnK
Bf7kRP3gic6E0fd+oSAwTXXdH+WGYJsziwcNFzsWWmkP8GPp5geTE8J9StbcyIxY6/Cs0iM4oYGy
CljuZYsmdTsL+i+lzrZMR0gvN1SsUKDguSd4azK3Bn4eeYtpBsKHi8LzDPFxTtNGw91qO6h2BjTG
cX4m/AN6t0oYT65yo8HYxghuI9qVhM5EJUWvkwOMdvMKETuvywgBAbHbt54iMMzAdprEcfUDBSIF
timAMNDusTLxXDIWUpU3YSw51kwJs1Mt14VRSZnEzZZvnafIeFzrNpTd732UNjDpgk9yq5Lchft/
5FnWNsoAsj5cLIcu9CUrAV9fnnfjDwd7TQC+UmctNAOhcjnQJkJ1YxqgmVXyZMrQ42es/9pDZgmC
kqW6QCaviGD4/T1cW7nse96i+CAD8Myu1R78811VagTIM1/edVtun2XZ2kvP4FQTBfXm8IsEPcYl
lQbnkvEdnoYdt1QhOmO/W+0neQG9siFEp7GFQvFIMjsmvc5NVyLjBozLLO4jok0g73AFGd5woQ2w
V40RwPmqsb0e4v3hLGaRFZ7wRN7NVMQXnqHHyJWiMcG/hk44nEJ7VyMCMpHroKcmiozOGosQNTgq
Z4vWWnmWxdrErFICl/kdO3uvJJ4LXkZz5cET+zfA9RmKPgpxc+4lGMVhdkI/rcl+QsZhLyDKU6Ng
v4S2UTLlcMgbyfMrV7D9zkuMtEjGNTPvyw7xs4gmEMasFiCgzHvohLtsH3DcfDs5ITFnVYPIKDw4
vsoj5AKaXYmFQN29mcbRmkULTPLbORtVoRb2ERjvXiwU5an1Etk5H1iOfjf62cKdQmueln0G2wO4
DdfdUptb19GH8IoEHNk/q3FYgXeQxhPry51Z6QgG2a+eT0j2r/kMHTokG1s/bbQLGejzYMiQTyio
Pka5Y7OeZL9Rdg1E/3/ryLrfmZTJDCyEL0cncfCJNKmNVFoxiylzt+tL6ZPZqeNqkn1zOFtwd0gm
HnkhHV3vysVivmpd5YFmVTAnuFSIeKiiT20Nzsh1zHajvaY2Prb9Nyp1394ZW2Dhv19AGdGp2m76
joe1ha+KFQ+CblX9p1vLM4w25nBIZknWOpqa5vEU0Ci7HQAxOJysi4MYiZOLN8SMRaUVu8l8A/aW
WpiMgmA+NnwM6FlkPIkUt1sYa4ENa5ejyAQqUKWwJD5gwIDmjdUbUdnxSNLIV6GQz9G21E1TnKTC
MEAOq9LrgpksvqJ0kZ1dfPxirqTxExTMFLg4gKewcJt7tRZyban1PutnavoXEJoFflj41rkyjdiG
P06im9aEvWOfx8bRQb14bjxKbyXlaNPj0GT/fq4y2u1+vpWKtE/LUfLwDBFFnPqjjApjLi8O7atz
6to4BK4HW56quwPdjLVPL2QIrR7+vk2qXuJ0aCfcOy5EXzbusCtadAnLDxKBZw7fZXPta5smBp81
LnSPEZMIiONumB5Y4+WguX98AQkkP+pAg/+Al6yOKFGWigf/iHdCMdBhs2gnYeDTguHhn652qY9J
Rj/1owmU67azJQNOUKdBtpM0Ycvf9/UxzOUvZThnWPVMNr0LhXlbgcidWuDBNLuGp7FA/6YMCaUr
60DZ2114G9vF5csBBb5DqRAsDjkR33TE3KMFoiVvhTfe7RcFP+85yMZ/k8Q70L710KSLzGn5qJA/
04uNQDSNO4i7DY80MMaDp6E6+5ClEf2Rmj1VWqMGjTBVNSxmY65/+I02zreEm3fNXjKKN076Dgdq
XChrOB0Kwwm5hy1eC05jpwK65QqZj562L/eiufmI4DiPM1pYGLn6T13gEymr+yfZbkzhiSjQU7tk
YQRjPIiNfOs9Khnz1FxB+YEeKOELok5WILjpMzAWfJMbCMHcA8A1iA3C88NYH1xAkZxX3SPl6ZpE
ZHe6kIAJloy8gu0inbztuPGLl9QZCRjHMTbxRQmyAqul+k+azG8qdOU4Nt1cbT3swV/TVCn5nbH0
rXQEwX1m/LLsYEFgMmJ7W4rFNwvUlF6bUUiFCa0fuXke9+PaLl9JAcFt01x4oOUuR7BN9bI+6vw+
jLcgi4VlL54dCWdP/BOcJ4uAoLoUzBW8VyiZa+LF/csTylOM7L2au3R/1azbgY4uDOV62eMwld2F
/juZUYC6gZl17WkcI0ahUnWnmQYhjGxKyQa1iuOPiFOsN4osZ/nFXxQjL+AGVkGwiEWBfqTO8bMl
xWMAJ4Kf3Je2F0N2EDaKD8DGPfVOv+gwr4evFrKo7Tw+5KJ/J8VbEBiyV9mwm/tPvQtwK6kkvwii
HlZ27fKeaHu79uuHua5OhSaTLgjuVjZv2C/Vqa97wjWyYDFLi5uSjAHDgnW5poTFLPPLPcLpv4Ek
WZ48J41eeteokksjcxHZB7uD8nhuwD8AnICZtspEEh4YmibrQqmXcJnAJ/7BnBwVHJHCIOzuNbY9
53Tbg6bEBR45wfKV5lU4cecFlweWzIVeP3q1Jz2GWxnvm3GLczNt/sA3qVqvLtulBTdMjdblWxwc
Wv+o0X4B8fy8oCgPBJxRZTRQmRxRS24RTTuPXtxoPNhshTWfiEHs5qRyiG+0dXOebpGbwgCuLxst
hbFLoH0iE8hqKUwq5DggfsJ0qLEabWioFhpmV0fgjAO1tmGYDWWHBfyiIcBG6dxX/5wfWGr7yQQB
ODlta2qvPEtJ78EtU6qkW2lSTEkbp5Ut8njJ2up9ewxR+YLjLyEqIcNeUyUXvm/rb/XpPNB3rnXc
3itjc040SS3Ue9srFHz0QPvsI/JAZoELTkeBqH511cCW5IIVFODNRcdfxJTUPEv8PvrxZOKAV44G
X/c/TIKXnbug7hmLc+iOWXeDaHS4LQeUVk1rtZuV3RMsjzG6qbm+SKFB6CqQH9Z5nxjNvI1iKKvq
G0REsqKQaFcRCcRvZ2O6V4AB0D0uILHbd+Vg2jzsi7dtlX/yxIPuecGEOE5HpdJmBc8KQ/fxkJnw
JreFHBXvV96rL5mo8sNDkpBmYrHdGnjH6UgxJtPaS/bJYJs3T1QvYTai1WpFkBCOnPmRA1EtPZp/
rKwfMdqLL0xwF+dt45nx7L9ma5RmRzITHl5GocTTXtzcDdtyZfYAp1spFeg0xXWiaflyLcYKN6EZ
wsF+rh+SF+tho91oR06xieTs1rmFIckDpXAX72v1dmpoev3BfBcnPPqEYbVrEOjLrpWS01CLI5i+
0n3o9aP5aOOw7aZNR2zlAd+S/pAlm4YYJvINsgswX4CEVF2uvGL0HZ5rvOkrwbJfE1JINM2PyFR9
Hk3WDUHK8Sq99Bn0vNAF+3AYWoreHBqaQqfoUZYPRb3x1bJtTSfzWcv+Lokv6ojWl+Tga1WSxY6c
0T6oFJ3oyPf58vsja8mLEqcoN/xs9MWl4+BCRpkgQL9nqJgWjclZISTzjPs3FctZcXWvIu7lZ4uG
mOm9g0EdFV2oFpeaI47cO/ktbjtE+YsIj3cm7WCEf0yD/leO33uB0QUIbtJ2nL4IshmOICrOJDfy
Re54Ap+4m57UKF4Q3JKSLiD2I+eKC2u/6bc6Fvkcw30tq/QK4l3SDpRUU7o1LNnxvshDqc6Tv3cO
NwYvmtTQ3v//mSqeKd5dLu/c+KBdwnmUv9bWUoMnAXcLdUvKHZtPuSfY3wEQKl+yQq4leE+NTyII
rK7LGiC+yvUEFzzNeZXtEf7MC1mEc22d0IhKxv0aJ4Mkny+tgOjAGO9kKCXE9BzSwxu3DrLnCifI
sulXm6+qoANAiOsllnKXwXdByLWZvxvpxb88JdcsBdxhT3WqZ3GvniGxLsxMjzep9j1SUXB8Z2PP
F6HhGDplU1N3jYt3EjOpmfnYMVYgGf89c3Ar5hgkcxUXZ3jk/4KwIrAfAjEkhmpAbEm8pCEQwy4A
Sr7fkxO+tWww7L7n0kHmbMGnOdqZZ/Q8/l7OBVZb1TKFC3i9FsmMTsrf2afriEqaaX5idyClQxC0
AbU54t0clQBIIXj/PVNeOIwaBmeBCZOAEXEGnB6O8QclJXz4Iqc7VIUboiFsyBJdzuQ1QUbswOqx
gU5845iZ93iGNdgcqfT2xdYG5l21LLGUFeifTnYeIKSDeJOcwEzeyN82EiFfOrn3VETiA3V3+yDw
wWSj8AOFATs5/k2COYNPLOBQX74tpAyCmFHZCLNrqLLod+orqQ9PoWCEcRV/bLSYLVeTtDO3JLQM
0IFMRiPjiSuZeYTGIj81ypqprL6PjHcdqbs5r6asDCQsYq/7Y6YLJtSlhkujPI0BVyBuWT+3G9Vg
WrIu5Ak/evdhmze1lwB97C3+blpTXWmtiZcAiqaaVuDI8pA45aN6BuoACNbXLVRjiBvQmJber2Yu
l/1EVfQwz3zGPMjG61SZE6MFxdq5ce0S2a2T6cP6n82Afy7q0Wwld7ZY94uldAZNuC1yrEWLdvJZ
s2l3QZRJCezdqE6Qu33WNdZrtkwVjvmgUkA67wM7F7R1/xgVysgAlAdeUNJ0KXTxJH6E/14qldw+
RVtNF9+FtePkhsDMJCE0CC1IoB5sj8pKwMzwuEaFbo6+m7dZi8Re0LNL55096rkRzatoGXy1VRWm
Ugw9JxdL2oCAMh+oyemCckH3/zpjSypsnD63kFwCVNizOcPojnur9ZVBJM5jL2e1DngkVlYYUm3B
E+95ASOhzgqOc6Sxhwp4pKfBiuEIpa6aa7NKbEAK9u/uWdK9e8qVtUY2H78TTJqxeEYZZtieeH/w
1IVk1V+J+fY1KOphNO54LVhvkV1/t8Iukx9+aCw8ARHgVkt6Y/wJgqoJKUzwOKMSD3Nd+rwfWoyF
PvZWGe4KlpqsfXNSe9OVDyoIXh3+UQnxnxHJvq5xHLSSfCOyikgvWrLla/H++alZWFmfjzi2BRqH
n/kgK88EnuAAYHbog29E8eipmq/QBaSuOR3K/t9nJst1l05FHgb/roLGGS8QRdRy8+KR/tt37dom
1XgPTDOP4z2j/CNW71MdqF8ncpNmOAGvogS2O58jGrikqc9+Xva4nvAVnuSNBPHsQ9kTx6syXCGG
34BQUWVhu7lTSO80JIvO45hebYwX01vYtIZyOw5rdEXZYgsjjzIXs/qgWHAXTj3RWYoFtuRSfF3W
jXvD2eNvHn8ipErCks42ck+BKCwXfUu0Vn1qS1QuzqINfgcQJxDeGLD3MNtHpM2+H7r3lRRByg1D
sbNuMdOI0jcUvkIcSQ7q84U22htoO9JJ/uLkcLAb9nRImraD2sCxvPmUGvFhPtJAAQpOUImPXU1P
iPDnyDUYfCgJtpzjJln23BTEs8fKvjFDJzjKAKLRUl5oBbIPPc4SBNDf18UOvgJ8UtE8uGtcYeRb
SwuetLRCFcs9I7iH9RQO/2bR+Ni+m/kGDJGoJMAtUtWLR0O8c/YZOF+JFsW4s2PISf4FeeqnNFtl
1PH1O9u31Pyukn6hdSYjQLKpOpx5lClm401UD+RC649g8LUB4aXCPA5dMv+mmSJr820hudmypoD0
OYLsAW7318zl7bEcoig2HmN22ICgHyBYXa+77W7QS6wOpO0kelfxPrjqFXK2N6BcSXGC9NFFfhl+
VlPP85sUOptvngTY2K1HOX0wnwRBtJJqm7g2dE1BEOxOiqWMjYOUOkxq2TBPf+1Q8MNgQD3/bJzG
dINKPZz7wlXwX4dhjLhfKjsLsw/OyrkX7YzvHLbtjqyiMI/Re5bDVzNNWRmNQtKOrv2Ndyp2dfX/
dZVaYjFmcGkC/I6ihcIZ6fX30lhxfGgbLVowkOwh7/ryrJRBQECiCvgOpgW+sgoKJainwKpzfIga
B+pa0wGSwTPDSPF2uKzLcluzUIFN8Usf4ZF1roKfDtesfuPrrXR2kgVygQHp4mOrZxhCCqAMy3UA
vYraoCvyN3lTzfZpirvfNVDEvRgRlQunkCtFYWtazSk36LeRhlzThAVSGkvl/3FThPYtG0pXu03Q
FLqQ/aBK5H3guyPBl1vNRUSORo2bqnsw3YsL0QYXFd1+AR/PHMl1htGpF7BDPQltShkvS1EQjVOs
SLXUwzaC+rMb6KWHJAr3V0SryRHAhwbVyVXxAX3IUOIU7uiomxMxIZcAlK/eZ4DzZDPZy5EUR+l7
NgvmaKgfQmU+hSLiYIhOu17zaSSspff46pSf5r5+ypfi9Fuzy3ykxR9nbCH/AOk5KaUxvjJ9O7Y5
uDLCgCwVCGgnfWq7PLAKGaMu9BqnCWSve5blCpHv1nMdgT6/OMQIaQqFYtfvdYxsc2nLf5YRiKlv
e8HdKruwHt1EGb9H7eKgPX9nE3iaE9/5KwBCKr1bYx1t85SnVubAuiwGvE8PKL/uGJHG+vdOeoAV
TVKZKr0FxeAllvfF+eBrmGWWOSEbiBt/42ZdimFy8LxcH1Nu6WGHgmV7SVoOc2Ac95ueYerbjz7X
iXKwzmBrQ+6Nm/rnFC55HkFE4HM8FnvqK7bE95RM3ApkVPINiZwueFvDnVv9bcjvDjW2Pc0IrbxW
v6Ozb1YF+9I06WfI4bS4ZBaUnijhPBoV9gt2n9H8zqmQ2AgnZF3c58wL4Df/QYTfIi1OCH6+k8KQ
AvQNDjJrEQlLtqHoy/aJPPo1Z8Vivq1C5TfU7pshlL9Ow2WGdI5l+KsGlpqsTOvmzP3JFWz6WFji
NfFprB6e7oLMbVtPGe9uZilvPiSq+eLTuX8lLLpZK1yj2IrCDtIyzUuVwtn3xVgxip11dBW+YqMy
rbWEVnDWXSn/FPmCJDEVOmyTbZMRdJwFgkwVPf/F/y5wgRvaL0kg5Ce0LG/5RXfLo5vcJrJHWsa0
PPYlSvvdtT3K8QKcjCCU2ESy+qujsZdkw6H5bgDI3R6WDWZy4ad7TKGeV3s0srkPp2zDjqSFONek
8Hb/pFzlg24Dhwa/lzEYqERv4/i+Dbjgp/ILQnbHJPH6mA59BlK+csEXBhWIR9QPrlYgnuidoE2D
DwpnzkAyLdJ3wLnpOBWAP/2194g8O7y/buLh0pt++MEEw6jf03Y0h6RdsQQa44MQxIgg8V3tPc2h
waVATm7rhrK79GyEw4zg9+s6X7QnF2387uLE0TSXc7j0vwLhkPR6e0aTuTbynd1WfC8BcE0CNdIH
TUs6JsG4nzY3HAEESNATsAUPu7sprETNUrVA8aEsFx+Ythvt6yHD+huMok/HRGMFj/fyKjX90MB8
yVq6Odm0I/0YiajuqGePCugKFCBaHd2kvbo/wZcu55oc50XDDofWlVlLgMZFk2r0fC3G/qqowkat
7tXgIpGHgvc/5MINXqM3odnniioTaFH2XOq5L7G8Ykh0ugSVKqhXAfiZJ+e6rM/tCCr7chaLAAXc
g6gKW1H+skugwa13PojPlmBTjoefABYpSe1dFo4nq10ORpdvrXFtCWU/q/sCsB47V1S/etyOKBPx
UtI78Kd5uoo+d3VY7wJT5yhwJNBDOm5Oe8dA6A72qBhNPOWD2Osan/Eu8OVibmINIuRNl//4BrF+
J1ECsDdBiBp2RYJ1gtpATv0PRfD+MpRpNf6fFBI/mw142pO6+z2b/UCDQpZfK5FPLpB2Xt9DmgNV
7XrBnw+oRdDJdg4dyu7NhWYn5tHHBBlTdOcOwmj/YGxxGUNLf0mBG3OUmlcOzbnRkdNVqkhyHGnK
8A546YLySZnwacUTOKVU9gFmUzkFLLKjfGizMUaoHEK1TAJVIufV7QtNK7J3MGJlctQE6I2HEyrt
JwT+ydbdbB1blEOxB2VkRz+pzlvTIMSVA4PY81sqYIB44z0COpMxKeyjJRyCc2cEdxKqbtEz5daI
L4i/LX6VnkrPP31EsjgDKacpSR2GNcSHjg2eyFBd6Jfu4taPag5d1n9KwLStIIiYqHdTJnTLEARv
qLSeaq+yoef203dEdtiasIKuzlVIMzCAnXu9tFOho3kRvhMbJpU9Bp7P6JmLWUCQoWzRHerSteNq
Wt9xrzUV4n9tDSU4iRvSwYfTpNyECr2XT2PJOh5RHVEURKBW0wNS16A6OwxrFVl6MV660gdRoYAI
PECrGWdpYY1DiVB1ZmPXWWwMo+XpYK63/cqDG5vuxVwWwhz+qmjHkd2MNDDqB9lu53eir6XINy/d
BSy1rM6nj1WZexiz4rLrX//XEco/arUarFC/ZpnrVAI45IcgaQHmM4uPc8Dy+RWaX4psafe4//zc
8mIVxSH2dhQX7CsAWK/zmvVzWaJ2puckOZ0elVfu2nzbbUEaZVzDIbUn1E8hRsvyFYiPY46Nh0+O
wYjlQcZSx2Nh4+1C1OREi6UaUqGDzpZCpsHogOrSHY65ERi3721psS1OuA70KxqYS5QEdnLcOTpK
6CyJfCPlpmpJNDArsK61289byp0gOzy0XtrOztpSBNEPXXYBmIoTsAQ4CdXEnwRsWcZ8WkM2Y13y
wSJU5v8/CCrFuoVhrc1ksYTX1hMiGINZjz9GZME8Cbj+n/Yo4aFDLZrlkbP9SM/R6dcIWOe9rdcp
D6aCQvPksPLpJmqYG6IqvTPtd1t9SFhItoxPaAIEW/GCpqaD/0Oaqh9mlZ4qA+brhD2mofd90DXq
l9YdLVB3HGBdgOda91C2FAVHamcNlTTvN8rK2MMgIjcOUAcR9M9sFCCtLPwSTPe6EUV2sDkyaukd
lPgd6FAU18uzviw+Lzpwss9RSupgMIoTgNEGKtBWJe1fukhKUBclYPxCjIbS1bZbt9uswT4Z3sny
7OTWYlPUzM1dYJO+155DJ8HZGUKgWAqRdkMn9yo5pGqSiVa6DnbPC4SeqWcVTo3a+2UZav4jBGnO
yXWGA+D1AWNQ7WfL9Tv1P1w9RwCYiP0fPxchky42i/TEkOZXsVvfydxnmSzizUgpOfn8t4ZiDJRw
K+s6P6w5JDXWytk4p/CrkbT9jcv9T8rAYyIp40ywNLWTzSEyILOiDPpgo+5VKBQQG2zPHvfxo9S9
R5n9msfbTFcHT5rzZ9X3bEogiWB/r8Tklugii0dBLAx0DTBu+d1N+Lrx/OI3hTjxCXhrSqWaJuqQ
C7lIB+RwaVHQUEfm9xCXdmxuYNmOmtHYCCF5rHM27rvFlW3oxbHo9MQAh6AkM0WyBbGY84zWXnJy
uFpBXtDfgrt0L69dsCOM7evEFS4Q2PeUlEzccktqCVicPKvIcMQ/zbG5JgQW5FbPrRBCuBylLyCl
876Id9v6PUUXGKJb190MO1U6r9D+d3yN4raolW01jtXxv3WJponQ4bWPFIxsbWE2wA6ADW8FwCCh
XHLMGh4T9OtV5OBTLDRMLi3zsK7l9lU2917U7Zp5pZYOExugBgvHsKZSzhPSsghT/UvgtW8Kmd64
p9/QYwoDT2gtfNxOKKSsXpA6UVZ0VGmIVIvI9qz7p738DeoB5ual+OQe9SVWK7W84hidyExLbE9p
X6T6/3vX1okQrn+acbawqmTTquNgc2fi46iX5zDeIFvvnxEseyPHqtvX7WXyikEdQrJ7Zpwb5wPU
sqmJIPzGBhyntkyNcTYmk45gZvm5hTyLfxUOuiwu928M4mRcaxbxJgYFtg6E97EeSqFQv8pvfAWF
lpDwTdZXSN8MRUuVsEum1UHc6GM/gJOqQIEv55R4SbJtnniGLpQu4IySSOrl8UlEDGbZUT3j7m+n
h0LX0QpM+Y7sqH7boTEkeIcwhbwCMu9b6WDM9Io7CIOmrvgjsPba/bnAviEINngz5GrVycMdkWfX
PL+g6gQbQRMS+1ZV4IupnGHmbu2yL7X9QB8vypoV8Wh55WZ6uoP4NqPDzIWDBfOD99taz9n9rDGl
HBctx1YHaNDSiKJl58bB7qjRvlDmCj3dRlxLr65jreqL+ONn06UKv+3tmsjH3LICe0MQUrTB9mwm
xNwZj7ywXPJo2CVdq+vNSuID87Kb5tr1vf9cSfKu7WBoJgu4VizjflO3xd2YlNGK0jYL/Oo3TF3S
I66nGTRXf683mDNq214RhYiwlA48QcGikVIVQCLDSO+CcMJ0gDmCi5SIVZIQQVIPru542lAtPDYg
oxXtYWzh5T9MkfwokhTrwqodmUmDZnSJEEUfYDidhoxTAOiwfEVirzPjy46VDqtbzKYGx1WK32D7
3VuqWy8sWsys5USeHJOfRi8D8KQ4ibLFjDVGO/U466TGAfDmKt1wEC+0gCBtcyCVRiAcyCS8yoaI
LmL0KtIndWtUA7L1IxjDUgLsHhclpJL8BUIDGuV/fTs3YtCPX1FfPP8VAbsDNt4vctHhz4GK62Xt
P8VF1IrKulTTXNBsOoIAhEcKCuI5jszly71yf6FhT2Fq5gzMXZesxYyWnON1pHuw93LS3y1zAaZN
KKPYLUBvkkkKnFbDFEi+WOWHKLL+WmJVBzkFqRi+pX7FN0chtCvvR3TkyPpOrshcnn9F1vmCMJJn
F2qA7dwKFnWAYdXZUYJ2IlxXOgXE9JXbQFWqRUMpIH56cbQ5xMhJIODi28l9eP6ycROgXwf/5/pI
L2APdUrKxCX0MLA49tjAvX49n/85rkCZTkJMKiEgiJRGhCoe86VjUETIkz4RLO53fR1w/I8Mxuh9
aIPtxBy2p/KnTNzD29QmD/oXbirVgDzU54Xd2BP9lo6yX6ITb/sljhIVRnUu0zfecLBTrkezV499
eQN1X8VdVDlGms9V5XnwWl04HUL/wqQ+lMxdWuqpnQOkfsiL2oPshhNcTSK6wXxXAX1sx/Dcupzn
/+0TcFiqAau+PDj8d1ssODpVJr7IFD1kvvgXEfq0iejqWAtVlzPoAE/nbHTRAVptOGYtwHujqSuE
rr/004Zaf7YRZ3wgRVARSK/tJ0Op+y8xGtDVQaOKyOQ7Q3nNq1yBIYirlYQ7ib8GwRU2UMfbsADx
wTeNTZum8+ilmrjudykFghzKKIfNpMEWWrtn3+IBXGfTFMt91YFfEJRGif4DczXHK/FTT0lMhqju
Je75Dg4RpojIXGiBy+GR20tK/Wz8DdBTVgk7IYJUfKNpl7Ik9aKAnX/dLKsmBFfxy5+QiAGt/keC
jFv0nRH5dAsp3Qp9fAat8mH/gmM2OTJQ+um82TYqsbUSO8k6w3G1V6wtvjU80kp5sYVarsdd0kxL
+2IFiJ5UDzHbRPvMaTeBL5Zb81UfJeOzF6UbGxCORJGS6ZIKaGjRGL5HAm14f6dEXgYezNcDXCQj
kMKXSd5MbJEoAuP3Xdj9tHKMY3Y2VAbSKEqRjessdVZcJvBOTAoA4rDcUGuA7GBuKStGPpX3rqKx
GfxvYHdMP2NGY9Ump7IqEB0D47cHt3Hef+PoZ62h6yUSTmzYn0h1546T8N77SIvrqWhFKcYvZdDq
sbYG5yqpNXJ+Vw9btQe4pRK1VkqYp7kZMSiZOZi3NeWT23Hlf/yLGrTXd4LV/dm7UnapSthIueJt
7TfDVHhcvRebFD4MwAQpsCuo2v7TpVCqitk1cf2H+zmC5dnykpEkP2z9KVQdTWlG42+r7vHuQ6jD
NZTRAnjmft1oXqewN8s0agMwBt8CQLBKXkHekFrkmS0IZQU4od/UC0wqnbQHndRPH4IR+/2BCK0t
+2ccb1spWItnSgRIRnt8GEFmb/WqZJjAit9h4UPH7Q+KtQlqsKST9d1JHCr9nxxkbX/tdzgAOF1e
tOQ2mIAg51KxvhRoBeYjYt+6DlL6qoNZY7npDau8HXGYRam/ac6MWPEYMiGruLVQec3LP/VzNqMX
d1aQCNkSTGxWUC+AlmPE8RFaqCAgX+XlTeFlbyK8KXwhe4XR0tsmDoYfY0RTsYFUVYd6UalOGRL2
AHzdHm8sVKtwDk+vIlXDLKT12yMKlF28ZIS68nx5GI/jL166MGOoCMjR+AfjCrIwt1qF89COSV5q
feMUCQ9JIXHFehfmQF+KicYJ6qzbjlhXE6kIcgM2dcRyCf64GBNjRoLaFiuKliqfBgKSmT2K6h4M
eDqFyatnl0f9vwBSUg6DE0HD2/G2Bd+dlmtE9iYOAB8HJ3FLf1Z040j/IRkyzmpYLAYly/nBQtR7
9RQuZsobYL5cr097O7M/OfVoD5VIXs1bPbikHadRv8fP4rxDTL22l6dYbc6F6HBkNjRN4nPo4Ud6
4BOzUofmMIR6LjyJXLryyRHYVi+RjIACccIeCooJxSbZGH1OXzzOrpRgnTIi8xHa5lN6IEeK3ukZ
/y3QeF3C7eN28mlJt9ZKC0NOUkHMpSfVx0gyfGQCDsO2C42hoopod6dpwa2JqefhnTmvU+USu0dl
EBpPjTn5QD4rG8uz3i/AltmOYpg7s1uS3/ne2zTAFJvw77BUUp9Sg5AoWNN1w5uHlAqkkshYPGWm
uTF6xiuGdeUl3Pqrl1AgYGg/dzD0AlJLO98gZzOC8lwKnUWnqLN1Ul9QFo1cG7dmNiWZqY//5bHW
2SX1l/D+ILbFC4pPAYIovn4JJHEsB3wbcCEqyYZkldcVFs/MuviigeeQAmBqnFDRYAR2cVpNrEG8
tu6xqpSaJMhupQLhTUgZJFNq0ggNQbqlepDYtUFyit0+H1t4bE3QO3l6LEzBvVBD8XYZMykM0LfV
Y+B0mC9hayWLTQbL7wObByObaWGU9fya1GNI2XSwdF9PN7P6nWXtimB2pOM5dcOazWV/IxApyx6u
idAW+bo0Xxr7qiFPXHruJHmCEWFCT8WNAc3jM1lFtGqlydpelwKYpdHEYhP9CxXK/S0sK7xlrTjR
bGAnT/wb+yYwhxKQCsF83BQW+jhQXHgxsT7/r0eBEYQd4oVcLBjjneToR2hQIdhaTHYBS6JDZLlD
TVCE1AnYWOiMdg8ztteLJRj+e/OlR9HX5OL5U1AwJEpfBL0Q1+Q9Mh4HvybydGQUuvCnGHuLdxTx
SIlSaWHsnJXaTl/7P6Xb1kkqpHuSs4VrG3CMpnCJhppQvFiqPDm10BpIb7lHGzQyggVlznEBb2xp
4ndz3sUY7BMGPOXQfN4IGbuXahuPn5Nhi6sYDU3Vrx81tZT4mTGNR+PmNB6rQrclhfncdBTl2G9s
Yg0+UlPbHZvfAAvg1spMmd6nlksh9J5pA9nYwvYWpvOLj337l3ozNEoSOpDQBSQOkAr/uGB58yF7
EHwwF7liJgFNnJ2rSDL7sY8cOcIlSSrBtKL6o5UGxkXQxyPGMpGeilmtze4/walxW8hTXJEzwf/I
B+lTQ2lHzPSmltEWty24QSQDhh5oP46ua/LO1cQYR/REs2bivI82Wfpb3AJMwgZorIAj217VQ/Q5
ykcLSpBoRF02VF7ec48tjZPA/UF0pocB9NejJf9QxvDygOdvH/poo2ihtafTlQY8Qzg4wQxFQ6+f
vUNXaMyYNnK9OOtbMPHzHhU/wlatquc+rHuHsoabxSaAUvcCLBcMAAyYEAQ1QOeuuUOWvTmKwCVG
OtQFj87ZB0aVYIwVAkTT0kN/3h+kbQehHTvdeIwZpk1KxT7fUVzNppRm+wNEpxyNf4M7l0wfdBZi
FO9C47geSSVJS8jK7xN+OiBYFPQkcG1j8X8n6+3FwtukkWCayog/t67NxI02dF9PBvMin8VP4puM
vPldOZsrmmsgoYXyDwycWmyH7uoK9tjZG9b+maLUBDSF/cob/xi7UlhL23ljAxpn9lSz766DqjAA
dQkvIl2U+kSQXLyjB5Z0bytsrOpLDsVrIDyvwvvbToiAFl+gso+uRuj6BhBSL+Z9MWv2Ikiq202t
/0A7Q2cjC4wsK27UYPfz2MGy48hdeXHo0tuilap/41xwfh6808C99JZlYoqClj+bVjjHDsjsA/Oe
Mv0hVrpopBW6XqA5cVOz5D01McCLgUKtF18RF0oRKp6r0X554mwpvI4ppMFVDySUwxiT6TKmiljU
DTl47dS397BKBs/F6qWN9I0sqqNCSraj4VzQiBzjV3EZB45C3qBT97PgpsSMTFCsIYh8IvjSxSnE
uHHZ45WIZqFZRavPA2xIyGeAw1avWSeZ6uXzcJZGh5umkCaBojR8Qrie+kIgWMrUVk0NXqzUQMs9
FGmbsr8ucT9P/YTBtpRVtyf0bogaGov5tsT9mTOYG6tPVZLmbrQGiWW2OQZx5FsYRG+DzlwRo1gN
gs2obKsAthTtl4uBl5yACVFgybbEqL6YNziSHvA/tfVlWLzkwkCt08KokGrZiaLUKJZuIjqviRfz
yeCTnajBLvwutfpjKHbTET7XZVniaOHqF+gSzvy0aMFHYV3N3rho5aCK/qegJkBBWs6ZK7EwL1Uu
dswA/RElRAlD9j7oeF+BBZepR+L9hbaNihnRFWeIvA93/eTW0RhVacGMJWY7elt0I/uW/y5C9HvY
ev3UQFoMCj/e3sKyZ3b7PAEKkFh3op1BTBi6Udjo6IiwSLM57wonMRucrz7qkRbL4gvOZnLJ0ZgW
yDXwWz3V9MyaCqAtgrqMVbO8lbA4lWqitlRZDQyeQ53Pya2MiVFlKSjwAcm3YJzzOT65IvlcHp4Z
zYyk64XC2gDBW01drcVhdmVRTh4/HEc2OEwLua5Oa5gW7xsTNJ85DEFvW2EAcXpd2X+P+6QWDXvC
NlUix4Z3mTKLRetWJlDeItZC2KGcByCOLDi3sk/huNJkDv5eG6KeJW+znXalWkwXVx5fqdxFMBSV
PgKh7u8zWsSdX5J+ZpvUW3Fn9qCUn6LYV0XJG44vX0tCmjtcYYh6D8mgmDogWZ00pfInkUeQYo3r
DwuuRMpnF9WIhyhdDPDcyfC3il34XnIwzVIvwRDEzQjdShO4D4i/F/DHjkeDs1o8GseoGbWn+uXD
IYOWXVYHMKQylbaKpZ24s1Ux3EPrfVE3dRrQusuaH3FPRtmnxDQUtTjTcfb6GKdpPqp5j8RagJqp
p7ZEpm5Q42IYnWHYtsZOV/5Ttjf95IEs/Y1KHkVH5vEp0lgsNUoriicCRHWd9wb4j8TAMVAQmsHL
HPiDKiHVu6LoaDWbOubmzlQ0COLwwvqZ6lOWNYhRdowOB+zoyS3c9Vo85G0NqgpP/Ra56Mwm1MPx
R+GkIqsU7cqTQog991hzWwVGbFOVMD7DeXxPhLO0HGaFwLnREhS9DqMiGfWozM2h6B2vRgAWk4Rg
14x490bAedezAxclUBCFYpVCxq7BcYmA45O3NT06+vcJ5H2VCZ3DCezpwSWB90LKMGenlxRNOHEE
iyzekvDbIvXEeyCZIA2fB8xmEEqsqnJn/hZ6g2Tz/EDizcLDH0q+tLjDQ33BwkrjYfjHcTEvWWaf
v6/a9L0hZoSB9R9t9n73SAwTkwPD9WG+j7at5l8VTrWN5MSRLp6t/JedPvoR5g58eUeGxH/EV106
44AX/xUgll/oS+rAQ/5MtwH/yg6P6PGw3RSdlq597htVF06V43STs/GpAJgPpclXkBfAiqf7kfO6
EBZ21uzxI9VEwNfqH2CC5U6ZiBFPqo+akp1eJXSFoNJA9IKwVX+qAUsMNuOTYkwzN7rkofAA+PtQ
T0KKiE6jfwmm0gih8sy65UxKYaP9njvyjGzBmtjen3Y6qXbP6jNOlgNemfccA6wJSVpD7zdvQmzt
oO8x7irQ7+dG6HgnqZD6sAFIObuEmfoX2xomE/M4yAGVXyZBdFn2OfQ39oaLXpChHqHmalobWcgD
Btp1CYkDOQubU9puADNfCQY7DMWzDhwC6DBW9wyHTIaF0pRtBosfaZFMROcZWpgp/0iXUGmd0092
lrN4uUImPxe3xZkxDsrZ/5i/fQ+5C9yPG5dSWhQFXhzFWSTKpaEMkuBA2DDXW6YkThv6n9y7Cpp1
sOopVTfQDoHKRiBlOXh0P1uH/E9XeN7cRsnb4nZC9c5RnpzTVTXrbHkXQfDSNMC9WcQdroSKMlqJ
6NdIa68bnLHHhntuqaizBmQdeTEpbqQWCphh/Dq0Hoe6YH1a1zcMFhJx3R7ioYI7kT/1eNVZiTno
ZIqFK4jGKr+9SPAyR+e0JpFSoUMoYTGkczK4jYJBiiuxe636SSA1CDPcJqegoQBbJ2cPuhJo/i9Y
8NAC0rZR0wWRCa/q9P5PnjMC3GqzU/uhOOifjA5jBft2AKGfM8EC+vLOY4joEoX6AGITRFEFzLT+
hpDuuHgb2+fjF2XN3WK3v/KyYcp82iNDOSVPUj7StZKkuNzfWrXuttYOOjk08QM3J81dJ0Obsq0Q
AJeka7FkWsuQ6dq4h5XYavud54CyNFei++/8/uVfQH3iGuKVS82aBB0H//oJFjsKpNoxtNWZmfOh
ayOQix/B0eE3FgpJZ0CZwmIyaBJfEM4I+1xtB673tIQZtsxPuVNmen/ucO2JualKmycGn5U+QwnU
jGq95jpyhU3brXeDHj/VRYsbdmclSXRQj5w0pYEdjPh0CR02n+Z1wEa2S1Omq/mHJif/5TeVwW++
+tWAv1WPn1mC5YYf1X8UNC/m54vTljzCbo425TYxrRTUnulCeI2yUEwsIJUsFxhR131i355YO7HO
u4U6SZUWroZlDHwc+c9v5N7UeKFN5vxSB20cW+YECfivmyq7Dnv0QxTf1FnpnliKrpuiauUjIpoa
0NiY7npaFgk82r2ns/H1QbNOOTMl3EgPcQeGYurjSEjdAA7JE16mnpCTYNE9IhZnZ59q8oKiU1oL
KZIdssqIPXEO0IZ39LLDeUXGgKXpskCnHoH+VmEiltEkuJALbsgr8DNYv/fNOJydFKqjGfn1JwVT
Q4ef/agIoEe5W17gZCw/YKGcT36MIRsmVuqnXAoY8NvsngJkDuI7fAuYBY3hSDFvjB4hpx0Gpx0I
QGGNkYUfM4aMblQOpsdfA04x2JbBLhR4IZnpig1wACcY2Z2+GrZ0WHPTjYpb8QU8IQKd6w4jtiKO
ssI+As1t/0ecF9R6ZUgSCrxG7SH4Gzq33PrlfUvVMO9+d4AwewMC/B02gYg9vF6ugn68BJm/Gwwo
eq0ZUYzYUgvc9MZ00yw+havW2ct+jY65KOm/PUQ/F6ZtgXHdqcl0Pe+CiKyc6w+ltZ/ydoIS+y5M
a3A/yjev8GgW0Il+txndM4lKhMIN+0cLdnZbK3DqRC3yWQWO9ov6wmYMFLkH1luZxU1SkNxWpFtn
3+0bG3bIE4Xh3xjXhibuqqcxIUCiAzHhzoEifnd2WE1PNI5V/uQQWMsGdryfScSGSfEH0CakgScS
MRNXMmse0DBlPesz8UEfr9yW1WH9XmdwEtdqglAIEqQUlbDA/Tqhioft6j7So5Pm0deXwja5MPr1
52EeQ6nKwYIYRQ32ZtlfJwEWrKQD64x+716vVKX7fIZEwZBipPDLMTMVYYzu1WcGJ3BMP6IVNO1Y
xIWoZ88s5M4lE/5IkloZHyjdKMI5TadCnYFZ2TrmQkzD98gz4S/8zv2Ih+dvGANYjtYaDS3DbZel
TFaBPFvoex0lPkXxa8y6MGZcSd+NtQDaxGWtwdbeUPv+j3TmKuxwqWCuZHP9Sqh8ZqiEjOyMrluG
v/ONAY2iR33gzcwMOiLVuv3m2rk4h7N1EOHzkDNhEtVf5aiLmFI5UGubqD1XNICL3RPHYoK2UZef
MoX/B2U46lo78JQizTxMlJCfqYs9ID53X8rmxOjr5JSNcc9wV9oDDpF7/XDfsRYH6YDjN25qO0I5
ds9hYizks61pQcp9hKHlbxUYvCU9+og8NYdbIlb0hzn9qTv9g+5pbiT6RkCUK52GpaD7HThyT09B
bk57bQCRA96e9WpiK+AdGR+wzXgAMjcykNqXOPjcpMoqwOyyy2GuPs87cIU0EV+3mMg1qxl2pfFx
XB7xGLDyQtAawTe6dA57C5nygko3CCOUA2pn6U11NXUUhavfDPl0F/CiRPdLpls5LuQ6M8SZJIA6
bn1K13VtrXlZGmOsDhP3GKCAokIKX4nIl3Y+ZLJ4XtaFK47o9mogHXuOE7xrssTQtZxKES/YlubT
2z6kjPr71XCGoX+mdloikcyyCoqoZ7yo5t7NcIHI04m+lgCZKLoFwPTs5fGnOTIIvG33LY0KJYLQ
wsrXUiBlBX7FJJFB0HpA0wqVhHzgv12sAVGdu4xGRVPAq47Ihl1siRqBQaC21QPE23bI5Oz9TKQ7
5N+mZsuemBJ7daWUUc05elr+gKp+NnCAD+sqQKcNrnFk2eEmaqedlpSgWmTRgEaqH09hVo2Vjw9A
CXt4yV6YHt8MbK0uKvZY9ZuSUhx5HyEJHgHKfUBTKv9GeI0HAl5OaA5L1AxaOnsBnQp0OetcY7G3
QwKEVoEo2g9s/Nn2UH16W4P0IxzIMtKnuvHVJeTuiVurwqCRZp485rW/yH8kHAbyIndJpzfTqsPq
GMBQ8g5/jgflZnU5FPLC5rEsjC2/ckJsr2bljJnV13uSSLZcWsawEFgfM11qroRqKHv86N3jza0R
YuggV6wdrQmfG4N5BElHEh+qOPV0N2sh9XXBYMgIvAQpkcxSvbXIeqku64kPed05krhlN+TWyE3l
ie2E1OSlyrIJrFVFK/CD2c/OETcDKS9znFMl0OxO+Ci/J4+tSJWDyCrbBM1FiRxzqO2DZdr0t3ve
hlo9mtEm/CsG/DTTrIrfssoddpGQsR2ckd3Xbyd5SH1OMUeLkUrch5L5SzYkNSCYcB9rPJlMcKwT
CS9/ceSfVcZ75o9qugmaOcl433BVmsNWxRa9P4s73kWfKqjZMYAbo2SEqphSB7VQBlNY6l3Aqh8o
oSeUlIpvx7bYs6mL+tInSw6mmU09TQnMB366rtKcbaDjUPD/L4oHVsuZt1gQdjByL6UlD9kgc65f
VIlOb4iWpAEp8NpPaxrLGY4t2qxOdkk5+Bah52Tu9DTzPJvlrE48TO2y1Xq6zfPvspzmcQGFneEv
RDAY5RCHQOMFBOuP0lY2WIWhJxoXf8cSGjcyozSEtzWbww1f6/nEk6fZSOIyut/i+lQFyXzOGPDo
aTk2Lxs8d6PxMARFscUe9p2q/HxU+mi3jr5uKpyHS7y9siFOCkIWqF66pPmiPTnehewduUVH1DRi
CdVIMjgrKTXQF+GUw5YDUOxqpH9iEhd/jB2n9JsuNX1IcrWgsWmbS7TZs3uHsVdEZPWAvIt0vwMv
udpYGMDF11tv8MWF2+l7Fm9tght9KMAjqFU4YoKzUyrXcOtrsT/Iy5t7MLMhIgEVGgu/tGYDpyQx
8uFMqpBkRJF9V1qfjGaIPcwxVNGL1DPUg8MUMaHGjkVqEtFKr0TSxPnhCY9Z1n+XOs7SRMV3a2ec
coAS8nZgSOQkPM0DR1flafUyI1xZo9EfkPJPYjwIUpdOxSo6t7IBo+NPnDm9UoEJKsbmgOGwtr5/
1DB6KE4JKh986fi5qkzUO0lfF9QiIkzOZFusdaai+0mFJ76DzKTQVg9eNYB62H0lBSBf0gYsQBkR
kDqnMx/wa9oJ3XRHZbxLpGNVxuRsoBqi9sGDB2EutYdcuaNm8R8tzcVw2If9ukw9AJXNK+gAKVF3
l+WvPVFiyvPlirq4MKmE1hMWdpl46DQD3qNJfrtR6rhsrufta+FSIxz/ItYCjDv58jP/WTPzFXBJ
k7yJlKRW74JrYjeKnzkkEbMWrolhI/POQCK9Udv7H+ky9P/3llbc4v5+vbvH/hkWKrYS+1LqKr9D
auDPNjauzGrEIXN3t66tkWN52Q7dTG4CcrnHiSrijtNyuS9PZQM5gBHT/R/5BHzB/ng2I/OQ46FW
dhV5ru8PJ9gQCv1r5sDICjwytirzKufiaDkbdkvQxZyGnqpt+dsiNHSzkPS9VIrl44EMMEApLHCD
262pO+5abggJaE0QIfdSrYv4gXVNltOYfl66ZiTrr9BOwMc1WCBf8D+WeMGY0JjOKM+zsPldTZ+A
vKPPMCtBN8XiUe76w1yR7cfckG/KJvh5IfczCO+IT2WwFuzcz93EvDHzxRE/kLcuuhOfLIVdByUK
f7a6ADGURKlrM5D2/FTx8gM/hD9Ix0AA4GBUAHonulvCdkd6MoTDtrFOSw0w2PNj7ByWtragLFUh
lAEivtcbUID0zJROOhT/f0SxMZVktdSjsc29jO3x4EFONTmcj5zkZoao4rglOuwIl9kiUMNufY63
LrwZuyIWTAeCqjc/KM0H4m8nS0kqNOqpviBvEFDETmB7EfrCpz5x5PD3RxHtEBJO18RMjUOLySuN
dmc2ACWz8WQbkkTwuEuzLkf2TmLg4tdBk/sriaDytYs2p6+DroYfuwgHBRpr8K6BTEVB2TRCjZIm
qB1E7r/FA5dRMQPwLKRNvIDFONb/0I47LTbCZSYZhtE4M06nBParO7Gs1tR3E6aZh1en4JEQf1ld
sCr+PNfmkGE+KioXFM5c9fRRxmaAc+MBmVrkNYZ/421t0k1b32/1kbjH2GuC5uUwsjNO3TQWWmbE
Wtnn+2xgDb4vBOEbpXlP6uDJiqBxfG9+Xr9psxvPkzJWcCMrrC4d484eKjht4DYmU5C3ZdbF2kRT
DW5SibLsP2N0f51rYKrz7R87M0vf7OpqcVFF7iHP3hJOsnzg6FdHC02jKhkzYaIyP8VhLtD5fS5R
5y+kfF/VYXTxRqIkyTnWGcNtWrumfiOsMa7m10E47STsx3zW3wbEhxwFXRkYUi40lMWay5vbS0AH
0UQcOHPU6AHeYU5aMQnZiHANq5uRpdZwWZuLhaxXpy95faFlmUuoV07ZyLQpjCKYD98MzGNiVF86
DPPH4nEV/qyiNYvWnsWhwZP+gSLkJDYdVEZhLkfvpjcV3nILTissrq+pl4ZWwTmDweMH14AIvFbS
lJv3GM+4+AhEKCIm6eMVJ8reSCsrZfLWKB216XFNFWfCaMuBJLxGq8xM5lEWavh/bxNmrBaDD/Lq
+lwzGSbTXHdhxaawWa6KzGisbXKKzynIhJEJvOcZS8n33u4xQ2yOS97bzPeCzT6iTFI/DpWUzdMf
aVS8v2qrX/y3Ng9fVHX14QU5g+Ok+vm6l7YInzOEp86jAEz9QiSYpdSuXUXHShegkN1QBS6Ic2Ny
tuquzcvbgGpOs5VTW4CAwBlYhHbgWDc3rSlHBQZeRv5dsVyeSZAuDg2W6HUP4Z8F6BnRsh2XHlly
kTTCFh992800uSD79NnNGJmDxB+rPyj7inrDlIc3BY9LY6YTo8yphsNFev+9VQx/ESbdVzYzcOlN
D7DNyO2p0PXUBrSGZR+u3XDR8muiTyyAft5M4ag/EmKPv1wrW3He3k93bL4ZtmcYFE2W6wBNwE5l
hSmtD0kp8k0F3u9EyUbthtP6aLoRq3CZmkWzZ1qqsyuEc2Oi0dTSPRfVrYJ5pkfpW9UyFb9MigKn
gn5PBU2hC0uZ0ZD2GEy5GVxe3CgfnHt54i6Nzmc0CnuUw9KPlH5Q8WQ7zXWwr10bPfPAQEma5QB2
OWJPglo5mAfnd8JXh6va9Nyv/mBziDehABW7M6Ffxa+dEixH2UNdD0Kp4gqF24kKHUgZo3HpZEFv
9pqvFIi/jh3qgzbk3Ih1/mAXq67YrlCHvxgCZfyXF07JmIBbxdIGGjfJXR8cLyVufPbXIr4frZE/
OqbJNuoeHJxFYePtdpHdeeYR5oBH0HaXjok8R/MVa2vKlOvaHb9DfqTKeJPbDoJ5sGxShEUgdXkl
PGyny4EjtWOvaatmU7paeciyb/P8jwYUkOK5W5AzgjXppXJ21EytEF/sxKJxijHIjwH55+1qQCgb
47YmGyyFjd4M6ryZNSTN9J+uakSyJQ0vkG3owjJLlL1j62v4qYy5XA05ttob9I9tPg6KZb3GEzED
tSEfXdgGSM4BT+kJcrhTx8d28OuoRFIZv9MfSI73RseyEkrPWTA0t+XfvjoVnV3+X6isduF2QmLw
VFIYK5eF5jBVmo00dpRAHB0/u1jeSzISMoAx2zm55i3L33a1FPUu/RLQljZoAAkMjCQsotbWP77o
S3UTkIhPH3Mlx/bUvu7+a8Z9ysqzZ/sg4ER6NtkAx9D7E4ZjxKlqNZFxt+f8SxfmUrrg7FVed2lJ
9aoOwNEOoYamZ36tWfbcf2FjnntX6Okfe8efnOw42XqAxiemwr0puvCvH4rvEXwV617x/PB1P4p/
NTajy643gqTga42PI1q3kbGKPBZNde1YbVOUEqyX51qpoSY6FHZgBZ9tG76gJf+cVbD1OgtuLTNq
1MH4UODMF+c1b5OBQE8sfzcOHhjzGFZ/kMtJt0xiI2WvEEDAyrA5yE9JOKz2axqTaQBsA8hKjfqC
nOWeKL1az7rO4K54LbRvuhc+zGpnQ035yX++YBVJVV7MNZX5Olma1QveeSFxMOQEhMPgkYMPIklW
yKUgT5ziLN4FnAYkbMbLk/vAT0yd9iXfUBbpnPorlWxpGMQ63WTHlxHGSQu8BjRV8nIYASo6gjmc
RvApWHc8xqeRoTmVn5Re2KRaL6H25qzpxPAKaDRFifFKbwu/LWu8sYW1AdxCXDZ+SmKbYTwrDNQZ
GmYf1uOQAZ7M+8gKHUp7OpF7gKzmGhJ4ljU76c3/cccPIjk1kWBo2zZN9U/2HTJbz3MlqngomUXL
vzSqsE5eEER/eki/6xxCu83AZ9fLYGZfPQKyUdVDLMDrgHkLy+on2AaamOWHm1Ua7UXHY/pNMN0v
J6cm9miFdc1T50iq2Yg2GdKIRVPp6XjxMUNcLtNiesJ37zVWONJd7OmnEl/kc11wDriwtN7VSw4w
G3sB4X4GzLJ2S3RE3EXfCz+hEr774hNUAg6JipGiUVu//KMwF8BbjDsmnsi8FN10DJ1S/pqMw4iZ
QoRrpRRA1gQfjFU9zd+f9EbKnczpxkyaxZNIgSmp4RqFfBdQtwIcKYpJ9bHeppkGeYeLzYTe9TFu
2Gic3L3ScvZsqQSAxviHKTaZckbqU+vJ47mvAExwrTL8wcjLvBz0LVe1r2gKZ3jIQpn2RqwL1AUd
bunFZFceCGfKjt62jwqrPk37iFmQXu6qTtZRIXvTxUKDERJ2bQS7cDTZ5cDXHQzUcEkNpvl0w81F
W/jVU2uGTnHsb8n1tO12kTOuTZYXXI2EmPdmRGCFTuYgYd48j1MKQjtixB0Lq36qeha8Lfz+GRj2
H8tTmxN5nrO2GD0XwgTMWZHQnpVvSRZUqoX7C3zPTNDWbjaJucImm0ZiLNRUC6OimBBjaFmb3lrb
JpzXIW3v/731RCrwCW6AIFaFBx9fvH2tipQlt7DyOPrNdZoH67xk5G8jdLG5nM8Sb4x1VLq0JsP5
vBzYCSvRRh4lr3yb6uyZApV3g+xxd1Bcy1JX40GEcCJwATTeD8c93HhheY61Eu9xtWtBMsCKrck8
wViDF8MtfdihUtaBjndXtNK/81t0aP/EavxVZLhi2j3qIBa8lVOyyOrn2bEq5IqnkTpgJEuo7NDo
taGzS5XtLnUn192fTyiJg4I0kvG2dshRZqe3xya433oWuw6z20Me13UwKURM3Q9Y0Wex57/Ammi9
zeISDvcPwz4hTi+R5SCyWSG2Ar3G0PO2xGFAdhiNCKeVKn/nDcb5NQanohonG06ESMeEoi2xcj8L
e6g9LO/Sx5eB7IMSI/7hKdMpi+qG3ZMPHnsOG43kdVMNACTEOL8QAX7XsExrlfEnzqEX3yUQpzzP
FTMmS/7pnsZXHdL2hI/5WhzfBoJtfE7MuW3d0BgTELxfC4gBwR6HSNKMWRI+YJFWw8Dmftid1Vna
3VZhQUthBVdMZksEtrGAXMlpHFYwO/uX40rpz7LRqWhvU1hJPTtUxMKWmjLCTF3WKcZUpshTV68b
ViWorVdz5TXOhF2SvV2nDdJNs6k7/fpU3cFCFsVUFRXGditEhHLoh+bM/TdcULzXtWDALxXK9Dmg
acBWzRiAqo6Fm4CttO1CjoMoNSCpeGp/e0jcpf9rCJqxQFjRBZ21XWcU3EQTybhgOBOfB2ppkHik
UVEg3WGlx4ij4cnXzgqwLvBWVywxha2q+rJb6wx1zXtUYzngX9nTIt+euWn/nEnHeaMO6nOAkXan
5woVra407l6n/TIbV6p1n1VADaLfgyyuN99LdGJNacsal0cx6lPv8poNjaxN09ljtF0stSowG2CJ
hFqnF45KHBMp/edECq8avOaTgirJzGOfBtaje3rGI3h6IlMAa6AuEFzvVJIEwnRyoy9T6SgkYB+S
Z38Ajf8BRk2mg1K1aI1t26niqM9UT6i0Y02V9Mot2cJfhkfilCIfavUSLKMtgS8GoCZELVx8MvXa
vzHtJV9iXQ9dPg6K04YNn7IzlNBHUx4KfY84s0YVOYFtfub69AMEfDsgPyS14tcr0bnEYL8SHMYz
VTBZzeQlcfI0GiDufYEUSrFcaMKEorZDyJAu1QjikNEHrTMK2MJROy9H/y2aRKlPBjI4x4GzW3yb
zw6IxPK7Mb4IZantuFYOCuzLKwH5n8RYFWfDXE5iV8ViGHsmCn8OW/ng0BtuOUh5JdEIXoE2JAGP
4CcuXfYYUDYSP8L9AcqmzPl4fyOFVPbrmrnjryAhZu2DQCsiwbGlIhGcmhoGrraewoeWmC90AOhE
9G12WF3qRHPPSxWoQMgxujo4o1TYXkG8FOeTxIbTmINixobJtyYYH+MRxAvozICV+PBw458y68ua
yIIqkVvxWnlx9pn5+so0E/8s100VzMoHNGTzXJC7PG8Fmf9980/eAyivd9ZIeikhlG787wl2TelA
egsXMif4KsfaHoybh/bQp2OjyDZ9L7fAN+d59YqaOU/sew6xqJKNk/nza50E5Vxj2jfvi5LbdhsZ
OVb+ILiJBLXNOJYijSGIF/2qPdDY+TNYi65w3fRvXQN5MydDstboIJwOHHqaD0Yb8ZaazNjip9bS
elnGnijFL71Lbf+XxktDsFAyVDhazOY6Kj88n3O/w+210ZkLKjqaZJCWPGVl1QduMzTfdJUmi2tp
ZCUQzddIjP/M/izpnAcLEVLJoSesoKgXw4t3nkDIKFyP7nxA5/lSwLCz7h0SS6ZL5FVR6WPbcY5r
BVEQg/iMAKW1jl1WzQ9iuBSq9k5RCTVgxe4MF4SxPgm5yAQp2JUY5tjeO3wezAvIze9qBpYIG+y/
9xPDEdgN5qgVWhdR8uy5gy+ar4Pye/WcQkeZ8hYZgxbD8W6HQIW+3fVj8Nt3mrTfJlqiHNChRwUx
v1A6dYbyvbFqdRML1sAStcBUOwoFMlObDBI58mlii6rRGpMKPPb5b5ibgsC4SOcba0vk2iRN3xRX
LiKvAhjEt37qN/gzyxQwQh3lKHX7l6Q79sCDSW2AOZT8FFyxf6CH11lN7O0Ak5v/Zs4gGIPtvzfI
gTtv3npqdG4XzSph+7jYNUjhbxPuZ9M1NzMJP957MHPMlNu2+CiUtzT91xgz6WAvLMg5JaBUpVnW
elReX05FLJW0lVhyvrFSX5KsJhF7hwJlIkLd52l55mYLXbId4qaydpzv4VYz2475nsKuPNWgIYDy
dFVSDw+kIFAu28DSEgLKR1CaIqDnlafrGDRriRjq41qDeGCXgoaQ0LuiAKJTo4J0US+kfI8jHkzq
OAPRg8LeAW0Wq6r/Ivvm3bcq2hnPKmAB88Hvj9WR50BX6FoN80ef+fUrVAm/rH6XAIuRXM3sbZ/O
y9FDhvM8iDkh9mcB3RqqyXvgmIZOZ7HxBIpebCnhyDUpIbw0UjWw+Iigex+ZWxMpO4Fi5Mwhrm6d
X+kpTGQ+hnf9hgq/cqzrYLy3gZG4AA4QJpaXBTxKbPfx+YjUKY8plglbobOiywdGbhTsvuRl2D1g
ZDnduTWbolbBJCYHhSDgRRv4TLB6WJ6i+jYF7dK/YYTNV1ML7QimcjIoF65XHdWDt7vO6Mrm5nm9
OG7iqKaL1wLu8gSbWxLWvHfd+TCa8kam1KhVzPu5UavZtiULR6lK0cifG3bTQHMRS2IZ0CVlTqIu
NN8Cy6rQIenLY1C94kb3ASVvfk31lA/r0WZnDgE+7uZfw7gx7cRyMBX7zKd2Vf3rO6QcnljcReQj
iezUTSwh0VHgp7fYOz3UQQa00bIAWUneSOY3n9mJY3IZDRG52/nAHuajIRoci0TidiBDIWgIogaK
NRMZhqoBjQEYIEufWurwf7Jric3u12iqeSgCTe+4HzyyPiNDJyvYPf6aEabF95oEnVvomklDUgRw
CC1Ebcygo4jCOTelQpKY/DYQ2W9F0sGw2nivsGeG+GYnZbtull3ptK36xf3jfbrg/3+v4BvEb5eR
AnwIdfAj8qFoXvahqWphya9Qzx4FoIVngIco/Fi4U68jBhmTL9EhmbF3sjK9uYjTfhzj+cjbCefk
ASekoLUV2LTxoLEiyr+Lq+OidHL7IJq8akdlpt0xaZXhamQluQXFT7YrJEw7Ggqi6KinU61kWriz
za6O/+rEV0rLXXXRs8n5/jtCKmICebK8oLXeUVR7JR5Iy4tNKuJ3VFF4t9nvs0jHbo1Md/oFLcss
uTNY+nnFuO+b7Oe2kp5ZBXz+rn2WeSaSz7VRTYp+sTaGWYRa0ppu81vv0LhDpniCuu4V3f1/dhGE
538i3WgRL80hEcZpRZYDYtnEjehdOi7M8geRFOXq6tkConVe1wE45AyRUniz97TqgKxItqYt8jO7
2Pn45TMgXSPwZq4+8mo+LkJ0X0V8k1nXQA1tSwRx2/IC7MG0jrdF7Ba1Gfg7e9o6Rmsvm9Xvlpkj
R05sJsoqMEFqArIp/U26mTJSJPCIldh9CSifSQ+RAjeHKA9l4gDYY4ocJ4wTiIbNJdd3l9RBzPvU
Yv9Sr4+BK+FWCWrhys6r2gj9jK/jsa3P/nN7qz8uPuFmQcaVgntB4QRjC4uF3aPHOqLOCPVf5mg4
Zi+k6l7XMfZK0x1eIbpXNv4sxMHafdmOc380SmtIZoftzTjJYbbcSHWj7sLARocTAl9HsBwfgKVs
J2mlmfzeieBHMCtmQwjYbYPVgur0JFHS4IjgrXF0uGaOgcFJ4WFGXRy4FxezQmgF8EhmwETJIF8b
btb5j2mY83ygZ9b8dO/qfqSEUANAemjNNyHQc3E63cHJp3BYLb313A7nuLbiOXt4Nlik550K1rN2
9HKWb3UBTj+rzYnziE7L3URhhnLennBVN+hCeXz1+eEzsSw91ROqQ+M0n0j5U3C75wSsG4hoyNJw
9YbKbFvlhfVLw72n6qeTcrFxYB7Lr94o4svcy/Vh0AalDgM9YpLr+ldO23OGBlMsK2c4LsDYXJlI
EmhogIiy1F4GEMd+uLJanuapFI/PJu+ItqZ5C0RWx614NnlEvFHBSAQWtsx3Jjapne5yNDLUfKXX
uxK5F/qgnWf9vEy7IWHzIr0nB22Gcm0zfolUd5swZootFOzcOd6FJbwqF3RUvWb/ZC2onf+/4ogR
gaoTPm+cafaH+5koQsL0q5tNech61WPXcLRNRY0FoP+9QIjnOZK9bjF08wiZATIj6v33QuwNyYEb
Xt5NQnxftwDHZWWev80KOCWj61RBdwZZ12WVsB0P1HyyypNz5Yn4Izx3YKt3g7Iasb9F2l5oJWud
IdJR3x/ul25+wCB+cg45CnabxYsP3w5ur7Oh84TZ8q4m9Cjqwn2rZqGt4lYqlWmnB4ATgeOyc9xW
04Mg/QFRlM9pr0XfCBzKg0lUuhtPdsVxKp2O6+gp9C/5pd+gRXAgbjB0RKcf0j88AWHtett0+MOo
E9TYjERcYwf8HR831mUwxSUGPyU9/Xx2ceRaYk9M2nLJXwpEwYH/OEXbqdzQWlvgmNT5bnyiEbbh
J313YM1Pf//hJvVNdJocB60aWHzEI52F7Au2pGHKfE7BEKX3NNwXFq/q/dNX1/OSOCpfYR97kBPr
mKcr3WBk7kupIJ1ECuyLZqleY0Mp5az4EBQvCX6xoNmp/rFMGjZgZcrgvXjzA4TrhL48a4j8usJX
n6uOHDSAhfZY+yhcwahXYJB+k45pDHhQn7ccmkq9ibvaC2dLq700Bz/ImM52xw9ijg0+7vqIlgjn
7LPQn92IbAAJ55AP0yIu8TAznIouFXaMI8xn7nEUiSllUNrTlbgX2MWHz8o/1QEIiSunyb+Sw/RB
J4byIBe7EgAcX3wTb447d+PBrIHDNbeXu5Rr7LAvT0r9v9Bd9CYmVmCTbD9mAq+3IzIxmHSaNx4x
guMAakjEV4JmKLGE1AcQw2B3NqGabFRs+lbPEKgqrtUzj9PjQxjeCj3iFqnCoHuQbFe4KoDuwdWi
yMpX2nDRJxh8eHxARwfGyUThWGHDCiECtq5m4en+LgbOgm6XNJSDhNh7nv5bOWvHiFr+Lud4ESyc
1PHHV52lrNVC3pm0sTugWlOWSrledQmDp2g4Jjc2hytQ7HQPRC7Va/iRy5mLQm035bE9eT2eRMxM
ah7RAu4R5BQSSWgHITJLcsOQB0e/HwyixVmiL+LaXzHfN6WNeVBQF6sFjkpvw9jSCtyfVG2NPkUL
KxtxNdUZV71pPg7IQiZh2qqjfhwEyZ68uUpqn3+SsJ6hC0TP1dbcOwpmYHkyQ9sNTQsBrCkcg/VE
YSMX5X5rP6NlQ6SBVhOGwAJekv2R653HqCys+elEID06tSsQbv/vdmPLRNVSAup+YZuVkzLnQ11i
jhigg3ASHsX3wiRXEn2Xp4n5mhNuQEw5vC5LWGbMd2CT0yxnFMQ3g4tftizA/pjKsQh5PUOYg5xk
dgh48uhtviSqCWkPT0Oy7SAhvESH7O6cPLXc5CY90Cm3kAD7LSiU4ZkT2LUvDAkfj7YnX2624Tda
C/zESo+lrWZE2233WbKbOdHayxhh9IcQw0hkjE2ubzJrldtP3pGjXddG5ssEOFWafU0VV6Zqvm1t
ELwxJ0lzaMcNEWWATu8PlP5H7vUYP02xuJ1BqePLrZdCgYVNTKpQi3hdDG1buQOraOG4osn0P1rT
OErUoYBnS+d/FKnVccv4dAst46T7GlRl2cWADW8ljbAlaSyKBIraHuOwHM46ey0wrddos2trDS5g
Jf7TZxOR39J1xS5dgkT5U5Y3C+TnlPLrEpxXMrUguDg1ac4+VTDRQGevXK1dJPqpXpOtmwLtxX2m
NHoYWBNF0l4cCt1pOy3EwiJSql2+UKnWYkGwTi6aEPpmmkwcq5pnvCyPojO8JwzmNl6V5aQpctgP
HpSqb+9OceoxlswGNsWE/O+RoJku2+QH5Na7s7jsAHI1uW+ufq3jq35St5eWOMC8YI8LPGY5kynG
iO1g6kkfjo+aTYd8tQQCZSuW8Pj7jJ2RgNwK4OTgcI8DDEvvKYZDxWxCfKpau7oHWuOzMEsK0BWC
W40PAah133gQWGjxeaCwtNsipmnLYDEXaPd6AwpPqHv/ywR9zOIlE8hfqqOiiLKq55JSyfxty7Qb
6WGBqGc7C+PEf36F7W8jwTCRX6ok/tXk8e6LQ3nbtDCSF1dANyN7kIVJOYAJtKkGXW1WTP7o3S/8
cd1aVpbYEFgx9ggc/LpUFNLQeQE3M2IIsh9OTB6NLGektVG8bDAsCWx2hi4izmtYf2ItftPIRhgW
zC/ly+TrSNlqFH/lPQxCU15+L57Pezbq31q9HAKxI4Yc3bJF61q9FW5o3ASld9dJCaA6Nc4hMkEO
LACMfDaLGoSLX3UDL+v1+KiTWb1rc5S8iSUoy3kEu2UGBrrtne9MiFYT82i4a6Iv5I6miLYSVCnV
UwXwWBIY8QKGsr420cFkzcWsKlBUP8EXVzpX0R5EPeZzqov+e8U629xGx6w3FG3T+T1xeuZXBql4
RpWihp3Cw2SA0+kK7BnMi92h7m4F28y0WjXpnK+Qsdp3RQzb3fXlkRNsFXooC1xGkqkxB34+uCh8
GDIQmVIUfvj8zTsYfLoHiABbHkY0RTrm326F37Nfes/sRmwrnQGXVh048CeHtPvPN+iNj23IoLpf
fNPoCVFYvgW90ruwOAu15Wr8UMdDO5s+9zvwMdl/NfnBX+S29W+oMCU+KInk7P8X9KOmPTUw2ERT
5oCwFH9yxj8YWeInr7HcJGj6ji5ad442bLThEc3g03Eug9s881NnDU8mSk3enSBPauzCpca6x9D1
1LlR/wjCid2tuUtywtSXpHW1Qa7+P8g8SO9dhXuHYf3ew+7TEcNGIRHd5lysrXhrsB5ZDnypBAij
Puc8iNz+5+B2+MPCiqnkyJAFygvF3nmusfgf4mXKZAA/RAwGAkGPukCIA+oiN1p+3o9xvWIvFKjx
VSPfG/7ltQImkU64q4uawxwoY7Ena/AkpdS2QaujbTFZeNVdrtzz8nVB6Pg+AUItVAcb+Rnq/jEo
OLLpzc7edsZg85MZQRwMF6tXdleTzh0fAxJg/6mNkL9R5gW1ulPfdQV5rIszwWcJPuf6g8MG00hx
/8kcrTyb3uy/2u0GA2fnvHB8WWpDxXRxC4DgoON6TQDrcndj4JoqobEcxiLitcqsoXEpAdSgq1KL
lXMwm/ESflYM5S2LeTzQCk4MNw7IqTZSBymvoVKHmyEGV7plyvaQ0/KmgokMq1IrP0ZQCRkUDMlx
oSmkxX4HCOrXknsNKmxSr3i5emQ+2JIgoZgNJC4JT1XAheZpijcwLG9R08fuwQGaQOhdMz2sTyVm
GvaHrVzwDMk7hHEvH6xVuhDvSeqsvPQ8urxXUmMtEsm943ddpUUrwjC4XT/35NMitSZmwCrmIw9u
JzHQwdW594fjV5rdkoC/zi08oi6i+BgK4XKOJwBvrUGYc/lFUqJaUJq0ruIYYEPJJn511krW2/2d
C86GteRvYt+u0sScLeqI9DMBBNsaI/wz4n8TZvM+urFzzC0U7WXNeRJRPmsGexx7xEk0ISkYEj3d
G1bDLUy+D/dfTW/zWe+KPxcE9uB8jluSXdJ8lBX4MciKKzjbTbpRBiONsleIUpFhQw2bzHdoIMlh
JOiM8J+JUPzBr2CQTdE5wBIBvVIrchcR5tPZAvrlnJPyMzLBPgqhnrPxwx4hh94morXjrSEMLtpo
fNreKFyFu404Ud/3vxOSXZiRcXDLAyOBabkl2atyBdfU5ysdW0boNN9LMV3d9Y9dM6ylLGWst4eK
58C0Hkv5Foo48EfqaRXN7mfpXsZlHPbWtplw1RVDSsjhMZqYixBzxR/9yOn8L7VEH8u28CUaq6vY
Wjg7gelvSbp4a7fT29sbx4eCdG7NZTn6HgP1A/YJT72N83ZCqd3B+KB5XPbQJYBO3Qu3unAL9SkZ
S+kvKC8SdBbvI5dibKwZZ8LN/oESWvVh8SK9me1p9p9OjcfHDmcD72RqVpoBwMcSHFG5aH5zH0eS
1Gk3K6qkX/2EdX2ByTn3nALcHlGlq0/jDv0z7QQJeTw798wCBl9YEaWswKyksZtcC1IE4hYlUfYI
9jvJFHQWmzOq6Oej8GVrvv81YiIGrYGCY6O9STCOJ8MH2cHMZxemjhN9hBt/WDj6bWRZzeXnZ++k
e+hX3Y6nQrtnzUondkPhhp3NB/f79X+her3d/0a+kCt0RCtpDTWUZaqScU50+ubSttXLkwjrBTrt
IZg3K3pzxpe8aZOQjrJOz5ws7o8p1dHymp2B0XMCCJsuUi0nMVj3e0I5QBos2kGlKRSEVWI1LD08
AFFaBJ72iGbt0rmXPgeIuairg46WcfXiQ4zRYrNlsG6xqSyDSlmERbaZe//s/Xr7azAxsnnOxkCL
7yvCPiLK0x4mq6ZXApNzes1uoSQMkpA4x/OJ7JQMvqqhxyH0No1pOEl2Tx6VmoOrOIko65LOCWH4
bFlU3y/KCwp7nvizvSmcPkXDaYHjSDKox+c/nulzCu/oUgRX2Pe80ynynJxo0UAkhWxr929BQwFb
6om0M9G3emgfvPpQJUMM4BC7I+W/x+PW1P9HtmHpcUhnaEM28U9jpjT75AxH1GuluexhIGmEVXRZ
m8qdW9mXDv9NBsn0cFy36HI8HNc7X1BPKjgfNrGKdMrT6yFAUIyqwIy3Ocwezg9TZ3Ksmwx5A9WE
7GgBXy+3mAlr9TVHMv1eYwvP2cyopu1orrVAtC0/F/xrFyaq9sEhbXrd6WQvcPLeDnEDA9YCww+S
mwfMlCHNxzIxI889PZeO1NxA4B1Acccg+CNIPTqyFYdYBWxLUuWrBr8zybC3m6nV71spnty1W57G
2z/j7+6yoE8WCZ2IlyKU0YRxG33wdmzAU/Y3MEEN50/Tsd4vuK8IDAjxT+kgCefHaI/u5L5N34id
wGQsbrjI1PIHcp6imf6d1w0Jor3CGpRXCW/PC0Lxnul1HKn13lUdKQYpHd2heGOgZbHlB53GzkSK
NI6LmQHWNcts2a5IqcGy2GrF1c9xeXCK8x4XmHUiwwVC1Bt0XhRMsta/X/z1eUwha10556y6bhmD
3f6HdOS3w4q3q9yHkdmlsqfhh56pKuIZILV3A/KCEfU9FAdltIV+gHRNdT76y4tREmQL9O39qEwQ
C3dSjTgfeURA2jcsvhJm9BSgnJxmleYGgTsd2xUOVfyYNBwjCeUtlVptSEtNB26MobjPAjObJzf6
5FocLbSWYHSy4DQeDfZ4hB0VFfFXlEqCU11So5/47omxgJbh2bG1wFteMNmHcucGLCK2kFjJyHhF
+1YafHj5EWe/VssjvjKaCwYINdwRF9WWMDk5W5RNNedtqRsBXpxTUF8AtBOFvitIrK71VVqkH6KE
kGeZzHAEgnE8BFzJv1gqi/WM9RDAsikapusUJZQoTUA3o4iSy1OlM1EuKd7r5Do45GbBs2sQ8Thh
qhFPsk4RaDcrobLiS8mCmfA2s5fKx8m14cA1LTf1FUlet6aVxxdtS1kzy//U4uq/JSaci64nHAb2
U2jfMmZoe2Pxk64eakehk0AI62g8ZD5A9bFQOcJFF6GJ+66vA4N4qn65vM2S5PY59Qr8jf2A6EHI
NfTQI3YnOBTMTUd7HJjFjMFH3MiFp4uU3bIk6VCVBfxlmju96B3Vsrwjo/mbXz7gzrFo4IRnoCM/
yCMnRtzILCH/1SO9EDtuhaeDclPPy44GIpdjsIVteAYhv4/JKcr9TrjFjZvYU2CQjH14Y7XV7THs
4Ko4zfrEvDEEFsAkYzsrJw0EVl3GiboMPRjLw/dH/+EFrpBvUOALEIebl8/wkFX0D1gS3cAawctQ
tszH6onSzZedR7gIBv4Y14n/cTx2V4RaOmxFn3t1i2n2436UWdLP0t4hCDNkNs2yyq4F5/tiC9XD
SO00j+LQATfM2plNivnUotQwpMgac0faDP1B1bZ6i8s9Douyc0TWnkAxfDOn7c2v6s0dHJxRDWEK
HZHoznDLpKdGEzHk68o9rXyPciiTDnDqTzXTeJ9YMpnx/DZMKRnqhrBOgd0Jv2ZjAybADtwre5u3
yW2VmcXHMo9EDnwNLCEBp0/nqE29HookpvE8IqLJlu28H2QarsIOlDzgGtQKzMrtdHA0eV8Qh7D4
fChTZSZ9VaiVU3+be0Yja2kB9gD3x4zDiGdTeGYSM45jPndOjsdcvtJGZAO9DdHSSRrF9GVEDet4
ZZVCHq2oZiMMfqlWpEi/8ZMFNQ8/LSKWkHAUph5zyjhtMI+9DqPRQXgzjnILk9AtxuiA3l0f8muR
WW5uVxp9nQST4uJVQfwQBag1F4ioNrLqntOAMgcZM4v9YcPDQvisei5SxuVUzjwg1GHLFEPQPYzl
pCTVArd0OjNtn9aBqzBtqhlcnRadI7g7eZoEtJyVjintbWbRzfQuZA1sLp+Rw18Eg7AjjXADuO9W
agYs7lBV+SsVXWlnkhJaIiEKO5vLu5QVKrBTMirHhcYhfLkByj6ynlGufyvFZ0YMLnmia9agWRJ4
IW/TUlAGx6th5Snk3+RRx/eRxUFbQqB/TyOuJ8w+qMo+be57a9tu175CCy5H4fcgJdSOwddUKx0P
zaO3yXfs+36IZD3ubGAiVfcwccPpjG0acOj0YTH7dA8P5gxX1NizeP1K6JGYoMj0fa+Dm6rYh5FX
de7ld1FA3JpSEYarBmSd8TtvnV/qy5LIr4GkZCM894+Y/QRhicfbxl4WbRwUSMio5uEU3avzZpE9
P2+siKbha8JFt+opl/WD65oM5ZZdAfFVGYtTUc3ZFgGjGvd8KjBG3q5VCmLIrEjX5lMzwpe6NSzC
MGuCylH/RcYhbm5D5AUm0uxE154F72IICWYcN3npCK47qoBafK0zyVkHsRmTKkM7R+2mFn0Qj3eF
2/3V6cqm4evkZLBRFSVhpOc77sNOCcVGC2clqygLzGaF/wyXOn7j2y8eRWjFLIhxfg/KcYpk+tkk
XypRXD62+a+IywNx5WF86cY4M2q7nuODfagisGuEhcFaThRiy1wxtNSOwd2nJv61M/1UTKXPhfEv
PU+FTsQnUZCvscHq67rTlj6vznGcUPTjXwOYkE3tdG9W30OychiTG4plXR+1v/J0zObEo6HJ9xin
2m8+iaw7TDrA8y5EFuaCI6ZuXPFn4mzu8Yr751e3DJHaGypao7CU4c0kMpDpyDG7fIXsp88X9lWc
vRhN+zh9EuaigjguXWHCz33itnfA5c9CLdi7y5G0CLArgyAPx8iKggbYt1NqHMzZYWtEUs68/Lr7
Ct8G6B/B0ZDmlK4E0D7d1LjczGMWLVUG75iNkQYJ2YZ9a6vQKkE5yVs8Xby+a6peHFw/Zaf4SOFo
c6Ep9RCxI1eH7MjEXTdXGgNH0jeEl2YAmKzW8PlpdYLXhBWx2DWehiiHKaim8SVWEZwZR/Ta/+yO
0EzfHA+4oDm13eFIUPcrwCCYA521eKTvu535HPYvWsB++En7jiSUd99+2y+a4gHMNWUVhyVTmotE
pQTJZAo4SgL00FASjMZxMGELK9ZksVbrtlviTvdGpLr/kP/6hN9EvQLXJdpPGl3kEg/4n1H7xF5G
w0nbw8vbcEz9NDxbRlKcsOvvOc7FMJdnibqwRQnCzHd8Y652St0CugbOYgVsOw78iJAFxh71XA8O
GHqBqaFYiLS8+xyxjNQKLfZchzyJO9cDvbZ4A9/qLQsFpwFt2gxRYIEstQHJzZPE6ggqdtIwIS8X
c1m4kwSuP96JWPdxYdawdiKnNFewI3KLQKUHLUxDRLPAgvnCuczkKAcWPgO42S7aBXyCxXeTE/nP
gmsqDV/lK5dU9H9QwBMiZud9sF5KEXxFMBoPe/aUEjR/+zXewwgiDzlWAnZVquIRJjR07a5XUmS2
MQai0gc55jvzyX1dRvadcpi4IWuSlFSx3ZdIjTada22zl4suTaDS3SVcOQiFj/Bz0z/qW+DusB3h
42z3Yc2Laf1Y8brtHqKZHzbQR9vKyUvtHk/0uUj6R4x/4CkVuGDUuJ5ozbXD4yJMmduvf79w8+R9
6ULY/naxAF+dep71yGFBCfwF+J/9z+75t3EmOstmVixKx4mNURefa6tR4C4lnqXx8SvXnLuLE8hm
VJ1vcJU9yn5kFWJXl2ipS/SweSVkqLnNexGhocb3SDY2vxdH5n48TZ5kdF5GVIYBDJlDQrA++Xrs
DmJyg3DQQFuRAXOX4OmsLQDKpRxP6EDRylk4iFqFf5XLdFFm8M/ewwrWXMSkdNKWn+87xEZLB3Ou
dj7jUA6hmm05nB15VJhzGEX437zT25XWe4ArRtzeDF9k15f36zKtVVFJYvnLTGlhFWK8tbvNgXjH
UkJe45pmCq8tTdDl0Nxy5tHDOH5+exLLPB5idvblgVlL6MuyHZFQeFGF2dQre2HzYJfurd1eIOA5
svytzUb7cLP22XByHwwjBcnIzQdN/SRopB7/Tlrwv7jIGEnOkfLDXj/V9CeewgQIUaiH72GdisAU
Zq3DuAByz2cEoFvL+BmDsktaVDfwu30LaaE0YX6doAUkf0zKSNtV/lJ+cA7cLJnrRBOcMsMwA6+X
3naVdPca1K10lzqrTi2Yv+GK0+QCw+iTvNzCC2rtjQD4Uvr2QsnXpLxVVLpZgWuYWa9S9lSOwCd6
tW1k6K1z4GaZYbOmeJ6yUzbNymIlNqzx/xknmXFcrwvqKhFbQpduD3Ws4ZroA37HyhkRI1GBTdUC
XUoX5Rw46VPwBdNIob9YBgQ3fSwnscs9bIJsQpwgtYWpI4d94zIrdw0rle+Lsdf9XHcqlH0BLZDt
8i5Lw9FJtLxJ7efbnP8JPTrxUkMsPVYkfMetu47N7msC/AK2JCSt7Bp9paTJaODnKdgeMaPieywF
QoYFVpMJyGdlVIVrQbQjgJFBrM5NOki0ngsszWduuEwnu0Fd10u8YBwskaf+QF4GpZeochaJM5Mb
5jliDRbysIWOGHBCwFz1cyWI3saonkPIWaAtx961dgT2MhptXA0J5P8TGErNSCpCEHfyZJdGLfuj
MH37DHwiT6nym8f5RD9Pv9j2c+r65d65s8FzU6lfmZHWzIEZrrvXh4tARE69w2ojoaBkWlyl1l3u
jdFMo0OAXzcJPnn7U9y8dhACbvnll8HMtpQe7WbktgcJzJZEBXIy+sPeCStdeB9ss6uiyXSVO3Me
dCHk4X9WdFVQ5bCxZwNN+/x4YPecflGPesC2TqSyEnsn1tvVrRl1he/irjZkqENbZWCnrk6U7YyF
EKklgdCxQ/eIZ1w8rzXAGd26un+guxyExp2S57VCyfG3BfDo9IWFpXrdFEOZmticiurOKPg5CPAJ
K9OvhAQ5pn4CtLGTlatem884Ugj7x7JJdCGssmRzXXh3LfTfbgKR0aXY+c2RPCp1UiA8QExWFI73
NMWqfEUf6N/nZHqtOnpuAwF5uZmdBKGjS6YY62OAY1MhjYySdfz+aB9ZdaAe+PF6qfxxg/Hc5dPZ
asKH4pst6btRHcyjuSo/vNRAFRxefQ8WyfxktMWW9ttiANIBOh+4RQFC3qZmFTtivpWQ6eQH/lX+
L9wFs6U4KO6qMTsLP9i4IbiDPRnL5Kop5byitlNNnvFvL5cWSQd0xOmQ8PI6O+JBp2Yeb/KY+G33
0fWhI1RxXEeMLepkosm+gAqzj6bLZ1GmfVRwl6uawRxRgk5W9vTMYAc0d8TyZn1DGFGEW+7lP5F9
tbsVN7+dPwYoC4xTBTZXkiJcN+2165uTIl55tXwONAU6Ss+Vr+ZzoIDrI2F8AJbAV5xrBJjvP28e
5PVTxYLQ7f5GIdAYP8W2g+N1pxt7PlPNNnW4LvcfLXYyCyUqevy+s9OM84EM0LdeshAmk20Ihcc2
GxpM/Xtdm+jRay32kOC+dnXOmGfpWkNkcnZo7xFqmQPeBblW2v0ksimDsrp5IWDp7wZ58CM451Ok
SEe7cyyTYcpZrD+vDFIpsbeUnKVPHk8uMkswS7NjF3UOvuxrZS/qySlZQl7wDjmNMTZ4L4JVQ4u+
h+XkOcowSxWqcYD2w+A53zUXizyN+ZQ5xO4SvMvBpXnNCTTdgW47qt+DS9+sTunBoX0Lt1sUFx71
HGDUoazv7u6vicfC5n3F45SwHoK1/eKr2HdetBwS5Kvuk420dbuAYwIyaloGHjxkgPycjhx7QvGR
1iEaoONuTYm4dgrA0ZOOTLIGAAkPIFmcvpwpcT5ytsoKjW/9X/PKX+UlsZeXSwogPNYacrDGR6Bn
wdApw7/C7swCPHutxZrrP+WkW3OMx5dRL14kh3Eu4jdhGhmwnGi6qA+T+guBMybqsF+z/4GNJIJD
907Jg7J/WvoPNOieRNuktS/idStEOzD9bQ/osI9cTJHX23rxAAf/+o8WSLujQnHnpLhORpf3SCd8
lFCs2hDoDiYr3JovUGP76NQouMld5lqJp7D0W75tiOBah1KTE+4F42F9YQbw1AdKUWAQkH+CwZr5
Gf/L0FvXiCJ9puTBGUx8CrLek+oMW9tmjJXuGCPACp0NyLfRIxydM/I0w/6fULaQoKf2BPEcKAsZ
Y2f+IZCkbcMOag8MP1Q0pskDxfrg1l6zGgi3KXlNuC+o11knKH4KkWSf5cUAYdNnEFXU8X+kJLNJ
5CK3iQA/F3q3Z2E71wEzGqKbB7jIUHc0wCNfWSeNUi6g0T7k46PBrwogMcaC42qgdFlCGXZu75ov
G0LuPENTNZQPkrg+yMYgfmzBtf5/OwVKN8Hg2p9x+Efp1Oa0n/LSXrWFrM8S7nBrvUnLgueFXcXd
HWo2+Qgcmct1OifrvkciUCUi/kmLTDT9Csr5bEmymtabprqtVYJrf4W29Shj62D6aetpp2jur9OM
MhWYchLZvM5NIiwh7kFayjuIq8asFwqu4mkVGcmklx7GlKqAp2oj3fN1+p2/Ja4Mspp9+KChE5OD
ZroV82Xl5+M8cv9sOeCW9uQgbDadD29SVdOXvBSwaMSdTxFuBk69ijBf8+5cLMYVDwjlgU33t1JS
WpnTUnMTw+OW8PNuMFHufWDf1KlCl8kNgXEvIN5nXp6Knt1FcD/awUYOqHMYiUNFTC1LFTWZnp0A
LaHE1np8LPKtSGApo6FHnd7xRucF73bW3Vl//BK43TCg1WJphAw2tLoe6EyPYPMXgCgN7s0sazHw
ySuj1noN26Lv7C721JDfYYTDh72856RSeHrZxJrDJUuVdSeKmi6xFenNSV+v+Nhj6hgW+gzuHkWW
PQe2qHTyZftitAxhNgGXyHVvZpwFhNe+pAMTLGqeYxQCOY7TePSWpwxEzHNfuqpt8ChRlqXwMco2
XIiazVb1RzBU3uXLGXj0AHn3XCyNWlg1cNEEkbTSCMdcQBqOtWF4KsHdN1pcebp2Di5Y20LroNSj
WBIMPy/cEF0K7kV0jZyUc6SDst0QJO82tJ+e95X5YXuwUolMyf3qkhCj03w3IWYoVuiClJNuoywr
i+7gCHzE6sE9JxJ2vcLN46ACc3jLhwun221B+J/H2TWaP0mNGo6e1y1ZtNZGbPUfOynCi99JdDPH
wacxsNc+DRZSeLFA0yiqgQ3ZWpx5F/4w+Ws7/nsnEB+CxiH2F5o+fgO2EKXhbQLUq1xit005BAhf
rLnFCJKdVwcTDwsg3VLvFz3+fR4De0Kti960Xg1Lz6hdwEC9xGEnBmXV9uqQp5Si1ZEov09udOWm
ByiIIUWe4nhdQDLmxMuzZ3GHrClpkgrufoAhD686VA9XLlPFIV+sQCYJgd5b6j+NvYDWLM3Ncpw1
8vZycuhMDOIscGC/79Y97MDmJF3fFLSXSvjWAXXDaCGmZgUeMDHnvDp+ViF2Iccqug1jqg9dunmQ
08DHJ83pv7BOiE4mwC0r7ahm2jY5TQx46eal6q94QsXyW+0iN8ZvxCLfz3XZX+Y25AHFublpIeEE
h4BbfSYrbF6Bl6tbVC6IUNnf3FlQkz3sMwp1IOm+6QAh8TymIivJ1y7VUkdrSk42S1sS64wD3IdL
wFp4jC6Ivdr7s9WWB1WhAM9DLvl0PIZsdLR1qEDiL0PVv4iJ6IGI1M5HjUAPe2DxSheqETViVYr8
uI1iDOLOsBcA91UQa9YoEyEioNJOVzEnXduFrM92QeCg1NMLsRkYdNFfrgHUtg8/k7Tzlm/3xNaN
2X5j9OMrEFny4RyAx489rUd3Uedk5QwhASgEZ7nRQhRtjt8EN7Tw+tyZ8cCPqHjfUkXlMWvXNGSb
6+jRLXaUzBe82FlEEozxfjeUHFrdxriquYtP/57dRLlxRobIQbKCeHTbZMaousWffCBfoUUL/0XG
baf4+3nHxDiWLrzrOlO7aP11SkeynCfxAdmAxj9H1AWU7mxNQ3Fu8agwyQH+HaLda/9SimXlWMpi
HyxizE1xsqa1gRNg5pXxBSE3Ktup58q08zttXZv9/zO1C3dY7O2NJrEiEL7cOXaX6J1FWPeNRsPs
JEjR2TdyAoRDqJhKvv/Ovgxn5uvkgkXRKPhayU2/eeFK8+p83S4BFz/t8YRiL/h0kcXhiGNWegoW
HnSmvsDuLDWWH59QT5S+mqcToOIfCzHfHNiG9CKaJEoDb809yHVWFznXABnUXztjBeuKDq6eryRs
r2dMhKfL6BLRkTGvqoB8TqU/7BH+JFsapm95YaSp99YzNUeskW80oM3IkfrEq7vwkYsBP0wJw5Uj
+tzSfX9hM2q3erO80y3Pk+HcaLlAmE2J07olKael1b7Q6c8IkdoRwnG0IqpQ+oX1llpyJi8jTbLm
MygkNAFbpWZC4YrQqk7N31DhKm3TQ7PTGgnSxytmgRICuoyxXxpyrtOAIXdEB3GDwEPVSajVX/Le
BK3sNJdhXrt4H6xAbCt8y2VpouYv4CigBFxEjeTInrPUa8a3GJ9UROiWjmtrfkqt10XbcuFe16bs
1kMlyTD4B1arl+xnKA2Iq0Jlx5fYSXUTfqTlRHxpA7hGwhiTF2AX6cDbxQyyxMIF9X6ipGLDHs9d
D6EFtxnmEhXBzDdLqxi8168NCj6GEqFNK/I8ClW+SWJCUiSrkvvrgpQywiUCEoYh/VGLj9/Yd5bc
6CJjyVQWFduYt80BoQD1Hi9ou4bMVcNbNV63izAcFa9aR9J54sT+4B01UQMcWG9Gg2EgyfQsRshU
FPN3KHfSdnV31tDZYTRnX/wOWtFqcRTC6Hvx2XfrQ0GPk0axm0byLWrMeJgglBsZIwZrnPQhknLB
n8iK21Zw9tiNlmlUHUXUNeDqLU6IsH6RvMLcp/uKTo9i41JdUmgKmtKeh5oy3mhaVHTP4XlL/GYz
QH3gDOTAAkccblreJRnOihvCW6Z2bXyMan+nZFDU0aCsKHSiTYx5aJnbPDsHvATYQMqEAbAKnSRq
9Mr2gzNVFxNk0u48HHxWsraIuIu6L0JN296y8+50nG0gIe+elbcjEVPSZhGKcHKTMGbuKUD9r5eG
BhWX0URcHLST8f1v1/QQo5xBiJ8gcmCnfkWhqyQVqgGhHKv9xhotn5Zk01/LiDU5XgOotgB0Olwo
Tx9S+KkQoLKZbzHe8l5Hs5P5ikvDbQyP/uuvheupxIMiSFtkVmLTPzW7D7AHlSn3D6EvqADZwFBb
tj0anSDaYl4qZUh+G8Y8/q2wzB2xv0O3zrC5jwUPA+/SE7qZbUi50SYltJ2hnTfKcd9fSFzs1EkS
KQUTO8Uc6+zp4WOUTphOb1a7buBojXfcxrzDIwXaY+m2a0u6EBfJQpXj52DpUwVmedLx+pMC9jCN
tRvwDrmqSz9rCJJvNaC083mmKTW0giAHFMIc9JjEBz/jXNgpRBZ9fUP6KNJU0p5/9wqRWnlwCGHT
2DK29b4ENtaztSrBKqF+nbG4fsdNYmsoZglii+NrERY2JOs5jkXfIAePdTCe79j5SG11CiJAA13+
mBdt/8TkMWhv2hpvxGdLBxbDi/yvmKoIIulMqjnRvWmg7Khsacfygae3JbXbT9lDOQn/lPCW8/6l
snk+ZlULyV9RghP54arvl4dX/VLNX8F8PEvYLw9UNzVHKSSZMLPpr5dXknXMA3csRxr6F/FB91Uk
8vhAdGtx6yse4+TBGB6gQ8JVMhYrWKLtnVWmyK2sXYDt0HyMFqPYVdC3VROCM6CVx9Rzhfrg2ci6
mCSpkgvzJhZA7TJDxQirzkzdn6MRLuIh6jPUm90EwQGpLZBHo/5lZ0x9mzMb6xlHZOKPC8Z7S/Dc
8gpXd/o/Xyc1WzKKEI2H7MFWAOJopcjoP4/ZZHo7gw66cztARRjZBAsMKzigtIwNRzEZEnX+52pC
B6SJLaLq7yAGF92pA3+iPuFQ4Rmrj7f1tR+V6s7pCT0GvpNYq5EZNHpKHL5mBarz9ssnm1qLwX3z
+Tq/eyQ77CRnyR7d2gipLkQj9UB/Q0SqnkMO4OLuJf67RCFDKFYsNW//3t2MaSXVSvIaW6L49FcN
NhMCZqV60gJVF/EHv4ldiSM/+QhElA2k49/QeaDkorkjQahETRM+aqJnzPLuid1PLZ1TwLBLyjBd
tPlmEzCOiyfi4jgO2EKkdhcFYoDiE0R7cSk4jY/VkpAqcsqtKo9NDoeSb7ZB3EQzwkYq7d6xrE5T
GvLRmuKucdnY+tCsatNckKYRWdoqGHl+1k5gNzT6Y8famlSMvrn19Q9EzNle2GicAwnP5MFIpMgc
alH8/qF5+lsfSfEAWlVF8K2ET6EmUlRgXZ9aYQVCo2YMnl2V1dSl4Mz0Tbswld5trXyrSyKTpd7g
rjBpyBbmLK7/ONZUnZ64eoz6tyhWc6qq1I0E0eF8k7XvRzClJlHfusdODisqXAGDu0T91eMOoZgY
mmXarjvLH16qr/5i7lZnTCLUsxtgxrj4PJhzvQmyhZ4mU1CRlDcmo5IXXgQROq0xwYFbRbEBGKAi
MX1xO1X5MIZ+bwEo1LU1nWHRppcYeaihNeH8XgSAPcjWPMdqhQN1yPdr/kia3L7IlnY6VxkBNmkN
Bc9aIsfN1fa0S0RFOr5mtg+T1by2tPNQb4us2VDNrsLUFCC3HCSfHDkSSwbFvtRt8nsRG78GERn7
TfFhAFXApGS+2VzO+Inpa+higCGaURlyjtoliK+7P5a8w/OTIAVd3mYy78zRg6Ry9dLG4eEZG09g
Rj0awbPO40+r2dgNj8KH2jeZm9E++1tzNLjVtmQT4Gs0BF05qjFHHODNfBwaSS4i/EqvPbzrPvtD
7uYXWVYHUJY6hLRu74OzswUbRYizZ7jEJdACztBgbEO3RgOdi1NPJITiovcSu/zSQTogv5YlwyTC
1DHL+9HRnToy5w5zrk/Z13XxlmQtw8quefNGx8+xdPqcMVIOjPPh8Q2ANU9TemiPvKc5YrwZkL8W
Q8yrY/kRcQtMaQ3m0xqmaEKdL6D4c2Yl7L/36+jTJOg/Zb7b4jJd2/rvlgx7vlMTKWNkeZ5iIh3R
YQ4TUjsWQtpUN2yu/bMWLujIELcp7MKDHzeKT4DJcYXu2mqMuqrcM/qvaR4/cPiQcKd7zx0SSAGw
PQ45QOh3ej2iHIHzk944q6vwEYX3Umr9BcoAgoH4PHDj5pV1buZ9hpBoGE+iQvSNBTED2UMsVIQB
a2qqLfebcetb5Rx+YU+4l+EAwFYFFNKirtAGhWw2jv9P8dn272LfEVasIEJmmvht13OJ4zwe8Rnw
SG3bsRXVzJ33gZP/1nR3fwgBJpBW/LziZu1AF7bCpPIISGX+KBvcwZoantVCM1yG0Uk/sU5AdFMW
YzoBIKyH7FDu/txTUwUcn0ta10X6ImFBQwLcJdIsiu/kY4Mbtpdp0KjEZ/S1zYh2KEXh06Yg6es7
1ywV81ZmmqngaG6LFcv0zFL5wmnToWMOeAUdaQqXJg4QbzFgV64hN39pV6k3derCduDl5FUwMHXx
OTDCW9pv3fsWNCQM/LSbQ1myfmS5m9S/7b9p/Q9suHOs0jGPm/1yaXJDsr/9rVkOz30dPhf9k1RA
E1NuanwTi3pN7gC7JTpywMFNp5/Cy4rCjVlDYmiiZBWgFwGXgQ/DH+i8ry5mpo0+Q+LDDH91vkCm
Zsjyi7FRJ756+VJVZIJy3QvigRl3Bgw1xpjPr3FVgtpFUQiwpdBmqWUbSX98VWlcaW/k7wWX40+j
vUW2nTdmQkfiM5H9Wb0DF4ujy7QUUnUv6EApLsq7SKO8j+A/tNs/4k2Bnt2Z1fDfwyvbyW5GJurd
YP+fLL7gQxtMc43onTUB7nTYDcNobco/58D78dC9bGpuvN0JF635Sem2OTAWM72o8J6v4Vl7RMGN
aitE2aODaHeXikv/W+/qi5nm5e4vRsA3j+QNXoOOySDDr4KEDD8NKUoYpP7/pu7nujY8nBwcAOkJ
X3IkzSgvvkd3pQW/FxxUoZ+hQaigk1B3qlJ+FRnmRelPifoNG+deJWXA88S2Lfj8srIl5H5C3648
MczZNsHpZNZMirOq/qo2B26v/pjwO984/yYumIiJbB/2Um+fFfpwlTWbdKtDLO182q47/3Lay943
vXcn/WGRIA1jymbIVhLzZWMPbRMrJdUWdqvTXOM2tBFORA6/mG3GcoHJmb1I/PC1h+iAvdvd30Nr
hr1ccTGr8ElWofho8ZNhK4ebM1nOV0hcFKeWmu/2az3MMBt1v7EVt6XOU7gPw/5Dkv0xrUWN3fdS
rbBWX+EzxNrNPrwwoP50mFmSVfUWLv045KOmaT57YnhOJ7tfDBQq10clp+DSQN77H9XgXgB4D5g3
1LoHzXVgA4Tdfx1zPhClZaihuLYtWwuyCIrYHlbzM8Qu5jDjGOtfJcpti+RuefkSwQKhM6EWkfnS
92lb8PBH4t/1gOkNiQg/5+t592WdzU1FVq+TltAyzt8A/VnTxPSiODLxeXVdKmA5G8hlorC/xtFO
tLF5MnkBfBktQ4yyhtWegosYSbk4JmRfzxqgD6G6vkzMcpqJghR5inP/B5KpqVf8wvKAICR/K4DB
5A1kAQDmHCGVYXBzee2Gx1CmyXs5LcL6IlCqo8eZOGJBdYoDjkULG0Uad21xMP2GDX7Wt6fZIGSJ
KVoA6s1FrF7fjPssuoc3VmNHdPiBYJdfCBZq1u6r96R1W4e901I7l5kFC4oN9KPvPcz5XlMhkj49
tqCLB3VKziEp6rKLGqVNNpDsUYI7QfyBbDMD7T8119qKY5n/8B3sVVqVDLt+3TZkuSFjdt4VFnWp
9tb/323RQKJ0U6oSHAxLwPxkY3AizEdEqgdXsSewq1Q+Zmsjn6LHXQ9wXCiWP0FotFmvEOZbDCWp
SBl4FqexPGKu2yprHfw2reUTQfAuNEQOWztj14blf5sa4BCKisTEDcXy+mcV+kWxLt/Q6SM4cB0G
rb7iLigGG6ZXgTGzgeMmgfimWRnuZKyadfMr3X+iSw6UuKFxpbU5tQ352BOVihgiDJH8bDO4WI4l
55UywQGTLWLqyHVS9J6oe7KynymeuO5+gVs492g4FNXMngWk/EKVPqBjrhkWWtSCOPhyusd0Xroz
rozNIuH/Zco/EaCZUqqXOU4BbJUwjHXPVWXxDDOnic4rjCvhfJjl7SP1bGSLGBhHW+SOQcHxHOjw
MPwT8XXuf3umpuXk5A77BpSPn/TtUDMIOJnW6ZB1lOyzNnCKOo0myPseRHcWjDD9TPUQ8tqKvLMg
XhEKUMUnc8dl+kFcv6jf+af4wl6vSqzjmKeYlDUZo7Ee6ecAQmbQbAxNzmX7lDz/irAyZgXSesXL
DqOQNYxJA9GUiwk64EcZBRiDbbj7Xi8+Hfw4ykL4SRAL+tVZDmh4nhPw0+VLRz1kcfAY7YENEQwL
aMjUndAMkTkPLNsyDUSxsPBzFQav5sXSnrabLJYhryLT/3G6UZzlAwJCSakO3Er6RDjzsS4Z7jae
rZTIeg6ulvY8jF7Xie55mZpK1cDDrd0LmlVG/VEMfnMgI7ISG/dSLXUJa8CHwgU9hNOAIWByheVF
iDCQPyX/rd1GOuONlEuKAQDC6x1WHO0z0yU+yTi0B9O41why3TaR5w8oS+qTkZ8yPqBgeaauMcYx
6ZdVCcU/6ts6vljeAXRhsnBLoGYanzEdNBppWW2Hl5ERu1YQB3Eznao5WctmMknCRbuvsfGvBhWD
14MlbtLVTDda3f7F4XVtk97FTClM9ixomIojkYUz6qd/jM+J0Exx4uivOtZQIsPYVGq4fGZJSka5
MjWidwUtWiKTtScASZKsJ8kO+ACpwhRfYTy2f3EqyR+S7iHLSRXoSipAgtqM7xqnKagvnKbKGEM1
k8ln5M+nbl9ViudDpORmbbo6BjPMS6c9L/6MMCihcVHZgN7SdHyafSUI5I0xdgFzMc0JbB5kyzyb
v0vbRlwx7PKa9SdHusN8j4K/ugXVS0brtleaqlCVhTFIv4aPOmQe4h+99ElVcncXjCKN2JzVa1Rq
ybqILQ2aLUk4a9AEzyhCqc3f9O5elEj6vUxY10CaxES9XlP8X8Fcfzd6S7owHx9bD3XBI2zfkfK4
KdeC39C9Df16QEUdrxmQ/9FqUFqsaUcTOUIh9Vq9EaRybYh7A+2th8lcUUiD7OHPQfYMGFkPGkkx
vGMiq+JzFNGotbfQI5X2SsRdIe5gWarCXnQWf2Rnk85L1JNGlk16KknsoDxx5BSoleqcfSFWpx74
FetbtLWyRyc+R9UM7FpX/GyFiOl7+uvT/aRbMKj1ALi/ckBcdFc/ffgJTTwDAvNtvdyS1y5vbU8h
moJo7BAcd8XwL3kOiFRZbpbJXAn3cllBOnmcbuxbwuieBpbMIhjWQgc8FruXCr0B+yT1BPHgsGJF
kOkt5ocds/rHxIPbWDTKfpCX2+ljT7+0vwCLQIjNBGyvaVoBQVHc1AGm+LeaPGtl57Lxxbs7VjzV
XyUxHLzhN9BCtTkPjldZXm7+fjfXQg3XOUJuZTcW+usytAQ6dzNomoQmAKJOtcpj1OJ7lo7AQeIW
7oPzsoOhYM7iBF8lUaxGKPDW6PRn4lXhRalE45dv4TdaCz5fB6gxPHGFWHXDqWVR1yYzh3L1Dxmv
6IZxKo/ARn/MQv7zZfeKxCcBitjieHFvA9LN4WOLIGMKFba6w/2fPKyFeIbribvlHtEbCegkh1Ym
bi2LfUJjHXkBJeWBIF606X5p/kybXWLWGatpky1/xhRbDrGhDYavr7Q+ol5P9jsn7vNsWr3y1MH5
HVKOAbdZy2KW5B6uNUKKfRqnrK8+H2D+YLQ4xHiLbxAIEsb3jdjSWVFZF8ro5AAWEdhnozBQ+GvS
8etyA7BozzCjhSjRFtTnE+d9DIm2eWF1HIS+liV0ad8sg/A0Dec9UVw97dxdMTAeK6GVg9hZlTVu
CYOGMt1XjGq2n39BGAaoTFP5I5YUUJz5i0Kosocc+U2b2IDPvaslSM63z7fiGxni3b9PWgBx6ov1
ByZ8X3Ik2GA3JOn/wjGATVzmk1snOkgOSHHHVpzUgfATb/2Y09wtGNVR8xlidvHG80ojpZJnrks5
HBG5493bOBCYiaJCGQIfDdC6tEcJoLFmSxwmwsbyUtZafgk4ZhaxQy3zcvpVlBp/trqSKU0brs+B
LII5VHlFdEsWpTi24oeWXrMOpL9BSsBS+TwjwaDxbEQzHds/h8XumJzk4njbPWw/YjFozKHZyrfY
ViG6thbL7wyPSMrVMD5YL3WbD89RvhFfcZA8kzj+iksqkIsozFhicmm+TEEs1zw7jGXPW5YnB3WM
D9VG6j/yvGXAIgGPWQj+derwEroT+g0eGiZXT2WjkwE+HbX2ELHOMUsmDZT05x9Yw/KW97rbfkyk
J+8oqfit9yUZrwK7aY0q8BaZX8R4ZBNqFxvlI1LpcjRqsYAMOzVabt3+gcf/7jspTLwofsNLAtZk
Nvd3q18kFtnI7B4tApxPZ6gUhLD7J6yweiIwA66hzZYGdZ6PQX5nZhcqkDVsMIHXWy+FMHA1mMtX
muaxneQJFjyeZx9dmTQnIHgLMoBlvTow52m1Aw9XXgomXB+IsNBEIOiYhpWymgCU0cRkFku8FzAf
vlYToIKDF/PHi00EMICvVmoA0SJthdsms3/tW2VBh197ZFsV1uFYaQEkD1mQL4knFfCNh59QE/bX
8KwTO99zy3ZT8/NR9do4Hl8Y1c5J5N9rWzof4+Tgw6i0Zn1k8ro4gLdqAPARV9bQnxsXt9yPd6G4
NwaTn7UBqxVY1SJYVcPGFGhVZeeHvcw/HhKF/DICMsK26Dyn27ALXnFmC+cMXlsYgOUV9iFT7NFf
8N3tQHy8IbTHIEVWJ7g4H4K8kteGDkVnk3mLHVKagDAguwWMDJlJQPKhBoV9zb+OTCd9I3b6T5Sy
pHSNszrUt0mdczE0upyNjlAyKvMX9ZgvVGLacG0JC7fGjI5yqbAPQD/7c+Gn1bqhdF4wH4JpkGLz
f35qMjMTiyjpOpIh5106Y4FcovAu791ZhHcnx3yvx+rDa6w9+Fh6Gl556iS+EKnn/qdBpd4VSv6A
oQHqsLzdyzUb+rI6JQVzq+lGebyFQLp0aWFYnO7OIJ9awvDVpH7gIyXy5Ypku6i2/K0kEoJZ/IwL
I1/jDIAR684IexYi/acnrOtTBBchCZauKVhUYR8Pgfmc4HrY6b9cTmHciRH1NAIr8rwOZ6a+6Npv
Fof8rr6dsjjuOrwrFFObkCH3AbnraLni5+kWJdS4s/ewppQrovUSktk3wYKFi/dAG7gWLlFNwhw9
HbUGXrVyjYyup/jk0/Ap6DLa//dWU6zShdMA983zimiYHYE456fgpBoDJOFPLEa+A3vODuVwslSV
oNs3GSGsfaqW98pjqUIKsclL9d5wZi/+Vh4bqaFaOwZCnGvKek8S0ddXFCwBQ5NcgmPy64TCWMAw
ZP+MHRhfAa0EUdf34ybOMDGYpnzG1Bk5yhV2eSEKRV1CiiJmqEizYDnyDKjWbrKPq5xEqHvtjQDy
rmxpKTohFtejieIcQZ/3D3kRcjKtd4WLRAZ0CxGaAiq4pT21FdASEtm8BDouAfXl6skvpuOEtK2l
2jPy3czTyaQ7Nxp9SM0t4zWnci+r2nBD9a89iNWkzsjxNyDEWdDc9xKObf1yGe5a+A/JH0PGBAmB
hSwu/9fsEcAmLkgRl4bFNwA6pipCjqZ44BOAIAg2WnQSmABDx2rIJpPJJzRJY5mEMzrSP+9LW46U
/7iNBCQZLh5Gp7yvXPapHSBkadj1cF2K1B0o//QqX3xtZXW3DrdL9pu+fye7qSrMKbAupK1Gq+t9
sxMeRTujMFuv6k5E1FeJJuphKzRcoac2yYj200mSrEuK32TRCfCgmQAcMcUZPIknikD5rjf7Ie43
vNyilKWrd29BEyfzSQ4aaHw8MHgILm+m8Uw188a4ze8FNgaGDrfZg55B4Mv7CH28nZay2SBPmhOR
V7yl0Ysnf7/9CXoMmanVAgb92FvX7k0Svf0rMqmSWirQ/HO9cMZtXAjNCZ7z9fQQczHuHGxH/l9a
5nm/lcbGhLFVuO1t/rt+ow8LCJqrTawGBao//ciimg7WAD5kUDlPBOusnXLWztcVcPSiX5Q5TEbd
zpluNv3aF3GhJQbV9QWeblt0Dla7YoEG/jzchuRblRkW/6UhqTDwWnlBfG4jZvZy1MAqku13wLO7
T7oSc0awXAwwrtHroUwxTlOmP5mreGrz5D5zKZQmXArKuzi7+TEbfgItm1sXmr/HfVGbHtz85HKm
A7nUWIcwMSIyYVxizsYVUbWY4zyIqRfU48Pon3r07ORewmiwEs89NeZvRd1bhdnjTwYIp1dThzBh
abjKoPJptRovY4WNuZfTMJ82KM0/uT9tGmN/e6r3kDC01ETmYhy+mcWHLl8SMBcgpeLaiJSvozzB
i8p/tZDHZhKFHpO8E05+4Mv1FMKNqzPQxkAhCgBpB0sdkzJc83ltj0Im3BxeTKG6kMseUG63Tt/v
KiHpqWxF/zSN8MTpQQ5+7O6x/jKyziLgMcnye8wKRVLu6mSpRpBoL3S/KvTW801ksfAIDIJ778d7
A838SPIvf7foC0RWjgex6JQ16RmnY3S6QoQG4FVJDm7/ikymCVAIxLoYCbWa8gVIrSAUDkebxPvX
zq09ttrwMQ5WvQMVoESk1MF4tLGikR9hVYLa1YyoIygWagPLfwbWaq3atT63xi+8v3KVl7m+9IPi
VylCdgeTxdUaSV4je/8OLYbbVHTWg1nBtIDS4DZKJ6eAamukicQasQ2lsgEPldqPAVrvtJzCCDyr
HrwbikgzBPq+24C1wsgBVYKhOVhP8T/I7qcFCrOJ191xpCvYWTWjCSFNJR3g+OZgEX/k/yDg5d5J
a9k2l0l7Rcj9QLARaLkRHn0GJ9+pokf+2KW7ZSh37r8LUOfmDf319EXmlRkGG2ezYLwAN3TdWcn0
SGASiHGe24zc8Xr83Qiig8m7e2TLAzc2VadG81aapAvczxG1YKa790eQSG6f4dr2WE4j/aT0mJgw
YStb7lA6C49rghDQm73755xashAkEKpaub335pBgB4AIHGvUF+v4kdatXyjV5eY8x/MH7l3pUdM8
n++0iPwAP20uCU6X2vbsBsz7lXI8KtZ9dEzLe9QLkOpwCW4EHCYSSI8kNRYrQvhGUqIoL1VMzBp6
W/2wK/9dWcbJkFxalT2j5ZmKjJElQY4FeNrpPN388iFSX6t/HWfP+Z4qqqTVQp3ISoXDnQ9ODVbR
1vS1l5S9Fj0o08SJ4ncHpoaRyo3Kovuejuz2E4OPFjZWFepkP/vbdlBmYN6NnQBWchjVMbrphE8+
XGwW0PrGfc50mhZcyyHfiiLfrIkjOVwVHXG3Tazm5xdiK+L9xJgE2GqguhhFRBzYkPWLec45/mAc
p3mAwBTAQotARjAUxZGV99qB68eApn0seJix6vE4c3Xr5kgXiPi1Cav5Z2Ob6tAekrR2SnrJX8ac
YcGWZo7ksclmEJp3hJXlCZ/3bLfr+QapRiWqgxYdSgD7t83rbOfBUG/+53HRmRUHO+pn86QTlmjF
oMWGBJIR46SdHMLLSEBVVYdMcWNAYj1DCjsCObYBLH58ixqGCFxiZdZ7wH1dI3NEZK6IPir2GP9l
C+UBR2ofQuaJr02FwENP8uXBpCZ0VSejCGbJKfSeJzSKEVUgNzs0rNPOksP204GMW6EG5HCjReTM
iUBf5iOSIUTr+oKkHpnK7Sd2vQqybJgHsM21W1IxHdVA5O3dACEupxozR/eY1L151gzFm48tk5bw
sD9LTIUQVgmVgrb1GQg6nOxMudiGcFK3tLPV62j5UMaCQLgde1J704R47rB/PjKGK2E9YJ3bk+6N
Omg4//Lcpg1RL+isgh2tCw18z/wIjgH63UYNq6PN0txGIgQThlEGbPp+LzYQxSdZx4LfTb3/Q6E4
wQ/OFFOQYtW4fdV5vLhoUXlJ/hui7NQnpKDcAD9W1hUR3cJJnRqzmvce0UxFKtaAkNBKPvxYRMCO
QzFnfd8dzVSMb+UGHbTKepbvr3sarLvSETNhNW4B1V5oQ7xszcxI5yWtgOxOXBD57oqlqRK1qT5L
a/af4eNeKS/y0ZCeDEvfsqy9KwjquVVqpHw+5UOtPMEPu04Odc/WWnE+rCLD3KMZ72G42b19k4Kw
FiyTrSBj/IsGZmIxtmCDYN3dQqc3kcfZ61Mhqzv2gPu0kQpBNbqJZht34Oc+Ea2pVkn78mGkJX+0
lq2kneSiQy0l+a97AtfVPEWv5DJVTeRbGGt2jI2Ch3tdevr3RgoEwwSw8OVnwdrlxg13ejj6Wu5y
vzmcnd+maPO3eKVKUk8L4xqmQV3Z4kUjDgn9Y2vEDNgw0pA8rC4KDBSRCZ4u5CIodlxQMBIt02LQ
mMfWflfeL+ii2K1x6RfUBdix5F11Dp98NslPV+kWer9ZI6pzSQ5jQ6QvXOzun2L+kymKn0asqQxr
kNQCOwXKZXv9PSOFeXT/ujlVqJ0b1sE7iNaK3oZH+tQAUURhB+G5h3ugnsWOV8hwB9RWEQXtG0sk
K72mqFz5KM9KP4sFfIcHc443w5pDUeYEBXdMpkZpKKhI2YC1sltnJV/VkNgqWZn9xbH/GpbxdF1h
TTfBhYW+DvX1qGzSFI3/OH7gC6i5b4UlcCxJIpvYAlx0gXkzYosSv7GR4che4Z1pPFyjGpcR0A6G
SJBjLoBMlhwqTJ8rhuKr6JEoeASRt3YIR+bLBKd0TANtGXL2K7A+I3CercMUuccPQjUByzkflDoi
5RUj2mP//umRVK/BQ1tXZm+mfBT6dIcHuuNRBk4TlbyyEePmU7KioenyW4PJzM4wC0ZPEBF2OVrK
yiUou6latc9ZqnVB+KnoPdt5Dul3Z1YwwLP7g9qT9BuMuTq3A3WQpTcK1GAHHOFPZ5Y5gJC76XPv
0s8hJCq246QXpPdFVyMX5I4GadtYIT8rhLy22AAdW9WxXvPpg0zaqJ5+b+ZoLAtM/5bTXjg0pLZR
G75mJptPyt9etMBf/eT3zjnHM/IcywtWRUrYPpjTMl/YDW9a+9usSQxzbu9Lr+wu6x3fdrsvmWJS
TITxY6Rupw4Y5LC0WtKtqmwk6ACrRtG/qYZuwDnjoq2rff0eP0QaxrcBcNl5ZmJbLwiulkSZRg/2
PV+8R/OxmNvFzZpwqTY8uonaFihBKJffyvjXUNhTqyQgBa19enstPt//4EacfGG8FLu45rCcrdtS
VPRJrhFNolA27OwEK4/MzTRBVbTZ862sn35Y0E4JSyiKeIfMhAXnwjstK+05xJHN38oFT/KzBH78
/A3qddG+vMxUZ7UfdQExJMVGo5/IziYQcNpdKl+UpKjz9XA3PoI0+KNNaJq+xVPKDTq+i2ArKt9+
mYh2I66eGIRv0Idsa5IlDNFZ4O6DhfyRHWVvyI8T2yNQy22cPEXQ9iC05/umVhIHV464zY3idzmD
oEbPZ3NdaVJ4SQDFtyaWUMBs3QBiPZpmuC6M3H2UkYfvzZUVvxYlKlcc+HtJcHQjGHls1x6oTKwg
0ikCFpuzyzuWAm3igGlcTT5mJvQ0OFUPHY99a8D5Tfu5bwcaJs2kNfKYsUi2HmJpMwVFaLTRSS/M
o2/rQeRStITi+DlV26xM4bpvC/0uawms5eOvZq6rXWRYtOzdaiqYB+5tql5TaHXYKNzR4DnGGg71
ooxbZ6bWdCUCI0ljV5hT5pBFdzpdZi3CvBvrD2HPjSMReouVB5v4j4bn8BwFHMvqgnrikd8aaIiE
qSRm9iXucPDuSxWKIKBHHVfSVmudxBg4K5gTw4/9Glgl5hB+tHJhY0ZyT+UzvNLhkKO2t4KJtt4a
TAzNpevmtipsr2zrK4HsqLC20vtb6noeeuD+RjPdIqiNPs8u99DJnLFRY1+SNL0t9325wzjWU5mf
Y5lLOg1vF+G8gN31Y+u0P+YfWiuxEjbKNVRDfiCwBD5DVPuT1LK++rPPDT6Be9iAh9zu61/dbL6f
6lR8lmwMwKiP8/RzNPnLcZ8CFlXiV8QfLvs37nDZOKOeIffchRP+SKsureRNC+yckcP3q5zhlcC7
/ihUneYMRUU9QO2u0Ie0ALFZONDd2TTzwqnexpJFdWmtUbVooIV9p2CehJV+eBel57JMKMAmjvY1
SvZlfvtuvfmsO/d1fS8a5VrBOsJ+6CPwWTnQnoRnxjh3mqLJQgH/Vgy7uOCfHGi5sEY+WdB6a5Gn
L++ULeAnDEeQyKULG8C8zY9stMXVdKoMQ2D9hInMxTcIZZS/OgfytZpz1y88C6VVqv71c6XOXzQl
uP6PD3T/R0UFbClPB9hOcn67qZKojnmmT5KQQUZDnPK/ekqPb/gSm6sxVhXIXtVLbOHYEkUrHSUT
iRQfPNehPzK34RY7tbBu7YCg5Tz3thU4owEvMiclWgegTN+oeLR7cSwVZdYgWRkHCT5yKsWIvVD5
nkY5KgjSaDXpPixt+doFSIPCxE2CyL+McR40OUJA1r/fkGPQc998m5V94hHdCB3U0TnyBlh8OXMD
2gqoxomfhimgJqBhgPd5ADSxtSCazZjTio61pcSVRsBvZz3CuizK7nOLRFBST//2PPRvbVEBJ1IN
99VurhaxJ08tsYAb10qWuoOIiQzKglWIEr3VpdX1jX9YD8MncS1JTQC+YciM83kHXiY1J5kW77IZ
t/XYTIjPzLGSHqPNDfoTe6nYTifKn0toqAyXeR+eEIkC1D4yTo6aoRKIURQkgQ9dpro+RrQEz9j4
aUugw4h0e6j5KlEHcCK2aDkY35U/NJ4sWAO2UFv+muxTrRFIUcHBGjLzQpIWEr6JrIXHptguq1VV
578OfV4Ws8jrF+pGn5U7hFnLaisJKJu3Wcg8RZOBxHCzIi9idzY5z7cbk8BlF8w9bYOqiCMxpHzR
woKBG7x+nrOC182KNZwhGA6HNipidzNY5mGt04U1xOAlwVnbfnxCZ2cZLPB0B16hYBLibj9vLezQ
U/EI5Xx9a1Xlok/g+ZdBUWTkQ44xsG4AdPBqa5YwUK1nI9EIs6yzbEQxQ0/BDeBELoIWOTm74zqt
Nf5sioUtCkKMTogB8neu59VKqkganNSYNrbioAGNXFJnGxQpvyE9x0Fk4Vz/A5S2b7KhsaKSv5aB
QoyffQllNUdJX8fRdgOU+97v60tfRg2LjViEsyUR72Delx50PR9LeqxApZDBJ3iI5fIWKJ9Wq6oW
wsuMyOzx/UIRZdZaAfDeMglvL0FYogL5n/sJ7XwWcQiQtBkaThnb66R77kVQLZ7fUn4/049U0UrG
m0Qf9UNT+SQPqlF/+57pC2WbEqikWxDdlNQEhfupxyi6Auw4ct8oLVLo7bxZYnPUDzECHA/lL364
QvCX/ZOqgAlgR4dODZL2YlYo0+agYn+be/2CT5YOaw4SopzP22KnOz/srSJq+2BaP/sSZnjTr6PI
jrKEfA2x8ESJhJ1iqbdc+z5uMxXIgSemBIUuQ/he2ftDXl5umCCYPoWCIyJNMB2P6dL8H8Bj6LY8
JV5iQDYGaa84UuIzsSYo++ccp8KjQ8PwmjaF/oMUF+suA7sa10YuX4p4KPrpwdI7PvRi6fZrchD+
vF/JuKr+8wn6HwCmJB3lqN4LIcI3gdrf2iFtPO8wprmoSUdM7nWhdHw1Tk5kPSPlsSOJpPmoXIN/
yL1aXAqhoqkajIr3Hr5PxeHOQC67K8vGo80PbXMWhi10gqVedOc5fGSoaVKMSOJJX740XQFsbvjL
uATPsZ9/FqA2UAOUPxHBBE3iEUbHfZN1coLlGQxrDTSd31+AAbYOuT0/G314YbqNBoofPneJnJXC
fONy+JP62ow7VTYibG4cvtHzL8lx8BVGKkuScmbjvnM5bxz8ZxJssst4yTufzZGDrj8IeVMAG8aP
bpxks+x7lFUZ4VXxUwcobj3w4xEebUzCRkaKVk2U6SiNuMJXKTfwpwXqXs5W8QOCmwTwBdTRkBdS
6RTus1FlS6kvpvrQ+v2BvSUAudD2aP0HF8CUNzHAyLKI0cI5/fv54HQdBrlUqWOdw+W6XfWGpucq
oBFlJMdCdrroX06z//V1tQrEVsgcMCJsWMQZ81+neve3eVQ6+vGjbKTB5xZoUIICz+WZatfLd9a3
pkgkMJEZMleMBKENxKUCxbFTtIrJxF/hGl4L18mUZS1jbd5VwDOjn+yVXOdySdhue7d4Vn2X2zSB
7ji+168b+G+HEd7kK6jFWmvqzFWP8g4g0E5DT+9c3UVzbJ/LZW9+IAxBXGwcVdkCqAq0ejDjNK3O
j9LQH3DCeXhsbw/Zz0WBn+SmwjMKGwofIoyJFxbQB70ztHMSjRPqbGYF688NHbWurm0HkO3J4Psf
a9JSQ0UFiHzDDn08sMxELjfmWksYp/lk+/sPVMV8zfIYED/PvNdBTNGmhIKdzmk09rCRudN3Iajw
NwL3Q392fiOce33IdqxZDJ/BCz1K8WTQ7zzrwcN/cYaDU3LQAk1vXgpS5ANaLWKXVziRp/jaEzqa
0d0F+z6BSRGKHMw6CGPuMXwvzalSlw1DoKkm6twkvH/oG7oCBnjhdhSYzNLbKc5+TkP+eW5O9KJ7
DK+1Z9f4kKoJxHqyVci0i4Tk4WyeavhEpBpPmqYf2oQDhN3gzgM8zJ7o2LERoG0SVKIpAyMoPAzt
4lWEemTaFLz0HQ5DZH47Svz9XkBwjpO+SqfO3O/pJmj4jnhsm4KZwK2ixj9YjSaNoYRNLqEBxlou
9Qo5wGmUjKC59UMN2YgWZrQb5XPduAFdyLAp9yPSHrU7Yxs1lT/M82zBSxCxJGC+MChNKRIGDTPC
tn51DMhhGXrTfjxcqfm9FIVdzmhUAtGq5E/syaNDqR222PM05jly8b5vXflXs5BHtDatzN2n2KAz
CW0hTlH5fEXIUbyUyXclp2TEYC4nWKz0zXL+DQDlaRT/aYYid6rZtGonVFV2SgVUL2CuJ0AUJPnb
U/q9AbgD7c/iaxEAq6WI6l69aON5CYKN69GVl5kG/5WG8iDZYWUMk3SVZEquHl8auVT5NlXAbqae
6vD8UnQ+NV3x5KPsodQoc5gbwuFoSEcLRyxPIm3J9vMbh/Lb0X+FQfLoUkf+6pnFCfquGsqQzGTD
auDukrVonMkH1YFTCUbfpEZz+kg9bhXkYs9JeNFKRAfEMzskP3d5wzePrRjSBX1VsWhRkCcma7Kb
5Tp+jNvzNauy1e/z8ONUxsh2rEZIltwy7+R6vqV3GsLVkMxxI58hNP2sj55CjYxPNlxUoLAVMnEl
40IEwVc0jroIyLBmZryCCG3TXBycIrj35IF9VF7N3O557Optc6sj2vUUVG2lYDu0lMxcVQOrbFmb
1MTp0WcLy9mDMT2+D2nqkixNx0dcl9aII7Jl0hQqXVPxrum4djY/LJ36r/SC+tuw/z2OavmGl1G2
3OODOnIGmY+A77ykAXQT9L1uTiYc15+MAjiq/9muADsyMrVNNXXkU4aofD/wP48eSpgtjKKJ4/Rn
ueWBe192iXn2rW/rAE+/WV6B0ZvCpSS7OeeyeBXVwM7qBZ2ewr3WTT9cGiAE8OZ8I1TJIantci44
W4Uyw41NpAxLbayErQRQXiukFpRdTc8Cg6WGGLq7FEnHJ63H1HNfZ7QkVPuLQRDmPnC+7cD0hE33
ib2cidHbkpby1z+a/GHMt8Y/RPrhBAijlO1LqXQh0DaO7D+j+aU2ZMRSWIx/Z12rmcfp+E9YgBR9
zAbJLJf6/LhhQan2NQgLAnD6RZyZi10+Q+JtvsIsikBR2fTFiTXmvBIT4yT+ywQPZEwZkxDzt2R3
ybzQZykti34Gf7bjWR72XTHKfez0em4zNFJpmg1cYSzp+DUyqh055qO1Zf50NyuDqPoL0q7n4Gj+
C6vSCcmpQ7EzMBu9ONUVKivIxYTN8hG9sIoL5qY6JJGj13BH94CnI0a6R63GKrZvaVgj5MYJ43OG
hPKaQnkid8BLoZah5KuADsyBSCgSyP22nR07rHV1S8djnGG6QalzmE0S/7Cbzyoaw/153zoPY7UC
Ll0HG3HDaB84MsbnVY2qZuxy98zpf0VqQEyfgYBJWrbUs0bjh3abBGnOozcaCf61tjWhr+fs839e
cEHwDQ4e4IRqR8RBUppHNvamAMWGUgZiqgYnZ3xHsxQFLdmca92mkkIyb53wb0m+hVdIxXvkC+0N
mNCb6k4MxpFc+4DVEvV97Cxv8QxgR1ZKuWb3PXWPc9BxgSgaCdXQcobp9JucTgW/xl1lLXCMYXxf
1x/Jal7nlC3FCHu+NdH35lSdY3122c7HmUm6dhodTAj4eScSb3jzEzfDPC2rxD7IdmY9UjH4knfv
75/Yx8xDASdkwvvrv9BYPRCFPpSFXwG/tXSsnH/QNZfnMmYA8UtKpnk3ZrqWKWucw7Q7b8ZzFq4x
l5BzIiSk5J4H7oNwkoWTIF76Cv+ToxUVYYYq5+uknqc2QmucADRaMm8qvOrk7mJZE5aL86JcpPlr
70WW6QGUHJ54cFhHAgX+bCrCiMA4pGZlQsGzPQa4q1gCdyRux+K3JDMqUCCM2aym6fuGlzTS9di4
pAaANoj9KIqwoAaEw1ZNDk+qURTVX3YiD6+6cFXqd/ZHEa1WUPWoCTGLAv02AlLYztwHx8QkM+uL
VNe8D0W8z72BhdgkStFs9UqH1d+Nl6vUcko7/66tGSBDOy0KrJkR+ELPsQ6blkv7lcPVHd+gasIE
zCCAgCrAuyKofkePSR5wCw3vXzOjCP4/q1uXMpBY6gUNSyys1z1FO0S53dpVt0DortvOoXW51VTS
RodjQVSsAfVpy2QEu+bzkT85JSvhEPo7QaA91wEBtNQ1gG2zy5AVwMy87vnwqwaDKN98hiH4/wnQ
iT4UoFyzNrOclly7j8KABvkP1e25OjdjKMdx7rMgw6QRjOzrKkfjtnuugS+2mjfM3kV3Kh4ZZH8m
yhcaYrBIMWIaZ3FV0wdVuMbUkMvy8/uPH/PpJUvUFc5WFcTs6XMhCrHfJcvMhX8ROsQBrlSm0rXz
w8tpJxKulsJjtUd6u8ZA/IIQ+eJa+zNk6OE2mdAIoOXKb1T1QHWpfGi+jCZAvrDZ7zci6PPag3iE
Dsra1XP0Etj/ScM1F3SybhD8iAKMFIKyzmQEx6bJP/40ZFvEvDIvpIcDEx9ltPM9ZZqHJ4YfOqnX
XF2xNb7KxpSbAVdQY9V7D4Tz+beOWgVVTUo4uWLlKpcKqTgnEr+K8mRRGk8+h/GKcAGMfFGXwje1
b6g6gS03yOY2UETPtto6hwQI50jEajU1fW4xu3v3eXjZ2f23fmx2UlkmmzaRsiFfvc5SE1tceBGw
8UYzO+3kfFiZ3aPkBJSeDjtDyWVTFuTfGvVhuVA6C5BnTDIjerLaeD3M5vpxLev8eUsDB8nk/C3s
5V0ozopeeEtf7yWbOt6xvt5wP94MYw2Ay3moYESAuwcqgOjzl49dxGMntnYMSeK45kDzXrPBFhZg
MvSRTGZ73ozrYAAuksr92BVo42+La7JLorEQEU+nN8u6d8Y/lTywKhvvEztYwOy/0CbweIjqAyDn
vX74wiiSzEh3cwhP2OyYpC7yOoc28LezX6XFjy9eWMvrMxdVyl1EAp47XGpXHESJRJ1AS37P0ien
TRmRpxad3ya+ENJYUHnLqXeIRuhgahm9UvzMTA08ctUtS6/6/eWmZ0Kamc/prrnqzlvZyaKIodVY
gjPuRaMEdFbV7VJIxTcl6KBeI/aBOrPW5WtB49HZgBsiq2716dxTSLVRjBeZ86FdaaJathgzG11n
5xyNU/GZZHdjWxXqPtIJIWwRHa2jqur6y/4eyXVx3cvesbKo7FN2ZyeDvh7d0daH69ImPSud8eq7
zZUiKtj5Fg9vEWhuXJYKQUvWnbMOK65kZS5Vqi9YK/0AaRC/pIsXphMD8QLiBiwpgLQcAExUr5fe
vmNWExev9L8JZQFF9q4dDmRgo2cG9iwKVjCih8ruzhoGLq7LmO7zHMIPdFXj5vvWZqZQdKyxUy41
MEpZfmLt46XDtUIIImCO622eRyzUAlpuBF+zodtyF6IFaGUnK4WmaVYmY8x8WCbaynL/ZG60Trnl
qhzIjuy632VZozZem5YlhfUNLSCgXavR5JP/voVA7OnZvt7ha5gUM4QVeLu9v4xVPs/M0l+/H+qJ
/TOQo3dImdDlcXBNLruVHQ7O459pVQ/iuxzw2tLOk1nBXb0A2/HYeNu838uk0xW1Nz0OUGX9rvXq
SNLBOUviFawl88zEffR7muo79cd9dwHuncpTWqrVN1K1ANATpbr0MOqZm8O/vk632ukRiAn5bkNX
UkvRqSHA08dDNrnXQqAagwQgWpBD23qCd/nks0nsprZ9nlT5X3tMeBA9/Re0ViOLfgMlrrEbCiMU
yrnOn/rAEiWN3yGxp8clMCG1qnKY0VS4FpgByRslskzIj0ggUV/NSe7TU56qlSUAdeYtO9wfmKOc
WKIdzQ7lCTqFvKV4V5d5JdENOAshDHD9ILUqvneAvl1fWjmuWFkgcoqkWZpX/8HyvuDdHvj+z429
fwliI7g6phoCGAikfWvBvOAqknhrhWjy6ryqurQ2xIDRduZkYkhbjkyahHoxvkba6uyOqrlGH3LJ
eDBmk+4aKZGr8WgcVCatr/7nFK82IJyIRrmpUk3l4uHraPBRbmbORqpepC6Cxw7CUAzQqfbdT93B
T7URRMNT4MWsnr9i+szgTOhlpeXfQa22qW4nMVk9BCon8IqC5ghR2w5pPfBrRcQQo14U7qg52CYm
9Gh2Pw4vi8YdLXlm83YSWGRrW7Nu9DqkN5ngubX6S/lfng9XwK7BvFK8AVLhRoykpytr76cqnZVO
WEiWm7Tq9VotDrsCIfkUUElZpbuHs1GT/RLUyEc3/5j5sHgNClm8vxNKhVTwc3Km+1TXqQyPFb5C
I0SPMLbYDk0h6tJ2hsfVlgyQVTAP7+jYNAbb5ygdzAHPqDIxuzM6QS0Sx+vuScARh651NA/IfhUa
tlCVWGxXC7myOFATgYtz1uJzyjj+wauzHt9YzoimbNijxykw4wLOzTtF4laVQxzaRjmO19HIv3ZE
eQPk+EDMvPAmFukWsFlFdHRdr4S3qZRhoYGVPnLGsamvtbLPQqizzJ82+3McFekvWRke9yGox9sH
8Op9lyHXcg2ZClC7d25I2ScM+oWpdWAWzGkvraWzCdysRRQ7TjQVpD/eJ4H3+IGyK3VtnOwDcszg
VhucPPR4fvsUaX09VuvQew/KHyV9ttuUBAT/7WwQ0vjwELWpGSpPWLY9EEFOiy7eWfNvuo6nSPAg
v/tj5WOPKpuRPPTHdQnvAfqyLBNPVBIwEeTW4j5LDCOLA2goNWnetPcKwHu369wrW6wh6p4pws/N
+wg8tpeC9j8koZl/cV+74pllmvshqcnhANl/bcQzpYytOEtV+maiX+QdY2S9tzsTs/HPUJsunp6E
sb63hf9pqWyQOqXg/gi9sa+LBKdkmwYemMqZZjXx1b/89jo4s9KFk30CRQOfxF8LD2rXE76IMHWV
CSc+OP28WESuhJWh7lN0tfKKpb91wlXbK50AOIS2MVdWy6GT3s2xXeSZjMF/3sHO97GHcOC0U1F1
xHhqHNTkVokXDv3r3Z3B2mTMyl8xrsvzoPopnHyvTAPsuiTcKbK1OzmCrLWc5lEAD8mYfnPiHwpF
2W2BV3COxqcUJu30iGI8PJr5srRERRF5DmnATRdNoQQ5DTDOgxklXsDPxiCCgS/dFh/BZsnzZlHH
Y+b0wmImQmKI/FjQZBtA3v92HeStVSKXvavSMON2CqarrAzTKZatQUCqTPBgCo6iO17lzcs/7fvt
tr8gy0t2cjxeilmy5KPHtS3ZvvOTT3Iu/s5h57vclXUo8Bwqart2PHxbKfbV+F2eI8XmZ6/rPgDz
liMckFr6pOJLLxWvwwDHrq+j6jO6DiJbgKDxjPL7s/SoaQhpW6WAicAxpU0k44V1y6hasJ60kk3A
PxLSyryKgbTjlVY5ue/9mlvvoMLCpMCOXYMW/577dHMoDFroJCkWE246qOIyAkG3UxXkjjE23WZ9
xuia/4ebyxr5ReMFhkuSAa3dLpQaectavfbSrgmOcbuE+rDwVy7BZJe3c+GeDWOlISDuI/aNSHey
m20vmQVZj45LJx3+6UmUkz4RhXHGUUMPLFQd0IVQlNHG3xV7AqTtt/CdCAqSSFiooRx1gXnheGUF
CU5JaK36nIPOPsmgTz28ta/U9izudqWObrhdZFGl4s4syYL7lKAuDUnvTrfdK1vu4o1wB4x5TT8g
dcwlccRgfkDJsUm+0fJURg61K4aLmctNED3W7EFkrOWBdLOpMS0Fbxq8LmnlT4cMb8nGBEE3PRbi
8COisYhKbwmQmY5y4Vby5TK/QYzymQkcITRGB/l5csNA8GAV7CErHszeTSNEluUXqZRH2WEPBA9C
XP7F/Ys31zddf8vTsx3TS61Dc3XDzY2AJtjey8T70euUIp6gXWswFSf2VxlClNUmSLmgs853py6Q
MMiCHwh6vkm//W6/jzHyh1x9bZVy58WPHLDI5YvlMqnLERoI9fTn6qb5sXIff9KLggwBip5TU3NN
+vPZI0KZCTR2zo5Q9H0XP0wbdpG8J25cFS2JvbRNLFTZxJcx98+gifpC0njncKCtLxSP4LuodlOv
uW1BCnKuHnfoRNGbBEYpooqIEwnRQsiFk/ES6PbZu4ZHOOJ6vBTTKxw7N//UqRs6Y4/z81rqvM0W
5Ypsz47y8Se2u0Q8ThIW7G6Qjhh8d6afNmXBHfMWo+IjhevzXqm7BIexPwCQa9u9WCC705rqlXyd
u8gthVlFNZ85QXOuA5kf8AhDEfCm0ts98YkY3jI98O44lhN+MljInJCh5YuWjlnll0+p3mPDFNyv
wceu3SdO6yJjeDQ1kwjzBWdCnJLq/nmdj11okxCCyj99bMWrdaO48QSJaruO79MJA2fsylHMpm0P
7nouBzYLngBCbXcqnQ0flQBLpysHH/aYKqRgj1K/jtmHPMoHpOUs6U8eDAqCEdhkeowdPATf6lOr
LEr9NzFyKfOr8kY8FQuUkbNxu4T5DIVkI9QnLOd/AAHx+Pppl+agBuVn/ZhiR0opCM0L1WZKb9Hr
c4gvUFjh1AYGIHBInDIAR7wABjlYep28Ejsqh0xxzMKTzFqdwXqBDqd/Ozg+svrAejtcUsjJ0N/B
MFExG72u7Arp565ZSgZZhBDgZKQZz7zeUsxAsuwno8iltyj5dhqIOCqJ1/IJEfyBH2j0xOkz67pm
riPOg1A2LgNYP2bklviO7lvve723vgMHQt4Z3UlIwYMm60BAbVYbabhVyOdiClAQq6SSl4O42vA6
S1dLHxzXyWNODpyeqpqtnm7pYHPW3qP5Z5ozPkAnnQneRhvUkkhvVLYWHTLmXW7r615rNkk6XTqN
sBIS6PvtMZ/E82lDeN4Af/ubOHZapFqdTZNHKF3Dk/kUC496j89D1xAh6DPUu+3LboXGaggnnZnX
xsw5Iod4UzFnMnS329P9ScYzJfLmSxMmlexdX2Xp3qZ5EhQeZl4aJKQnceOvGdP7GBAnYN9q12pX
nvNhIJiRDR1vQmIaHnIHUlcmzvtJUxD0Nl4yvKH2YrgJg0bhiI84ayIBeWXwkGrhzqngu2RCB7AK
K6u2luJlhtqBQR58sUt1oooHHN90XMFANPa1pTwYelxOW3TT8kwCNmEqkBD//PP1ZulWOKplKSHI
l8xgnCwBoy2bW8GLwcj1R4ViL9RjH6gtQ39KWy+MDVJgM9cPoZ0BMu0Fq17Bx/5Zp+R0mEumtCnf
pCkvLUuSDlngJDUURUy+aWHS0ta7TC2E+/EYcCbLUFGP4fzAyUEnlqITYlkh+zgx3mcwNRUoIL2a
jfVAUEms2DafYY2HolRz/3hWZMD2bfwxNQvfcIWTmx2egCpJ4TYREPtLLd0j4krcAyVaanhR4SyB
JVnBG10Bb8yEx2/v4S4b2+fNsX6W3BlVDRoyhYM+7XoDOUSU1dtKNOm3FUceRAuGYr6Uj2WZSVER
kTiqeiAbw5BcIbM9OPDo60H6uPJ74jwbrbIWu3hmRua7h+4Xpo0SAX+Ajh8oYinVpcqPezTjHyrH
7lSGgMz4H0y0tjwd7t7hPS6Znuagzxr7UalK0wiN6wTlfK8/L6nO9U5xzAnlhtRu9BWOB1xoJdqD
bFOx4n/78+C5QBMpcbHjhD3Xs19OwR7wsWjGvHhE4h4xOmpg7T7v8TdY68b95Lr4T6+lI4b7UTPG
fizkbiNRO1LgQkz2hH02izm57567kpblpqHwFsbt6EZktyuZ+PVBeKc9rsqJUWFei9/lFsyZZyte
pywQLlTi32snAZUCf2pwVAGmMYV5Ub9NuSFYqLmoMpduWAQM5RYiFxxnKUn+lLSMQ8BFtGQ/o+Ld
IGfCqAXBJLdPMhTu40wKik/rdfg8zXlPv17FriVR+1rH/01IiE7CagZFPONH45DFMGAPqrAz+5Bh
h5qs/csw88dOBiRCs1a2lK6A1kp50eM4h6bHwQFV2djtz820kZs5cbE0cijeODTagh/9TAfb/MGS
O7sMZoGvH2OVFjqzMRJvN5Lk3Vl2Hrl6unPLBDbDPfxccM8QHC10KuBJ/TOe5TUxNNNuPXke7AZR
B0er0U6N1N79BYXsyG6j08aDOyjzgqZs5Wchw40+iPIybyl7GsaEChUy7UK2LvPOzB/qMHjs7tcR
jtnN11ZLwdo93Nl7Vri3QnY67eS7AlDliNlpyRH+EaDNPTazk359DABs8HLcMEjI8fXq86oTiKvW
oiDvJ+APCwIe1tPKmja6NLiEFFUvLzbSk8h/E1RwsZ5BTGBcbbvQlCCRu0ykl4fco0CEc+NeHdw7
BAY54dm5Km4WHcwl3Rx7os0tZDkmeGzQ2Fdf8bZYnQ/X3oNZ4eh1EkMzu0tSprixk103uPXp33pP
+X3n77DBLLjz7/3jW4fpDNIYi5+Py0DdszDx/mkJb2g1Id3rtgZqmzGECzFrb0o8LOUNTHiO24Ch
zj5SVkTkoeZsbre9aMbFOflPZ7AHhgz9rETKEjAcs0rghN+lZGDLVdpkT1P0YGkG6ICDpMGTO6pI
P8F/Ixw6RezPo1fc/c4X3AsVZjX9iomGpmqAt8QTpP5T1q/LOFbXY2y8DuZlees2PFk1zOjByNgL
Uo77Eaa+MotDfz2GKa8/AwlaY9CwgWjNDhdGPSXAQDwy+OCjLGwVeHKiVxJYf4IU7P6hGB4QeoV+
r5c5qnNZiXSiqBJIn6EEQ3/xLO4TLkPxYOmPHq8XoFb9lOn9KujBEQDzTPATro5lEckF5ELi1nh8
m2BeCmvz5Ly1sKPEkQSkqZfnl1IVqu60CjnZK9kthVK9IRpcNf15xtLFy+LRU/qkNMmmI9B3pc8J
XZcU0b5YX2GAjMK8S4vnH7nX6fzWl6qDvtSzQ1KAEqMgysvXxGIzAFayecoA48LzqcH+4H9AEfT3
+iFGaAdrDvwXKL7mbwcTCuq68mt2aftzpj4JWDj4LruVLSJTw4gig7FEEirfkbZ8usEIOF3cflCa
io/Gu4vtdtHSk0IknZnYVecwOewUVPQGEsfcDBOqbD2xb/gdUkPzBv/My0JR98eZj5FbJCDGhPjz
TDtDIooUXk6FEchxR/UsmCwk2e3mFOPjwzoOI1pzE+Q0EGHl2Pi0ntxM+AGmdu1dCu0r6VOpJ/gh
9cLzma/lrBi6yVKVZu+7i8p8WnnscoRfMPmfvqAXj+QInE6S9c1K4v4Dqi1z14Ipq3tBSkYmeVYu
rFRsrqI4oYR3MQmKJTfCeQSsuZDPBNGK87lR64dX7V81im10Tx4ExQSWHHzIh6diw7JZEPtrSIt7
WkMIdwzDCBVnB5GXRKTiIP0zd6QjWoIywg2z2qH7q4F84gRYkmMO/Yv/85wLRG50tX8ete6jlao7
jwVXtJ6J5VJEOtO1wbnDHtUFXELdO22y3wtFi8e6Si+WvvmnwVO/l2FzKSAx5rmskU0hRK/mTOdG
RF9BulHsvGPuotkX70b7NzvoohL6aTEoEcx2SPrTUjCwxtT0UCYq1zwuxkWYfS87k7W42kFcVpre
Wu2GrOo1dx54r49W1FwdUXg2/CycP9PCOhwQnT65fbFCuAGMjvs38yCIgzlPbP3xh1B5ViN0QCWA
OOJWI5nl+kvARZW2piKugu/zLxkHnfxk2jYR8tJkNfFW5H/divEb4i+8TI/vp6FEvAtUbb3CTA7L
vbRhA9mTmlGxAhxqAlBD52aPN+TXldIlch0uVFIZUgHcEYDFzLBZjVCwsHX1UcB6icHzFEZWxBe8
hKLp1cZTWcT2ynLMxLWTTpymbrNBbMI5uRj3UIPNsheUNfA6vwz5RQ5WUzLcXl+Tw55FG9KFYkLc
a1hPZFNUdon9xMNZcAxAEyLJ2gzOJY978/6QUzhkN5DpZ1Pyfq0TAW7FttYn3cSD7wQLteKo4acl
FyrumS47aAgcpNwcm4H96R/oJdhw9FHfSYRois2kex7ej/YbRF7mIafVULqWHMyqXkblwuHhOZIm
j1esNKCNyLaIriUHa8OdiyTVkfXOgC7hWfVqfxlfOGZySVo/3tMwa5uH0oL9xNhISXPzO3Ja/Grf
cNj3zLr//ztTnJBdhW+OzP/Hu/vz9r0occ97dKzGlxLq0JFbYmQI0fIlwHZekQvKGVZb1xDlQC5J
8LVzniM5bRFnGU7J07p6IJRPQ9wN0CCRydvi7Ou4y+yiy+pKI4W1hYgezqoPq4CEjZfX7purY0qR
kl7+wK9g4xOm6ECmHDAyQd7NhpjgrG+JoezdwaFDBFU7KheN6KIUgc+Ui5eCvcV19ISsKdKdzR4+
A/Faiz4iF+fZe7t//fGxyDowRFL5JHS0T4/YhZptQrPh5SR7JQvGuq+HfvawbyvmnpgIfzIV1Zrp
iN6buMb+IIuipdM0xdhTZGOLCTWy2ARnIN5UkVE9TUKam0xncQtZNaSLFWxFSV1mQxKBPm8sFjlb
8IxEhJEMRkdj4fDmXODDCRaHXp5kThwWEvGx6G9JOXx6sXdi0j4RNU24YiXY4RYXWjKNev7znKG2
NgU0AG2X94bDITqoiLK/VIoCn5YwvcZcQJMmPUDoFi/49ibCzb+LTCoqiRF7o0kEla5FFKyJzkVX
+3bZpVcWa7E1ftpsXBuKCqRDNHlKDbdotBEMDkQacCLKObqT6I52J/U0qKUJI9cOv40Oku7Do2Kr
cavkktBL8p/kSppMPRJI4QB5Qx3kp9Bf5GEhrfgsjA3uB6y9mOuXQuGXeyTDiQSuvpgjXfxS1cLA
NRWMDSCwAa2Evq+SH4a6+jbOsgcSAstFExVKIIJ1YHV4jFeKsKk9hy08kmygseQup7zW3gqiFo6z
lCr2I5t8qCc7+8Q/QPMZTPX483AuzLrzeFRjHb9kwlsc8DceBJhxyuhQAptAd8pXhXXkmbri+Z5x
ndWJuazEKXXWygU2b9VUdO3+Hsh4RkRAJkg1ZKe2Q+Xambo55RNu6LRGMdUC6Otjo0zsxUzD/SO+
pY7xy8uX0I10AeTa7V2r3oNPQVza5VSJlTSeJL3CG9ZqS6xfxR4bG+0H1RrFGyD4ufPLdZrj70fk
9yE/Htwi0CSoBnQpwtS3ChH5y7h50uEst6AWUOfdlivgsbnytMGI8Cb8d9BupMRT+UaUf6jef6Vk
AdWCf7yS6hRXaGq/hv5TlKNNkqYhwIOzxS7kVGzYwIVh40fKmH3yQJzBru5NsnoyLutxkJCH3vsL
PvDL4fdQzwlmkYxBprbbfCA77CvVyeNHHIY/AHDE+n40pJPB2KoH9o0vlDxyIIM1KPeeBk1ghtOz
qyFkpmCQCLe+UIt8Ww029EbCno6Nl5r9RoBtYJMf9hmhrYiMflQuUqd6zS7Tmig6kmmpddjmgbr4
KfMhFhhHMlCGozew3+1pms89dOL5aG3Ye0G7Ls+pVmF7fx0mvVSMWUAocfUPFsH6vVmZ0l8MvVQ4
rd4QLtcrsMbCfwCwBbj7Vhy/asJ0AFqWwOH/gnOHWyPcbqgbZb5LyaiYgXhfCAtuB0YNCEx1fWbK
BqZMEghGYfeoFChidsDhLPcGlIxqQTXc2saIQoZUd/D0EBBT19Lr9+kKXOR+aWBHcD/OsdonpPQm
ltAv/EqLPi2WQvCICmEtIt1uWV3aSJ4t83wu35upgfRHdtmrRH4A1aaIxkssHzQ9vmsAjp8QpKaR
rWGgl7KnI4MZ3MrNKAJJmabhEALuQv4wDbKF1XbfQ4O1ggS3KtOWdZrE14lklB2BmMIr0qRcXZ5X
E1SB3o6ZgogBCG2cO5AEK8M/VDqmr1H2sglv+ERPg3sSuntCzg9GlLb40pbNyQo4n8+O+d0nnFe8
yhMDvkvciPAr+z88oMnKQ1HnVJ4r7o6XSZKXbA5GRWpc9umuiqjHZn+yltYhlcwNF8EEfkCIwuOa
qSueVaGL/M0UMzimjwUh0S8E4oB2t4iDVSkvaVr4VMkmN/z2a3kB2rdHsaxpzXHa9LlR3g7RY5nO
jxs6dIZ5RpAt/YPz2kWecCQ7vIoejNgdh4JWPs2Kq4CaGbk4kZPszJInRt3mTflLGRJu4PqYANJ/
bgG/u1MVlI8A9Ckfihffp87t2EGYbd39Nf1oQW0u3srg7JqMyyvMu8f5zJMNBwiFgmZRveqUTbAv
ShJvGDnnmkq7jRw5CIGan4c/Hs8Dto3vUytsxW6qJhftpdZs5C3S3fxSSNVa+XYsie1/XldZNubO
d3A968yOljR/vVQy46BG3r2u8hcN1A/QbXIEeNa4VIzgOeQDhk/oJT3TNRS9dFVB9WHiFn7DS9wT
XzIJ8KLDe3SPcPxVtfk/AoK2xXYIF+wtAJpJVWuEzJpEPPtN3t3IV9AXvqa6QkZ+CVY06gmYlmpM
i37S6ZGOj7Ran3k4aOA1FobqPEDgDNSW/Yxm9m70D5BL/jVfKalwGgl3iF4IEUVaisjeXbLZzO1H
4CbI4vcbvYBKUvdoBz64oRwVzFEBH1QB52I6ZKUqYRw6r4qrdKCvDoszTYALHRuDqVOWMGrnLNJf
l5XKtxz+4elDuxu5zRX22COE/Z/jI/dFqzsTVC3ksTTS41aKlzFU1cVuip5dGnZ6Zpv9a4r62tVi
tnPi51Nw7J/PWzKjGYJmoOUp+HJxdL7M5pFXP5U5npBhN8YqDrLzNuY2iCKAl57aqNJuh1YdE13G
hST742d685DHgtDuV1GgbwYaP+7sjBsUK/+Y375yEs0HUBQBk9x14LjO0jxJWqqYsu2v/oR9vdXK
pYjZ5nyrcJoJRnfI7TcHFg/VRedlmz/+eZFHEhRT1L6k9eL08SXEWt6UNwfwIOQkxstplMr8wM5a
Vn19lmE5PNTShV2n6dLPjiJ1ppT7T002wl1szekSqXYTVMXwTCqUP/DfnwIkSl98gEY+uiSCjQVZ
i0ZiTHHR8+c31vYkOWAViJGAG5n6rMhGSOk1ZvmyyrTG1OKPBzY4VLA4NBod0Cu7ttAtN/rsD+pF
2j/5+7r97pAIeEbumdR5u2CDpRXHMSm+aZ0No7lU1FIAOBhfytn3MMLsJJT9aFgyc7Ie2o0NrGhj
eCli4m7xdx6EvnWrverl+zt49K+K78IKpORObDSXz0IO71feHMWiXfXFJkmBfKcLVzWFNZLf3h3U
e7pOGC9ynzuLmQfjGG7TPLXnOR7TyuTJZiDtObmCBVkxHg6XUeX7NoQrNmzOD/qnSkJ8AezpO+yI
XOfI6BlG2zt02uo9JRu33auT05F5npAG6wmFzECRQDGVpXS3SgHVQMtVnN5JSPEioJmnOs2vBllP
UibW85iVu3QxXO1ZT6jHe6E1gnGWM/Zlr3GscjoolrxZhvywNQ1i2iKY7EWXywDBhSLQ1hdszCMv
7T/h0AvIEsLczJ9UObn0tiu9ftNDod06wBrUClL8ON8ac4qpfcM/NAk+Jdu97zk8e/Wl2ThnZWNU
T0vsFUinHJ+kOLV65q9xxbNthyc0QhYbtTaCdDfBif/k9Pa/cjulfVBQMzsf5sn1FqkEOPsgtHpH
HMY963g7bJzjCjZawJ3EF5L8omGchWzWtsZaxQU3LlOnrUDe9gu6QMzTHYDwHJ8dNgJ47tLUx0Ty
AfSqj0zTOQDCxIjPSPvBeVA+Omncp4KB5c95BB5ycYfrOCKypUto9eDm6JproJn+pTO7WbSXgRua
s7gN4p+ZTcYxIdOZoun38y+R+EkvhIF50r3US6k2lvvDvupV6p/RRLaLO+k2kVXR89BYdgTfI24J
Pcn+zT1iX6CbJzkJ5g/ImS7EN0hBlywqhx4TSJocB1UJoHNmddDsp/4y0KPStc4ehKarz7fgNnvf
UcrFZ0NoEox6E7sJv9A43kn7YY4SE+g069816nj2zLQuJd37F78fuiO0O11My/BqqASrV12d4Mey
UXLTSwYRvnKD0KZZ6y75Di475wgCPDjOo7bJqFl0BBCW1jTITdXk5L1XJDlOE9tqo3XB8VMEFnxR
sP/2OGOAGN3vWbTVXJedM6GO9PtOlpMcSSNJs7XYvuEx3skeys0uOogMfdPijQzJhBOEek8k+kuz
yZJl+O38YTXktxMQLGa0LjAqHuPrG1GJFOMX+pY1adHgrj1FnH06n0+g7leDI/MGMO3J0tX639MP
yZodtxcnKq2BTaE9YNt6wszachFQ2cvCLlzvQh7Juo72Qj8i5VEJfO13JLiUMpJUB/j7tMFrmNRX
2ggsek2NQw88EGVmlRDoEeOnb/ZQDsLfHalk1q2FZ40l4N/tWcSTafuPcDsJ5na9viYSx97M+5D0
v7hjMfSVKMDibt6W0CfJrD7UuUmu1C7PrdZQ8VYFC7qdi0FKPBwpYJ0RWEkIqr6PGHpsNpptwF0A
I+lsOVTczKemcu26Tlwbjrg01iTvC0/5CXpVWMyMLUzyNwhBBiplXiFJ+KbExE/uiVbKFYdWQk7A
yAFsti0+4H1On6MQpRUaTHxIOtnQZSVFQJiyORJgKLwM9KD3G7QRZlTkG1MAMPavOVsHU/XrooUD
TuB1wR4f0moKgzUfpl1lgjMZO8alZRmwNYKkYMyorqd0diaArrYZiyxrKvn5Q4VcT8RUGk/UrU0b
qw0o63XORZUG5W1PjA28yigt6FOEkLOhAAad2trvZGdFOkWe5Lsz/R6jgywLNeG7OJGiTgbry6Li
BYki1IKf/mJDWhBZ4JVY8DnC+3/LmveXklNt0Qzygylpsx2ZxFVHb9XXsAy3yVkeWt74UtCwf8Xq
0w/5yvE5pWgvwk//5OYG2mAzrmgXsaLkMV7CBDvxbkkzZ1obwryTRf3glQr9Maqq3vEjQcqyiQ+p
9hRMxue7tW7piiomun3jrxQdsTrCGCQoWh2PIZY5orsMZM6k7hfhsj9Zmm1bCK0TbifoJarT11RX
yIlqt4z5a1UW64hv8N/muEkJ9WOvPGrfErS7YU5TveZHAUDCWDq2+weE8sT9uYvdlddF9IEOTOUO
VOopoQS6S9uSKpNBPWxBBM0VGHP26FCKLABNcg0g5RKL6fUs7AAUFKAhScN9sA/BySdOaYapHIU7
cGiLTOuYXT9tpbI0AQN6RsqUxwEXcf7g2OWhtigRQzK0aF9RT2tzK03PjZTI/zZThZmNnpWC524o
lHEB2cqQicSHuwTZ0x4/m/08z9d6BzqXCi7K0jY0SGgEMYhF+HTn//DK5rgBu5AHli7iGMZKAFXW
5eIKP5Sl5+LWuAIM2SYIV+dercDbCBHsGDerV5TeBBEacxaWXpHLgNcJk10tQsR2E6DWGT0r4zCT
OTZakiX60WD27IHN6skUc4iMNP/2RfAZtfV1HnRNrnaDLxBMK4LO3BWwH4X1NWCZiRZDRK897Qy9
/0jFQcgfJIkIHbImQXCxfmHaqvKlja5S3rjZucfta10TxUb5tZQrVCioWLNF6lfz967yiKAt9BFx
M7TscLlX5EpcIe7oMFVyNQNQZHQnaltILAS0u7dvd6E4SJGwJx85Amf3v40FyuaGBsSIlEYUkBiW
w+rpvu+QJo2Dudrp60407VpYHARsuxb5Ui2dOg6W8jZrcua8lQtyXDgwZWDzMniUM42f65YQKBmS
PvebiADutNoDKd6XpsfdeKnJ+BuhnosTT97h7B3fDnLDNak+IOl5jkKmMhtruIgK85OorqCB5b6J
t+AtPqrUrkcxdfSLXffeNU49LKoGMD2sWrFXtTANyOZtRUPB50FRd9QjLmusVD7GTyrnow9o0n8S
r2pPWU2n3B83WPf+5tBWba8cH+s+pHYy4lTl1r3Qk8Ut/xPEO1mFNpR+UsH+az/g9s0PwFGm2Tnb
DVYoA63zKhBrRH+RroILFZx4GAVwqGwZYFzEnKCHKdbW25iBO3YP4+AVXc6qQyN4GqLHHe551A+Z
JbXepRJw2+j4TZG31nRSg4yr4ajtUiXs0PtLvXTq8Nn3EWPA7A6AoEKYwRu4cat3QHqwavJS7KWI
0LENfpy1ldfi6wKcX4S47QVPpQUalnPuQxx6i0OAa3ctRh0BrrZ9Y+ReYHprW5Ksle6ougmOGoYR
bz2QJab0iXKT3et5LTmCWNdNd/l5T/1xQH2+GKZEDeEwppb59NrkADLInudng8MzN/Z+HL2g6eAa
cjvUT6T5JRH24K2JAtlmyQc1SgbtaUaR+ZcxqElNv5E61IV7Gsi8cd96HWX9sNjJIILgxZ8c8Jah
jVGCbSJbZo+Z4NIWYLwhPY4phJ3OismUAhoyLEmA2ncIxio2yS7mckIVp6XRIFOdjZpFoTiqCs1y
XvAsj5EQIOhBUfqOnfIs1gI0Q/cESLNjJPDsA6lNvzkbYayTUrF766AHmho9MYDJFus/c84SCjj4
Ah0WbhdWgRf/3cjlQccTuVxNVRur5KJ7HzfyOxiBjZN/0bafbdLDZJE6b3KxAXBcM0qCopegQ5ec
yKNmqEYfxftOXGQ+FsGnLBhmlAOcWD/NMbh5JozHkv3bzqswy4D12EWRGBgchkBfrG5ONgwGqjfz
qa+kF2CIF34hsteoCfa1/86EYPmsyappqkXflU315FthfAg3fNoIiBMsEbH1tL0uiXIYc9e+Q7TV
TjnV1/yAKLLnQM3EhD6bGaKGjRDag10tAP44VOCnOSgWcjCe5L3M0z5UjYmgNsQteXKmjJ2ZRUBk
Kla8zn8dWnWb5lsVmpKN08t3bThjywFiqfzlQ+660Re9T4L7zmgu6XagTJj4D5AYnu3PTghTI9bX
jVmh4J9Em+rJGknvCauVgOnZcdToXkIpw8z3mqaIVbKH1dM/8oAzELUuJJZpLgAqaBQIG7cB01sS
mwUV2ZCH/xfz6Albh/uRmejNISgp2HpJ3C/try9qv9+vpxtt2maXETVbgXLo8EF1a7NXAnGLBx+r
M4KZutrzxHsHbut1hK5VzKUqSCNQaSWw4sYUKZYYJxNHCpQal3UghFOCsaYjnuMPAmdDhQlZ65tX
mXGa9+VouKwuiXwukpJm52UfCFM9rSS2yd5fR+Se8atMAGLUP/qVLlXVfHzE0IjOgggeqA0Ns10j
sQnHB53gHtymyrlJvq3wPPrEO/1MEeeTK16sjeqlgPLzusVeKlNJ0znsp0g8Pyx4qX2+JHthe1Hr
3OBehwln5z/nRN9W6rg7e5JHjvi3laAnrKJhAtA27LCm2uoRlgVQFZdYa5/z6s+zmqJ28DRM3bRI
JZm2+SEUp2e4vxAEf/SRdJBSvk/l1adsSoIiUz6ulcmWNg8lJ18zUJy0ZRZV7YdJmn2YdOejq3jS
s6SfWtlFeNiOE6K8gQg6ML9zUDgqfE7k8fZDfnRdzd8aqFX4mYxeTvNpPyFmPugwDOLSKQePUDhE
JpG07sa33RPLgpUn8G5J6FXKqh5wZuNX4DL0wYxbQto41NlbfGw5j9WgvYVF1TZ1eCG/F2XV66MQ
9soZceEBeyRFLWj0TBWyXC+Ty9fsxcCVrVZmZ/zxAmxSFy0N+kJk935cQuAEFyx8YDLpMFYXlvlr
6WWCuHnc6r6K0HQpCEAAA6OzJ3/oBrKE5VNbS60TM3LnNq7pi2f4QJ8flzoWVZcWkI6XOXMjkvr2
O5wVUWdli1K9tum63ykSk9ieP/C5DeAFEXxz7drWdlH8M/c0FlH5A/QmoXbVoYJ5vSZvy7FnS9jU
hgXvAEmTd8KOulQ/VhBW6k7CzdfNUpH+ktcU+B9AAGsjdKeStUj/vmIEQsCAl6r8x233hkX0tJFT
v4jW6g9zp0IETcptKo+NyY9LX3yVs9SOWRh5Gjc/vQ/C7WCEXHixWZ6+aj8AFqVtnj+yD/Vwianr
1zEnxIzAOrSZDgPDgT13T2RgVqR8ZtirI2NQp3J29z9JDHWpF2HQFLAuGxWkikOybX6lkJQZphdC
YX1eJltofeVfZwE6EQm9EcV0U2qX59z9+ubYrnfaqvYprk9EJFyJA5/+aSY/Cb4gcWrmHODUkXjw
U6xvoucVF7d/Ucia07rD04pL3I9LtDcqyPvcxbBjnqDz/GENZPDsHLFCw3cXI4hbosKZ/wHyAr3A
QIgIS7sXaYvXdvTOHxukQmoiymP/OF+93l9jZHxpdngyT4pZ81sQfhPE83rDbJ0Ikbv8AeiLpJp5
tc59fti6KS5AuEfU37V2fvkmLwPKf0M71Z2xuoRbc0BMs59PcPLhNabExsz/XDNviCFnD3QgNhhk
RYW4XUpQUTsrGqfJEm6Tn8V3rexVeD2ufqJetmJsKNggyjNy9K5RQ6VT/wp0SvoLB8aMnxrmbLRb
HFgtyaaxJFAvurUV3G9oekIPwYlnlsKFG2HHkHmO5ut0chaqMvAT2lj3UEQrQ/issCTW8cNl9q0C
We40eh4rJOHKw9n0DngTV8OJLVXBh3Co5DfXg3hNlMezMgc4lJ3bkTTSXmopDhE6JBTRd/UVIqqy
pAcjE0KXuDFhFXxI0NcanGWMoKKKarockQhCVQkls/YLq1OmhfTw3S5f8KI1gZK4rH+fRsADIpK3
v1MzisWpmh/n9jFG5zXO9T26DnOWdcUaODsPlIZtOhsfLrBCYOmuqTVNB0YsjBWxb/UYC8j8KgEG
k4I6rYt28sZi96+KksAiTdKMWyXRi8Glo71h9787RLLm8s95c1kWDRuB6a2wgAs4nmORgS6HwB6t
9cljAP3rQLTqVEZzFBgayUMVmIUzSxnjZT5ieVkZY/mGc0efLbONoUgQ8EgShmuAcfkse6NiINoL
O0TIm1PjhL817pgqSeb45jWpmn/ILYoXThdCixLRyT5z/8KqgodbYMTKDOmxMIu+9BMrmlnx+Fst
csFGiHTz59ZMBYrgcnScI2YWCdYkponSuXHx9HQk7XkIAZhlHxJ2XvxCSw3DepibOkNCFZQURCOk
Scnk9zfnZOqCYAH66GG03Gb8gi3nSgAmXsL1Uk4Hw7VCvHHXbSTYYPVCCOxwgYJy9heYSnOixX4s
xj2oJ7VzYaEjt8b2zqbINFgVjbBeoZmScZTN9uharIMcmjOHmI5v/owo9ABj9jff8WLK6o8BNN5Q
eN8DPwBCu9WPvr3bi+mu13fgD2A3gj3aFodpKx+C5SEkQ/+jwkpkBhqOMGZjo155dbgNDuFPOwAo
gQMvxQpAN/A4dgOvELlxjGcLOX+bPP285r4lJtll+FGH7lkXsySNR4qwGJfrADBleGQJ+qg9Ig7C
3MzQvjgC9dVL3NwAXvCpBBZqzbo+qM05emL1m8f8TXgMyk4sozQQEQskaI5k51ESmOf+maNWROic
BJ9RF45X055qM/f4X+6icd8ldcnPbVCdLtcVVsZ4+TPj8CKamA13z6U6t/RdomM3ftzn7t6zLP72
VMdCvXVCRtgHij2FsSZIzGGzp4D++KCd84yqpZTHStgZBWlYJNCV6BfYmstep0uVbN6zybuiOONU
AgS/lMA5xxX2oIjIwiuQtUP7oW4dESXoGgGO/KFBDvJnw+iLFFl8f430PneDMDk6Fm2mknueIin0
FMvnM6qCB4GEJVc2sc1+nCULYFV6/uyp1TYlRLaRPi+HMKZVEcKyTVMl3tck4TXo/XVHe1aWK+er
iw8N7iPT7+1ky3g6Jt5kRspAzvtNF6bBhhdrbzF3chaucBhpCuDOQjePL529wV6q/eE/dO0LrmUC
HrFeYQ68E3wscG4/mK2AhhaUmmPmxUSfzfotI+KEU9numOnrQNeCx8C9CWbKjOYeulorFE3yCT5F
vdlO088v0d8p6XnfM71iu7VB140se8QCEulwxizKp5IhG4riymjx/xK3XsWb1ciFOPhFBHVcMXSW
FbakzkSCvOr11lTKwioSlg8tusQiPab2lCryYI1qORcH54FYUYHifA1urG1KVPCZ+UuZFneS7t+Q
CLCYtpNVJOufyVxJBxtpm6qdhpqpDk4Q4TgNl6efl9SS9l2JkoRB/9M2j4f0oRK56SVD5BIbyFYM
8pOzi04fYWbzPZ0wE9MpTZun85bjpXSIEoj06rl1h1IXYe9kTMXmUhOZ0N//heZbjsk2v8tox1gH
wKj73CQXhf78uW7SJemscDHAa48WPixvLp76Nup+dVui2mJQ05YuvGzmCotUg+vxn+1ovvGm5tkL
xnMClwtJEJ41dXzwXU4A3AyLloxV4WLGBrZIOPje6NHGkDLLU1T+h691MIIMue7PPGr1M0FW8xuS
+Hl7n/us2HAq/MsGJOCSYFs6PwK/1jZ4bgtpAQHswvhJjit+5llgDI0mCR0tu5obx+37xhbevzJe
Nyzh0jYXuEQlmNnPvyOKsN9aymlZO+a2ZtY7+Meyi9fuThcKo2fCsy/OUVP5SmTT7vvE6i2Y6Q1G
m37S4JsYLRwUm6CeT3DeBNMQRp+Tdov0Pv5ZiAffp86J6tDfyKoXnyfr/4gkNth0u/xo3MOgYK12
Gl6PfcZClZtjPRsuFDbFqC3rnIFDTWRTZqoCwzXVTNiBynLduadwpy5lg92EdbYoIVtyltsgLJjA
X6cjZ/Q+TAyvbt2SKdekYhQMTfCR0dEpFHZBiwY5Dgw/BMLHlmyn1IVEVsv8Je4RRRNEH2TiG74F
LVFDZGFskYqCxPg0K5aXJFimKGw2Ix9xIDgybvfL6qWjltGy90n6VG1Wx4g5aw+RDIDsho8GhctR
+uZkWpe6PoU+QZ3gYKKzEdIgkFxhixxOcXC9SIw60WatLK01z5iPQypGPS9AS9b8Bpj24yg8eJ25
vgK+CrP/wPIg0kipgluERCtUGJ2IVyJaYnZ6IpU7YaysODQWx+OlEIAVZFKkn1gEvxwz7aG6JLKP
2lw8Vd5fuma+WgrrIeRP/zQYkvuzS6cKlNOiOhALa4F/GJ2HepK2/czJ0s8GFvNWsjoIfEdSUet0
Bl661QKZlENlRvOR8C/CCfpy5w6DIa/wBdFCAeFdxySWq4XRvK8E+HZpOnZMt5IFpD08wXbHRskk
29j8vb8QsXd3jWqw46LeKmu4gqNjZGPfKgQ+p9i35fexKQP9uqromz8mh7qZTJahh76zEG+aCFkk
lImwomHfMthRzvWqBHF1+fdX1JVe6rAVL2MFraAqFgowqyOlKxRA6zpHGEBQm3pCfns+FA1GnaMs
h6RYGA3Z7iQLocpJuugDkfWQRhCF91GitDnbWioxn5HUapVCKrFwpIFWMZZA/P93qACSHyHEuxBI
CL0XxGU77t3cSziMwhiCAkHWSGD/9c4NvskkzHVeKX/pShpJ8Vi3G5gTKxlv0a1/aCv9G1gRjNjN
UoX4VmLx3OSiw1JEq7YEGectY8MtAsUnua4YiF6j1ioAclmIdcFQDIcwlIcsP3SE9zGt66NAt3AI
xR0x9Wn5wBvL7syQLoBydMKHOsqyAVUoWN+TwpJ26WdhOhSM7qwKlexnrpA1QnIoAF4C2p2WDClZ
e9BoHkHuIbR7xiki9scVa4o8gIEVIJA9+0vS1xOyCqmrxCuaegzVzA4ygoKgYrggH9MPgOWsYbOT
KiuccZj70iZztZ6l5ywbKv09gN5vlHvTiQonBVFDBAtAmovghEhlqvZQltW/bworQUY4UsT776+G
6K3hkdNZyjJEvXXeukiBS8Gufg0S532718+oORb5tB7nXuvuVpN7qZkCqhxS+9rGiBDrhQj6/m6Q
TknXciUAl8Bd8F1FLMpJPVjNnhfss86IaUarSvFxVYtDQoOsUE2BxX64h+Iu3uUdVm83M9AjJIuc
xRdSDHY31GPvCQUFtgGsDcNmAkaTMLhVyH4K2N9i4Gv/NUULzFqZ0WpNoAH0FvQETGXu65qDfdF6
qeD284EWQYG0pHbSCuvyLjjLnFgyf/P0H0ho5Eq42eNKxnJtFF3EsLyj7m9y8/Zd7uLiXGRugEIR
VLlcxS6mI2M8dRDTu8buHo2eVfzLo1NJQaegpykdaMnPrAJbDGW2CSNjmMX9ZmEbNLeZHO4EG7yp
W3Kf0wMX2i928utHnYu6G5htu07QdbnEzSE3NmEQ8NZhlenPubWakZ1YH3ImKU0zvuv0o77e6baB
YEIeBt08HZUfNC8JbzkMPQRHM83ADzCySSi5PGOiiYRXDFHGXoHmSDWWKJJuwryVkL4/1w6BB1SR
+qR2SJvzqn2Q+R0fWvEYO1ZrPBr7Q9iN/NjZ/n5mCrVBSj+HXxwldM1AMPsv2ZiqRTdjo4A7k5tB
wiON0Qx/z4BR3+5mlFGTOMo44GWWv/hJMSAGcKdzDX27jfTaK+/E6oWCR7vQvieF7CrroF/X7ztm
cDtNYaim7PhWD2gDRcg5ryENEem0t5EXHJOxLWy/iHKaZOYfMGvXLKlVXoiDLIVer+8NQOzkXGuu
j5UtpcXhMy1YEAGL6ClKY+86bQTsja+GfisiYFveRsDFS9YrvEkeryCOFg3uw064YeL8b0lZ7tgX
EdE+NioHsPsX8NE+yoEVAJfcJP5ZwVB9vcUWMQ/8B+XMJNcpGer+j+3kJS77SdFnAOJS/BfBGqZC
1YljgVvl8iDpbsNkFF0zR1sGCjn/mhFWsV8Pf+ofiQn9xfz2jL7VFtxV4ZlmvZRjWm4G+jP6NegH
ES+R9e4PEM6/Sv95cN3h/SQRdB9TlCLj0IC08MTq3902AQeNPCpUfu4suG+VgmI4L0CrDPxxKdNm
+Ar5LeJU1XXKP164Ir8uh+CLLXZ6q+SBidZVgYjHG/QWz5M+cDGKVFmn5V+QWUej975mZvpM2bmE
7/xYKsdkfQhxcD8rInk/pK2ppEYXKrQd7Wd+DGJwfXQjWNPKjf6Gwv7gM/TzKonlly1OgeB3j7n9
caXO5XipRl6mpxGaEWKnl9e8AYT+vWvhkTCWH599tJp6mFihz9+QXXkvoEL/++lm7BiHE3Qwz3vQ
BXUy2GGeKCOKjXys48ZHrkD7BJzxwMgBXDUJhaqmhCizrgKlE0lNw5g2OyvQvekWoGzyc9BT1A90
j7lyemecjpDRsAZVQLatii1fy8wwH3Cn5MlPMAK5gxhvpzc7zT3qKkU17NyT5QmM+xN3QC0gW1IO
dzN92lFKfi1/RxLaheWAmmzEpYKNA97Q2yldiBDb1ShR9opyZMkdJd1pQbC/qOhhjbOO+p0/8tgv
hy1+qO85MZe06Wq8gsYgiuSyTXD05XgGpzamhRYKBIoca2w/yODgH/gFoZqYhvtWIwPJNdoD0VRT
Eut8UDZ0pVKx7OkiAiGljbcyJOXpztwIrBC+7x/f9ZHxv/6SfF8yK9jQy+VId9cC2k935wyASK+v
viPHvkwyfYA/HFH2MVOOpZKh9u9t6/Bo6O0LQG5nHYnr2TQSsBVb7MRLWozgVrchB4gON8uA9QwF
JEkim0nOeLHuIOkdO/r1CJ1xjzYTSU+4HTIYVewr8o9KNUVZk6nYt5bvqGkF8DrVJJ6CZNKdl7jK
yhR+fpuIMwg0w2f0rWm8jJYgyYVmYDKndgSgsv6zONtJZbFImAXwHR6oTUzWOCUGGOi3OHvBBnNz
x/uMlFGunXpGAM+EZGfPYEhnMIlBp1zMvmR8XLuAxykrnENIV4D+1YxR5YQvTwCpE5The7p1ZjFV
qEKgzWDAynehufDXS1APzIpB8BFaiNQrnrkffl0FxnhHEi/C/qw2hmmXgzLdf6UWLMgvoKWenhSn
HstMUi9gfdbzW6VLoCXu9QQ+h9MXGClhixUfoxzOhdg8dooXnuTPHcScS9cX/pobniaZgwXpzTYC
NrcovkFC0lYF6D4jfXvtUwYxtHWacFoIwOeIhYemp4Dnk7lp0ZMo4VyxVCEYT+UEgBA8Nadqxu9q
9YjlvYB/+jBh4XjQFEQFkqwrVdfQS+1I/Y1sx7m1e42UwQS2S1x5IWDqp/4DzP4CoZTObSYzEnyH
EHrtYibgYxpl1/2uc7iEMc8ruUWkUrtHyyeXIu0uF/R/ehM31mnuX2u9fNQZjAIHGcqFN+u6iOkh
+0tTcQq6t2vG2DNyGygTUbQ9YyMbbmeHApIHVIdv2hsVKWnTo3yN25k8qc9JYrCPEADfo3JWubOq
49rnkkWFpMIXRmZpjPdhSStyC71tg7MQkvDSSoZLCVj0Pw1Q6yjMKUzlvBVUJTWqD+AKUsD+FKB+
A+92AiEw3cMLa6YinK/qBBRV4iJ0xmBCxh9aTpmRYRX5J6d6jrt/rAlrF8EuUiUPtGjFOobvLokq
HgTWcD9BMY8L5ZiCuWPgrLi86WaGa6sRFwMumNSqLW8eble0SZOnp+JJaOFbEI2FNgPQc49zPP0L
WG+QiWifj8IEAMf4epD6Zl+QOA3d3VU5C3N+LKRCqBM6yL7DG5kQSru54X270mpJhzkQvcEMkgMi
LsnuBvwgTn38ufkWBBMgiD0GqFLUH+OynPcwzHWGGjbpH1KCCOsvPKOWBL3PJm+agh/uIfs0BaCr
4NPhaTK19XI94Va1bET9BB4Cz9JN4FIJ4q/uGk4ZimMpsxXdS2gRgdJQ/nX4Fn2azYtS2WDOrjjM
awglJxONC1QV3jGSqm3HzGN7ZiukNpF1t0OaCiO9Z/HR9RR3YdmZ3OvcbRnnL++z0jpi14IM1lz5
cNxa/SH4dKiTy+N/2QGPhaueeA22aqSYf2i14tGOqzy1N45s5VKH+JeKRIHD3xEer5yCr3vpfWL3
ugFH9qLuWrX4xrhtwUvHH3cwRrjACHSf7f8KCIZkUQPHmmutEhrBGmRoTcbYA13STimx1qAvbzkX
BiV4ENCfNZyYdSFVHtDs1++UVbK4NkezSiXX1+HpRBe5HWGKd88sfT0cmAagAX7pm9feKRpABCDf
xv+zqpnYjuRBy4SQXKflEH/lBHKF3pYFfSLh2+EIYM9AdckK17kiCTstrUuGx07VVS12x/N60UlV
zwrBOKMEHK30k2CmjbiPFlTQk7YB4zoxE56Rja6novw4lZ2vHRRCOonft8mHn/icMNlQr572jjaU
qgvKr8hJV8Nr80KwKtfuva5bCtQ1l7qmceWxbVC5pfjXOVcFAy3iQehM0FKcXcvrLTp3GiaE0bMT
/eu4/xUR4OEWywJgM694GIWQi8g+nFgAaaDhjX2I/3o7D6xPZnUYXnx5d5mqk7u2yGY6WzaVbZGX
olHgVsTe1PL9u2NQvg2hSo8frJbzkK+5CO0w0zGbeOBd3PCHQmL890CeFJ/3YWo/kmoNboImB5Wb
i78pKWhQ2nJ8QFf9cYxsMghYdStMzHDVuhLnNuBP2xRptc25JEcLaTofmgPcoAhPWh6kTWa0Qd/6
NaW6c/EmI428uEQHsUoFjATMIyZdoug5s4Jb8dWG4qCfb1cT3RgcQMfIRBQKQI47H6OQ1uS9tHwQ
uLYBHGNjEI+V88Ch5TTLE+VphNItUBpz5m1/Ac+6RMLwLf1rhvX+hw2Y8CbeQaMnlerjlXDEfnIc
oKhhvics9S0dXu9X4+M+wjFnhewDVvj1ZmVVXRLXTTbx37NGWGXd1lfY3T/LviS9aX4+Nb02Zamn
Yl17CwWwbS9fi3w5XMt5osQ8kMSiIS6p6ZeM7x8iJ6u01fM+WFhKbOVcggb2s2tsnUTnoaphJxv2
6BCYhsahJWwkyI5VSNVmg3HZy4KK/JzQAOgkse8CH4lDksml4Csrv7gnozpzChJKTS/6Ro+CDe6e
UL0C7kran3mYoINB4Kj98wPwucW53OFv4ZSXuEIFbOIW5uDMref3StNQrsORn5IMIMMkzD53zijt
CC3Gy9Ajfk8Y1Skiz3TfS78pKhsGq+aBSAgTuiJDwmGpn4s4gT+2J5RnlQV29nyubkZ82u7npUem
4WXZXFNY/nDyK9s1Gm+DqfDBg98L+lNPUh6KsO98xjbu188YXpoJxItVXOwyiOsFSn1f3SrdfJOv
clmZV1wExuCxplBxHfzpOoTWH/rthyYunYcv6x/bO6HVIBZeW63VEdNZlTRZm5IUOdNFgaD92BsC
kQeKC2/KeRvayQRF2E00FfAnG2YbbyfAXjGOWM/8TgESzGaZ47FOqYdIEprhCcDKoZkiA9vOKfZS
GD2T4AqLMVb65F0EMQILqzAqjQ5BcGtchkQUyoKkQPelAo6SWGuyxtcgGWLw8xB7UTzz8PeC5UD7
YbkXylDOUIGtGPtUavXnwoQ8kThmx0GazzeswyD3xcLVjuweZKmhxB2oRQQ4dfS0cL/2mTh1r2CA
43lzJeieGAHeFgSP7l6KADrLEQXSqlPFhR9s5nPqAMoLxtWofM125mf5DrGg1/zASdp/RuKTKyLA
Bpz4Qhifk0N/blHwQ/KMjxFUKnXVmJ//L8/w6f4A4fsmpgjYcftdtwQlZu80ibRAfAUJcuLwmF8k
FpismKgtB2J1ijJ26U6MdPWRHcS+CokjCj01ALii2pm13qZVgcRSeK8fJhhhCFtvNMEMIewQ/p5L
DAR7Vh2sBpMH8CM2itf32W8wXPV0L91l+mfy/2yHT9BjunR2w6NVuKf2o0vnIlkZ03xWCFmunaX8
NhYgBXr4gIStiI5RP/T/NrvosayvdM9f67VMl18wimedkDC4kK8wDrwN9rDy3LuRx+lfRFa6TwyA
4TPRzWdscVVijH3cRVGSqo6FtfwH5myzEhDkBTwXsrpJ0SZgIZrBQUWc48Csh/XSE22MmjNRNmNX
xq909t6FtF5HmSPJmtniFxcTNctCOmcmVqJGqczVHtnSYFnrmasRVL1TTKXuC6DFS2vKvAKQcgD0
e20RPJvMcRHyMIYvcjLKu1c7TkjndgN2reEBKptjF435pc1qqKEwEAycmtnOlV5Ger+BojqDa0vu
IvWZHocooniOSCplHKhfFBcwOddmEptG4LHxUze02mNEqKv3UVKdZS+vzcfkcH4WMVsYt0eZPs6g
o8qA7HL547ZV2Ky2adciKnOq+azHEljeXtfi/VdUdAfdvR3irBzZlioxjF5HkYcCzlYEZEI+qA5t
KJ+uKaAdYGpbSOtKUyBBsYtK6BimfwCuophdTot1EEbNicNWOrRcGjcztHFumjK5AKeLd3SkbGDT
hEpuVzWfhGlCpMehu0eY0JXxz/RpduTa3VCM4Yk73IeYRgSv5JB3KgLfloVnU3a/bkwDGKXawKnv
CppGwqlpronxcerng1pbJK2jbynN7Z7xWRMKyL4JIzKBbdUUwxXXb66+QTSW6T3zwXErqsJlVgkw
eHZksfut6/9VKF8M12G0s4GQtmPIVmfZz6IiFGq51gpf+bj3d2uTzKiXfoep2pXmcnUwYcvd+1RG
GhPI/ykiAizfbdesJKLV8tbttvifwR7SZqn7XaraDT87q61BxQVDUXk+hKzNFvLRildEm6DPs6Ld
BWYJ31vwBYHf+2cZM1vzXse7X3wlpQhKgQm9tqovhfFfG/4vmLWdZnQ0pXwxQVZ3TPyYKAQ2wL1f
IbuPS3zt+F21ZogPzNZzYA59D8xDJ6Y1nS8Cem+hCw+aO9pe3WH13da5KT4iTylNBo15zqmzBZnx
52t/yNz2PN6XCKNTq4fzUQ/d/GYHV8rv3uBb2XLScgf1aIrJsqUz9HL2qEjXS7B7dT6+XL7zc23x
srKH9IVo4ppr89dXEvl87arxrfEnUStxzwF6rAq2mqDXbebYxy2qaQAozPWTAAZDxnivUs3DTVRX
Fd4UPhcuCAubSRiX1peza3rURtcW1ak/uhyflYj/saeUAr7AVysH59NklINfyIQfIPbXZ5nIFTfG
k+lQtQvayMxFfnXmbzUpnbF1HAed5M/uXWfk2UjbS798GVxCCviP8fx19Rpem/gPY/2hzCEkGMqs
t9WTS4aUFvQRmiWaXNYaJ+BtdWmgkd0oyoSiRQJgeNTUOo1h8vW27qtw8MemNo2LzBcqU+4fMbOm
tPwK1QVsyCHKnJWosH8OEMOV1W/bO9MoDSfct12znNVXvgDZmmpt2mOayl2x8itwGBHCckCWtTQH
liyEEC8BlyJlzHlTve6ndpEo6V6aiGVN5lwBzm9jin7EJnTbs5dKqFz3swIJJDFP4CSKznHc+uUc
wEeBWyDczFafQ2cS0aPhF+azZP4bQnb7traKQ/X7EVZY+p1kGXKANcvh1kjLovy2FiDWkoYDjzQJ
fk6fjTjWPkZDypED0DwmvMpyoHup6LDXeEAK3KFIPQMKp6OwwIZkj7/y1+ykqiktXGH3JNiWFbAq
wpwRyD8nbaMxkEeaJYxXzaCzQUPmcf0bQIox3wa2LdWxrQyV9Y+1RX3sQiMgqLjbQRGgtdJZNuHm
s8BWsleCgBuqTj/Jcs1ai41P4JyLGIvBFoR3nIJJx3Vm3yeX/DZSZ/HjLocIrhaHyk+fIzmbTUHu
eHW2TU3ZGOU9DcrTTDW98lsrN6quK+eCLbIzG+YfsinZ7DhcwzZpH36IPNVdxGCS9+8pFb2TTrym
eHQaaRhYejvxyiluTI1ksdodsxZrYl4XWFl1I1BUOlj6X30QNxJccqCG1v6WacrbSB3fPlf3Hxji
yx4Lt0PqN4arS5rW14ZdE3O+fgtu0Dr74PQXBsQkcOeQWRYHcvSPx2OgMFO0qGFq0UBsCraQvDxW
fBDR1ORu8GnSJIWZFNJ4HZoosd9aBh1jVWZ2pRJH50D2YXP/2mevxcWapw3t/LyDN8ryW5MZlz8Y
OF2F1mqQ908FbQFC3uvPYTl8PjukJtQgVKDZRUxoEE34CTV64KwfDbi+ovmSH0NJzuNJza6UUpMn
HB6Jrfw2soUnBuF7r8KCTLkGeUVyeVJUwA09GEBjN/H7FcDQ6Pr7xdB9xoCKBqt9iFerQ73HJCEI
J8JNGUy/yn72Z1bGzcH5Prx+VLuZWtg3hcwDxFgnxetmE8OxIE8P8YLpHDXN2PizAmDPLZVl0bKE
RP5J7QdZwHlVzFuCp9GJ6TuJ9yeqJSuPaMgYdLT0MDj5xar53JmlLRoEJiSJoabB6kg8scExYd7y
zAuqM81wK4gqxZ9DOEurW30anZpQJAPYHlGhdtmzv2vKRIpqY9do/ZJ5A3rjs1eMDypqounFE71H
F2vicA5WnDSwA2M4RK2kfka15XnvC0csDX3+lTeqmZV44Voe8y0yyRRkUSCH7VT9jEY5df1BRcsc
xseknJ0UEk7C2HYvFvurL/9GbwUwFkJtBiPxtXogf3KJj5lY13qoXwI6fDWBZRgVKdHVl0H3LliX
Mu2yBfzYLoMRZLpcT2FubmJnTTSgIjV+B8i2yldqwvw9cTwhBiLMAZ3uJK0m/pgewLlr4N11UgTl
hNWOkpxDdOafM3v97b/4EEPbU19dSxzuFQ0p025AtMYSLCOi1lKcR/hCn8ElPn1wS+ntC/54G8Ct
rpx3eFBm6UfHFCHSqugHOklucOz2xEVyG2b1OwJD2RO+5v2wOTa4tN5BjOwUmUPGXxEALcrD19uz
63BW3DA1n/chJmSwy6Q56cPX52yXDhkFubBxIqMlezU0+R05eOaLptkzSRtySmzVW3icrgJkRikO
kKGTCcSo8lSoUkm2hwDb2CvhhF7OQk1sTRHMf22NvzlTyTPOJcHpi1P1DuNWq+2jttP00qCZhKck
fGqtFGeLLyVmtMLSwsEf+BLjVgCppIIAK9pbtyvbFBqxR83KrS/gHqKnLBXyNTru/CORgoM3PPra
TvvPckHRdsFTYjylzeO0ygwbW9fEHRjsffKGSYbjuN4TQgvnykGeqvveyEjwgfaqDyA2+d+7BZB9
IRx8RrpvoXB0Qgik0D3EIC45nFrf7pwpbi8XSFo2xzlHysk1PM3XDUsCOzYxe38ggytiZikNhYUA
Tp9t2G6mSs1i/2+Um1cl4LTHtvinFGONJqParamG7iMIYsRDnVgvOz3LP87W1xb7UdqE0JAY8irC
hprtm/Rn1yYBXTcfw5mULXMecCbPUUqK4s3ZJkgj5ts9PSQL0+9k7QqWnPSNR1na1pd4mBL5WFoD
vSt5lHOGk584to+7L2vTn3jHysOTUEeKvte4+GY9yWNlbyMA46F6ld0cS9++TpJkf/vM8iaI7Mxj
Y+f+7E3r3FoqN57ZOSvqAnrdErcaAzAZzGIhppouyhvs7Cu9+8iqIbnhkcW+lWdkXLwZAmNnNix5
NvyXliDGw1jbihpBDG8Ww8+9InBJa4NlpxGpRp+Mp4bCsmxKg1godltZH88axvzPVs+WbyT61Aqp
QswrpSlsNAf6NNUBAKGaKv4RPq9jw6AXrs4DS0T/2Ffz3BcpdLH4plh8SOGr90sue1d5wKkWHhUY
WQWeZOIUFzEsRehnUT+JMu9RZBIrgtJJtgPDf2XOsEbHXm+qj9jjg2FCsYwJQsjpXkdaWkrFORq8
6BReAeT8yEma2yKzQbYPsQOzk98bQTkbRRWRqZBNXJgJDbuHLzAwO9PjgAIVEEogAaMjI3KTal+p
6tTOqDp/TV2jvDTBYw1J0zjdMS9yHafhkgR2f4eo5TIuZXgchjXkvfmAEgjsBeCBWYi9ago0jZA7
cmO4qV4yBdsAYA0O5ZJY6kOLDw66zNOM4cCwOj0CQHyOp29J26bIm9TkJVSzE8N/MHfOf67yHpfk
4NN1Aa/U5M+se3VDvIBaWIpzbvTniM2pLHmU7EbUbAmXJSfJdU2xQaubFcpwC+Z7UgufQv+o2ult
HOg+lZ2IF7bKzpCJhVwKxC/zG0evvXMW1gqgRLhvGxUWWIHwo65IbDYhliqPouPbGqy220VLeu39
FYYHu5kBUHhMJXByeRVjB5yb3UVaJWRiPJNAbq0UmqnNt/7yum4E2m3IL+GMwVjrKzaL+DvMiuyN
T5NuwpJilbeWHtwdb9dflOw97LDqTVjSAHPKX3rSewLXT13vcQTbUavyQH9B5gqRYXk3i0cwBJBK
wGx5C7f+FpARY8lLUcy2rsK5cm73T0udSaMORQYZZvULlLp4tBbiIq6BPASD/xEdM6+K/hJ2tQDa
FucvlQ0IBtiL+w5eZw/NHgqAaoxZ3R/tjip7kI4kkpnLU/Ph2zHIjGZUOdX44jzyNEjpZ7g0E8g7
GMY1Wi6MbnXG7oknlZNtggOtFLmvFxiDS0yxv9y/wJK5iGudctqCs+/vpj8+GE7jylW6u8+07iog
FDGGCOSExe6vi6dXeuYwbk9pouwtN6XIUrei8pwcVlXA9wQIj372YpOXKVUVSqdfA3TvGTRpVTai
azSqU0rnd67MMu5ReJ492olBmd6I6oZTDMNOv2L8oVskQSwmciJabou5O2eQzr/+kVpNOSFUYMOr
Oi9gHFMWnm/N8J80bd8+15Tn9+qaoMkGdtfLeIayAVziwYYRSDmafvNRUfMawvXFGRmgSrmCE2bd
G9+xwG1gQOCE42Yb2VWAbtIFtPIVpXOFS9PDMUoJ+z0wtWmeKT3DKcNds/TNU3fYoH9/0J7ESNOv
Miq8R10oVzvjNbF5PSa27Rbyde+1R/0uEx1vn7udsZ92wnYgrYJhEAFerjfJakIuThos9N26qPjH
CoHviVPRXWHNx/PMCB6sJlOvegcCulrtRK0sRjM7eGVFLGg1ZAQv1C5SzFmdKAcxmYskPP3ILE0z
aMi2uUOeMYjqW+V9WKlt5M2uv8qX+ZbSh1aGS7F60WkhvdoniAq1tN2Ik8ZC4NUSvx+JhSA2qFvh
1jEpU4Xtv+Tf4MQ/e7hqUBSLl/X+qW+sDjNO54quNdHSMmO1Gx6U4k7AeGO+8GEzMFDbk5FtQIM0
kcBbCJUdCPunrkPsqwJaIyD7BVXrZv5jFCAVhN6+jkKi3A8sKHmT3U5rM1GAn4/pAAG1S8Icei7Y
vyunzmM1EJqXtR2JJTO/9pPkFfi1ynM/0SKMM2xVJYzxi9Zd1GWtFedbKIHpg1gmqnFlcBEaO7qM
mUd5SRZyVVDSza7IMNFcWjxxcnQWRJhSOxFX6E6EHYq4hPjZjUQrkTIxbpCAq6Czba2E2TOui7uc
2IFzsMvxgnxe8hmCxCf1KfK0mP5z6PC0RCFgL5uCu0bhvLbAnSrzDuVJqubrZ8Ol4lzoQ3Bi2uZv
3xkvr/ftED4BCfSfffgBdZOs9kqjKPNQVzrcSFYwQz7NTImi9GIuBA1cWfDh1qBBdoiiPaClWWlo
YuucXYd9i//20QeJAxwAAWBLwofwT4ouasG8pNaDZ+3xl9WsfSVfcsCCv96dkD6gDOXZnA9smZEJ
xJZBTNufW9XNhLFXm3GPZdezeoU0Jxosq+KKzqCZCNy211KQYRNXc744EMOspp78Rbg6BBLT+kmD
3smc6HZ2T9FtwU2/pgPEnlKzGdKyRxzXnjB8VGvYHTXE7goZTQikO04/2D2FE38zkZrQ8hjJNhzz
LcDtIyvwaothSz+sLobO4fq/QcTE1Xjh0JU5MwJ1lP7+XY0CNtE+4P0ZvxnIryaw/4WB8ll6FxYC
mfygI8BD5EfcWGBtWpfm7Jnca1B9XLiF2u+yoEpVvEj8gteTBsex0FkqlvWmUh41+vE1K+Ln4bCp
jGC1mvQnlvfOzw1gzB0vPmuIAn5jEBO3PONGZRYxRHSo/QFuFGXxT6ZzC4g1SrH0xWLdTAtxXhwm
3t7YvWizQktIfnEewWtdBzmO+c2gETjY4zJ2lVOprN9AWg1CsuJbE3FQ75QwTJTy0CccrzOZIRH1
MRA2X36XkD9pQFHokkCo9kf3YATE4jPGbz8v75ngQnKX1QqsZgpeZnMXDRY4abJFsnGzMBpk2Kho
yEMAKVoO3F9/cowm+mGIi1rqtMOE8X2SXARFa3jIqeaWyxuWwyjrzLv4Hnwwr3a+k4au7+1X9qEE
x2yX7TO1PFlVAHVttjN97GjbCck4liAaNiCyrj5PrQ7QCwniQC8u72ipc+nF5gRV5P7hMP84+hVw
/DOvQqeObto2Qv9rnct2llAiXGFtJI0C0HE5zEx0RLMke4ymAOmL5JEnyY64pfV7snqW1IVVStJB
wwiJv0hhq4B7XUCbaLc/bzyvjytMYmJRo1lzh7jMSUDC3tKg5fR1tEao9Qqv0OiVWGQA6PAb9rUt
0psTw5bVTHmJZE6L6wOYlkuvDgeS81StNZ33ePwrcfPujwC2IrV5hjNBMvMlzs1iZVxvCjmZiHnx
UJKmLCpmZyz5MjDgVpTyFJ8t5WTdpu8HWqJ8vW+uqnm6cttA9Rg7HI2vDeQ8T2ig7iACaTxtwayT
kJvoLIDPTacbr1dFwisZfNJc52h24Z1Gp7c1MQurthZEzxb3Q9MDvMw7dpqHbPSj3kUQHqHKYgDZ
AHX9sZdKISR0VCocZRs7OyvDFtMbZ8t6TbisR7slxXMD86UyIn57aPZotEigYV5sKzO9LlfJ3pwp
UYi7ensmfRujYFH5kYLr9Kh+bsre/HaKezoXR/euBBtnulczQdE8TkuMlw1JyLnrkpcKrPwZhAgW
Ic12WGNd/PCzDfsUfoU6o2zoOSXvRo9A1w9iHVIXhzFUIAFFuxRQYHt4yisztQU3S/NSlEXF0D4b
/8ukcmoIZ2wW1gNh/05Jj8D/hlAVCN3hxH2XMUY6kiF9s4yTFy+8Y3jk2sBbvX5EQPArGH1mJ+ac
mqpdZB2U3rHFihO2SgkKtoRF9WrT6BYOmp8H1GGMOlwxJ7RVrdSHe3H6u/J0NFZrFOOVqL251p5S
WmPczxYptH28XIIDF5/rAdbX72s8Xzz/M74AK1cNrq+df0jxaQwOxV5J+43+t5KGu7xXoDi+mvgG
DHB6NoF2yP15fwYgztFN2BhwvOrCyUSvjxeWQ0GfSmUKMy60pHtXczP3pzOJUnik0tdCI864FCU8
vqFtLNxIEMUgOZ45x7KcV0VeK+o4R4O7F7OTxL4udOYW8M8EQOvQ1UgIT63R20aKZJUMV9+3xK2Z
KHRhBX7l2fvcAI3v/uiVKiHBOzUwQwJO2SqNMj1FkD/uq4yQnc2YDrZtsAsCae+OfLzOv4YIPvMM
M1oIFkkAO1DgvvyBBSTgltZ4XzWh5uXko+Rce9wWUndfjlftCqbEeFg2D5q6kuU3aiJvboDNBSml
0dNkwTolmqt88VEKfeTTt8D/LqR9XUGBg7cHyf5vHxN9leakOhCwa+EGlQGXe1i6DR90LnNr6Dmx
e1H4fY4O4ETeS0EbVR7x4BGrdqmxcrAMvgJtY770cygBbh84bp2omKaHljgsQcndyLt+IfkaJ6FE
xSw81+hJCWq6TT+9To1PYLYSLV38/2d/STPykehaoKul0J50vVw3eMdUhmlSYyR2B8YMS086lDgJ
R1dg4MzYVmfxKptebzHVymaqmZeW+VG5HQFeYLFc6jxn1Twv3Y2VAmtvheQxucU1vGNvnLjJzG2A
yyUTKcfJzmjXWAOoIf7xlDQgAU6Q/DuTAUs/uoJ7nJfXnkPJidKONU+mSxMurbDQU5fvDTMVeRr8
BebVHe2nuBaNm97RBiqsgDwTvil0TuYkgAbHQzVflZsrS+KQTvQVQXneRsmeL53SqaMdpEoi8eAl
SuPVvgS1S0uLEhhsvQCZkJP9hoaOsp95MX/3pKmEyYmdtxbQrqdDVA9SHrdL0ycvW7r6+GWU5ePy
YxFKCjbhuzV5IMcVx4DKzggn0I0z7zKi0RWYz5++rAZvRvT50icokAXWwDnRbS7xs9hKwfRlYIer
IBEScb/zAJo1LAAGczmCC4mIU8hsXXhg54tl5J9Y9j8WSzJHoR8a/aGLV3hPlu3Ll9QCLc1wY3os
NPK2vjA8YDmyalfJ81puS4cKg3wgdyCXIgGBYtKJzza2roA4mbPP7ZZiK8eS5ViJjEpSmfE+n1Im
DW8Z/G33raJdCNDLqXk6ODLOwa2MVWPoR6vxHLThvGFvoO7UxNixPuspv0nvC/k6FiUYNxisRMt5
cGrNuZIplROMVYHvBQjIsAumOKA88voKKO4k1hiXOUpbgl5Eiy/jRoQKbLFEYrv/RhCIWypGTIYJ
lPs9ZYwBammD3XupO2TnlYfjSFxRO3xiPBIjvc2FMHEBYvkl0Mku0S8Y+sLV65ufgqlxkRX0nGqF
gpY3CvaujoZcZC4zRQPD5nJStQG7poZ1AxIJMbFHFQa+D7yw4H1gtryBtq5oQwQ7urOYmvOn17YG
vGecUXEedYp65doqArhM/oqGhVIZHP6xVcRCULxsSu/WkHaiy+nER1/3DckbZOCnqfN8uhDWn+us
A9WAdyjelLY2NVlb9gAr4eMJXnvJ0wLG77nF1FDMvOTAKZDS1JgGbG6oJnpMhEIkQoQVXfa4CtKa
8sJrXMtkAfKJuthcGdfBc7K/1bVTsJizA78aleX0EcK9mdZS75zL+Bas93U+zrKwXiCCfc1+TXwu
9le5R9Klrq9Gd4i1bJAAtlXfauYQ1ke9EHqLGCc0HCX/lNC9o/pPZqKktooJfCYVk/1u0tGuY8uN
4CPLfTArydxnyxHKGzLGw8bfwfT/VZePCjnh4g3H+kHADtdEeSu762hBFc+Vb5koRrnZkkmDxpNQ
sjoyJNjF/OP4BRlfT+PATQkU0831Yk7nVf5CrrI0eA4pJhAQ61UKyR4tBaU7cvfoCGhRyAObEnYf
6BllPppPLx1PIWVy6hzcBNHZNg2zkkh1uxEBz/0D41AK8bNF+YCcUGuB622qVF0rRR/HYLFp2mC8
DXg/3oyBy/h1MZKZ4CP42CneL57agZ6WrGr0sGqlI+ZQjKkA7lTZB0Oo9+Qj4OqiYxNArCuYbxK8
QJPe+zaqclwwSuJIDwBC5taJNERSJ+hbxveGyWGu9lVIXBU4zl42wWurLj7V2QgmRQbGD8LeJT1B
eMt0gpeK+X54ngSTqkej2SMp9p+W3KzcG21//bGQnYeJKisgZZJPtfHq8q05EGjck3jDWAk0vta4
tseZ9CRSqNv+SI6C6zslHO4yh94NvN4xxWpTk1Qu3+4PbYdiVHiRT31tdLu4t3s3DTWYZgZJX+lA
iCtt2KlnnaBh1mRivMIqPrajlFaaTPITQI3qd6DKvf3flG4hj0FBT7sMtvT2JTmtF/oV6utnTvt0
tOr0WZ0FxsHJ+AcIjrEWF5FQ6NOor9ZFPe7bLdltj5WMdsZxKdSu1byxaLDQD/oZeC3Qwwj2PVLz
LnVMhIBb2vEFfSUaujkw9+R9P2DdNTeb6tdYGpIr+ZBlJDVjeyBJ11RswTQfP4ptUtTb6BEa3RH/
ia14CETL4fYpqRLyX3wvOLeqt3zAGBWrsDOoz5wQsNtISUHEqavskVRxUWt97KuiizwZMtXRN0UH
/r2Z51/juCLgVgN22DQeVabXqgaG6AGxziWN4NjyIEmgw6atns6O2+6TDMre9c3ZwwLt2o7gvX8z
g3+jjcRiDpn333SsYXZ0QEBV9QuGLNgB+OSSRvItUfvfXlwXZ+0UNbzp/lL2/SA2AIbLQqKsw2gQ
vudicYpsefeXikUCL6tLmrlq4zu/gbD/MiscENYA5vFnCqB1LXbSdJrTyeHRruEhhKpYYdopOXbo
AsLYH6ORNjEIlgADr2+aSc4P0hZHFUqyCgx2AQuy+UtdWiSnfc4yyGQZY6FgL70OPm07416FPMgp
3LyNEJDPai0+MAs7h+jConDIk6Rg0JJ/XMEgdDJXnlsgsXVbb8cYLnGr3kigk1JR6XXlnljc3s+S
YoX1dAvH1aOioUkCGZuWEQdpPbsdYLqHZ+rCRVRWlsRHh+Br9TDv/TYqhsJyhRbUfxCephbiULQJ
bc0KHRj7CPuAlo0svFaXWvVTNfiALfUDREd0dagVgMt2BMo+Reon7lurUIusjKPR17nOFQrb+Hcb
ppNDchHI+QbBn2f5NtUpHFUXbcurG5Naompsv1qdcT6JEId74+/qHxtF5byFTwsC9VflGl8oclux
x5ewfCCC9qPa1mdF7qV7BDpEnJQSuO5OFG4ZcyAVeJIWc1HxD2WUcAPk/iG9HCC0QIsSjoWo5VTy
a/6daJj2EhDLUfSrHmIW5f4mZWC1+o2HZrPbNjEE/Nqkkwz0l7t28hf/lyYh+3SrS9Atr/zgH+yn
rRG7rvIBoiBeLBZh2X0RqLs2ZAz1BTwNUsJWhL+Ht+guTgLcA+4MObNti+nci6gy/c0b4ZAf8C+5
jYHX3UCA5qZS7B3xOH3VQbsmfhrqC9XM5diAaXApBW5aKh1SzTur60+G37hUSHcjIN1vbNs3jzL3
fS7LVeUH6RhrcezXWojR0xS9QWe0dKrqaMosRR7InCw5Wi9wXkvq4TtL+/muYOWEILapHVEOfrxU
MdC3jPTZSvjyFowQPd9G9qEibL42/qM2n8AgWlf5zL/zWC+7DuMyqyX3K4UsQ5Zr69/CB3gjjCNH
mI9DlRMLN9uKhTviQH5xP9xbynHWbHJNb2a8LGaSOSUXlao/woWeHc6h0q/kNZi+PFSWNU5Gur/E
rah8fa+toRLeFGqV2r4X+wQnpd/mFYfbgcw1IagBXf26b5JyjUxy24tJMRcr1T0p2DZBuAWQ4FOv
MoQ7r2gMitpelUxjw2r2edG5XHu+0PaqR+hbXuAt0qMCTbXMWHyC9KzXuwm0hux/haCcJ1szfkug
d6Ylk36O7liBiCaSMsVoovbQHi4oHRzKzvQ78BzLezRbQV1Pb7ULGY1Mvh9Zzbv/iS/Jc2cfy3bj
eO3MsxGAlEnCre9ihPVBDpyFzgvJQw/TjDWBjRxEWMVJrV2ykXY3vLV6hyjoKG02pQ9shYB0HjcO
/Mn1ji7vlr4tMf1NElb+BCTJDGefGmhSkq5mTaJOjRUC/BpSXoRahIjtUZQ/qWcwasdXWeDlEwVS
xUDCiexlgcRCAVLfOAx7VwjE80sejWTlZDfTf8Aqq3ZYSBMuPnclRnOjnGoHrTwdAzXjGPZQCSg5
Spuak7od9elN3rKHCrE0CZv1CHOhffF9U7jS1qm/v1Lu5Drx2DN/REwq2oU6//XEkfc+i3W3xeVr
DnLMdYa22cGQTotEm/oqMwpdeseaDlGiJ7+th7BAH0+InuSl8BUNXkyJsGWroWo58h2OBCOrLptu
EsJkGjsfEVZH5wKogcR2rHRmjDCF5okrKQd94lLCU/yIASmeR++EqtPJ5YnbB9ApiPITyq8wfFCm
k98ZxQUmAjPaDRdqm7HuWjZITqWIgFU79cue8WdvM6fJG+0iFVeiKnuGCTu5LhGwt+iB9gSMfazR
J5ZO8votQ2wYJZGvsYIECFN2l5ljs/5zm9CpNQXEBGeN9ivoZOvOep9mrMFoDE+6JMJpw3TY2sRl
j+woBZULEuLxGXMoZVnks8IcX1Xq+NpI+SH6pLaWrN+5l1WIjJQqRWmDjGv9D7cVVm1S2uN22mvt
H00J8T5/pmIAnySsaYVYeFaqM/ND91z8hsK+kP7rT0ZS8crIpawnUmDiq3xrTfdYmRLsySuLsyxG
LMyLb6Hp6/gZTP3a2g0LkNZ5AhxBtYcPj9AaEJKDgZvxd5NcyGyblvOamYLRyGzrIs5LSpjeHKL+
FyJOgvwwW1Th4OGOlPB7bP0N20nk0k8LSak49CxkLsjETDphK7MtxI10oEhx7RvOgtcwedykr65K
+i4GhJzLekM6pyRftMZgJtULHkDNrqej6ZUZaR8JGsxNiFNkPwEH53Xgi3Hvc2Gl1hkLdZ7BzYE2
3GhnuO4pQbrImvhV6YkoMKULW2CNCymOGFSeik6UthIHNHXFdI+GvVQuEcXAQE+UFQyKjqo2GZYV
saC9cPKH2kreDmKmxKvyv3N/nqdZIvtIn0YeoZyqyyj+rRIwm/r3UkLKaxToxA16iwc5WsfSGOnu
c/SQ23N7cQRIlCVoAEgpvIpOBou3H/0qpVuk2Z+cFRC/gDR2e3LiYJB/Bbq6yitJJF/yjmeDUTxj
p9XHp3K6Zad5GjW+ZE1uViTd75ApKt4xjS7c6696VJAAqRiOCB6LPrxba/Hx99qRb8rYudtVPRln
Ksy2ylCTZ3Wp9WJ+HfuPNR0FPUYxlYRN+EOlxmb6A4WiJu6U4ukk+xYWdEt8GIrjG0a1+lZz3G4d
cwCg/V+dsLIARgm2AQjausYBGSicz6UG5o/Vinqv6Dr/7SbDYo5QyGpzdnZSuNpi+f/S+QXCozbF
+n51aNTLRfpwTM7zObb0hivHfMzR4bGvkvfm8qOr6xjyM/USqdZNfDwTX9KH6WqaPYRqlQ3RZSDL
ujiJu46ZNEWfAjjQ/5bOopLubWWCRFDApcxTgjAU/soBoEUewOcD9q98n8S4YFkPtYapjNEdm+D9
+2cILfu0jARxvo60a8ZPDeKV5sKnXB+Ptj0y58sgl/mEi8mn7AyrhR7RR8T87CF20n30bJ8JmtWl
+33HXR7Jga9U0FHLx7bcIbqIOG2GVBNzGZc+wCOM9dSdgKwiJ8t4nI2avZxTZNF952AuqKANon9M
gUSG0QloAtNfccShd4/21r82Pwc41STl72fOpCpV8RP3i/4WxtrieZch3Djm6Zk80mJ2DxQPChg1
wpQ+AmcHHVB7NkYA/99hVEsqW881q5/eoGOsWqC/dnPduS+hz+bl+8X2rKfb30GNYLuV+2jusiZx
SpIBrJbFir5Exa3fVEauiN5Cw3V2AGxh3X44sa7/CXXCkxYQTw2HGlY1zHJOJAnT8xD5bK3pFp1j
OlLlbcWdGCCdfKn9rqI4Y79MB6gZA+piYUhQhjfvhSfwJf36TqMCSfjuAX+gvCNCJxLdy/LjruIR
N0Lr4s+llcSPB2nqNaKamosQAT7lQgxiFMhIm6h4/NxQlsXhJ66t2K9NXdmMTDoC8El2s80HzL3P
obAbSulP4yJqRsXUS4KcXQqVlO1CiaErSMAtFHrk3HtoYZAO1xwKBCyxwLC4YsBGY27HS/K/KeU5
MX9tp2W+HnexH1yPMLT2fCSD7gHGgV8lbh6Bx5HuQTwHASI0G90pm+mPVvjkLQjTXAi27U9L+77x
TuIl8epM5CFWkIuAZ0EjuOVOoxrG7cb1Ed7r7BPkvT0FSjuzuWrVm3OA/GMWwnyolLmaOstbhm0C
ox5Ybh/XFwEyrvFQO7ihtr88JzaVgiL2XRdjDHIDbP31yzLTicZbqHo9cW+GBpEB2ofBGbe21puz
aGr5MpQ3f08Bn+Wa4nO+7s42HPoLqehwGUT5GBQEwDDRiVHv2uxpoP8io86SyXZGfND0LFyR09pu
X7VKQSBG6pKCZK4/XT+jTEOr8hCzHojq94XgTzO7mZ617ozqK8r/uxJvbmTqlR06E3bgZn++Dx2w
vuUvhOi0SUgGN1cMXWhUvF6r/J9MfS9rO1pqhq2Rp9LrfGIGEH+ctdMdhLmrdeC0RIM8SwwxjfLU
CxwK/mfoSln1GBz2QswC6ED9mJa/UaFWH1TULg3yVVRwUOzoMlWdomNPkKSIEfUhEsZKYiYVlF7B
3CxH4KzQbga7BvR0/zyyEkzT5Bi9ANPyv/ewgJmyVZBg8bCBkyHcduYbx02Ytz0nnlbpwJkurAuQ
k58bF4O8XZ0HSeuPMLO4+TIiHzghEd/Dfjeo8Mt9LJV8Hm5P8x6FlhB7pyDY/bd/PpnKag2sifGh
EGyRLZtmoWyCTELmFF+T0dnGpvzUru3Zjwcl3/wdIjQwLgGxqL6JjnYK6f7rGQeFUOamRmOFCbrZ
xpUldTyqeCmDKT5yXZ02rx86Y66itjqd8IjmajgecezQOApjz5xwFjCufH1AkNYW7QOewHlRKhJX
YcM6OduJKBCDaau8HBuDzp79yR4MdltzKum4dw+TUoDw1h1YzHfcSlixJ3AEJc9W4+0OU9uv6czK
L+Ufln5ydmGaswmo/Uby8cuTsTSN6mdoFn9ohx+90fCcfOJ+dwMFZbgcG72hzJ8bjhBL0EAd0g7S
yMLm5eTiUUWs2781cTpOeS54FxLX2w03CwgcW8ZSu027pQdSXJaIAfo8mwwWkHijwId3vP8Totav
zvn5b5Sk9NSud4vMTgAYNpcNHIZ8AjyI+bm7MZcZFKSReHmT8uj0824uc9u8hHGWKulYOGBUnKmM
uqQGMC92F3NwjEqZBSjZruUJOb65jxq+oHWq3mvlxNJWxnkTHGcSua75bKXV2M1ESkze044dJPxq
Qv4WXYNKonxT1qf2kRODZ5VcKpbmAOWRVjmUgKUlty/bXrtjeOE1o0KoLSHD6k52bBqCOYP4nwzM
/h5C6GG5IO4Ml3HPcgthgI9YF6oPv9m9zlV4sXjIMJd6IhOAi7kTFTe5aLHmNsNXDk8JVnmAHW22
jh3SOw31aKpMJC445qvGC6ISMw/S/Tcg+RmC0dFDywBIVwc6U1U3PhZo5Bj1AmXJgNjgEGfB7r51
zlV46XojX9m9qNRjWBp3yu5E+AXPT8URM3TtPuC9lKu1Bzs9wIQgniqe0IYLiO6pOaAEqZT6ROkb
5fZDr+jvttlm03J5febHZ2MHLOld6xFA//CsorYZ7LkmQ525cvBynQwyEnKuI4TVBLSpA9HaiMNs
OMSCEeu7VSiWYf+BIlh5iH0XKQEPkOc2BdP1f8KaZT9ZggRi5zGdiYnnjmCo+iiF/FHhRuDLgSb7
4YTa7LM2qsA66hKBVk2vJccjdkVXtdKYQ7GAFXSKr2klInNcdNV027mPYn7XWX8+Bgd7XFaC7VCi
p31hAE21jGHa4xtw1YXDd7FoK8wgGSufTsW50N5IpUrNkFrH9FxtcjrwKMo3DxeFCL9I33e5Q7nv
sMTqFV0UNNMIs3CZqm8FfKBdY+JsD64FtnZbhfcvjn+LckaYPjGsj36OxbRObExW5bh/nTLzguCr
j6l17cPePhWmj8D4QkLiYZG6bX6DgJ/g6Uk0NH+g0CM/tX/oz0zSm5h7w40H3VgiT6KCx9naK42s
Jov1FZmm9dtLP2mdEBhHLKs27eANezNQdGVZDAFhBe5TLcxS3bM7j7E32e2ZFdEUHh97+u5UtvEf
Z2Elp+X1b2knljWTz3HbPJcmAZ4NoXUEyr+Cv3wteIE6ry5sIBiozr9A5mFcXlDa5F76SUbedVPc
iT037iZElOMFG1dQaYz1tcRe8x+fZbVxyhsEhrpNL9kzzD84p/89Jexa3GgfOGGKozFvihdq3rq4
whDSgXKK3P1JScBAjQAEQ2RA9TQADySsXG2B2zBsfjM70CNRm+NXev2WTr1dWADO9WxArLkewQ72
XadzHQX7WWxFbCE8ctc+QBcUXURnPbrpOWHbfXr3SoS2+lpis6R0FAnPW8JaEqhzPlnDqa/ooiZm
pQHZdEC3bpTfZSbI/xtmZnZYUWhbT5UNfGZcbT6SdeBktoMmlYXeY54aLwEGOU/WPF8CqCAhObGL
gaYm3v+rPcTQNbMRw6EkoXg7gO0ESx0hxbu4G53Py6gOr+8BlCZfU34ksoAlKHHChCQ9jCc+7kT3
UYBg8BNEjE5BZiAZ0UefeLKiqa5Omoapj+Pt2R2eW5wJgQNlbrVsJNsq1SoiI1EqCHpnD+FF9qpR
gC2o0dPfsUIC4UrVcDtTmORnV5bzDzcgRabszegd/tqAZMhDSDIeoHgbhqwCiRbl9N4T5+XdkNjk
+W2nbilt30TDL1hIHYTNnuehocGZO/CRE5cyE0QOJmtS9wkXoZl2wJG4CP3WvhXVkZZ3OOFNkXwO
pz0u4tfsddwCyePRq8//4NJmhA8Fb7ymq0AhQ6ZeC+F8IGF0QKhrW3alRL94ILthHEv54ORlGnmC
qY/d6CFG2CJgpmEgjzABJlKbyFpcX/sSVWvXKVNNCWD8L2OA+4xx5NwBZPeOuEuzH5SyiObmjuHe
pECJijI5YOaVDpgP5lCXP0tHq3tmcEkgpZYtfjsuywlDmHZysTIB3WIgCMfGBHpCi7lZ6pG85Dgj
WdX0XQFoy6djTWCMmP+m8HQ7Y5Y7iqQ4MKu+cm9BVsNpOj7nL3tgKzgzpTolbbIkdoMg9F+hHyJB
2/EFyqeq0LVx8su+BwKkW09JWD01LsPj1FHgEBVmRyxF7labeIvMKAMDXIwOilvklElxumQV3BMS
IUCGzX5wzh2cuWI/F71NRP26dm+nNJ+T5Y9dsiObz8n0ywtZ0QpJs0AQS6sCkl4KfsIqw5+rtbxe
IvRnkUXwigZ7LlVgJ9lysYEbxButii3v6bT4vLMc7w5CIVLCVfQJcVSGGXumNMABp0xS6mlefQ5v
GfE1ZY3AbxLx2jB/5L4PlXxBZ/jnqcIgo9IWx/7e4Z+AFM5f53rDxeDv0euy/9Nc48z+Z05tFjW2
7XxUwfvMlVH/RUkuEosScvjgxKhAaKlu04mMsXh6UZ9gz+hIz8DydP+o5CQBu+odOB05e05tE5e5
IJxLYNiIF+bao5angM1CLAh1LhGZPLvc0c5XszywaUsl004Tgr5DNDEZ3rP1JwRITjdhaDJuf4Zf
t8lFQ+64ncPuA+tCkZ9DOybZRk2AqJ3JOrHD0zI5r9bjhw+qLiEyc3gjO9xXQkl7GNiL1fAqA0/z
06HIHGG63MmEsvavxHvMlBQvOaE0EE+hU2Mjwvh1iWg4GqXDHDVN5bJWn3sbZaVazh0skBRSi693
5RbuEB5DjWMpW/NzGXgNKbCujGtzWmTaeWUIoX7mXU/veSQkHSnujtI5asEPbKj+fne8HSAOCAna
sZFAUjX1AxGBdZnic6RiBFFvPuy70P+RYJPedI7oyPWpVRs9sRn1pAqTYEtm+iup/zCffinN1Tth
wRyi4uMXB67AW02SYhCOMQ7XI26doiSC+l9BvizpQuSaHoJq2RzezBqh1wbxWc9A/cpwLpBNvWJu
7XqYjUbPh7McFSI3VpL8CZY9QL5wZxt+QrvLZRveFQ9AqrUdZVeuaQl9RE/cU9yB3wVxF5Z6LqLI
cc+aqEs5vYma33ym7Yd/zsK9f+KyVHUPTI2Mfp+So7RqRr1VOiKOjEpz0HhnNPeCbK/2Go41BPEc
JaHXOJzULkQjAPPKuhqk4WHgFHOTWCid6IGIMlvsqco6XcJtguURQB1x9q1+iZpL+g2E8Y48Ruw5
kRGzZY5Cw6tX8zkUdzpZ7LRYTR/TbggPpeeA+ojRdsK8+aqlzQUGaHcmAuSJ3zy5PGbkB2maWmAG
w0PZZ3d4py7qOkrDshDLfw38a/zSDsV9WcOu6gSI4mVUJPMFKac2DvWsTmt/pd0OF6m3LKXebGrS
s3A/lLgMDv/4Ujl0Y9StoFwxqpc/5G1kFqQobJLMp0h/2sC7tsXirHkvn1EC37G81vus5UNtOyBM
ZmUJmwPcnkWNcENWTBFBdIAyyPyspUweAXh+MM7OetXa3Z1+W4RPUs6wgDC/iJaLu4cnHXKpSH68
gMa0/EcOHCD3MBtj1U8sdPRNbC4DERvgGhJDpO6VuzLeD8otnNMAPGIvUT2tr5JUYnwP0DTVIMh6
DJ4x0N6+HBrmjJDzqGU1jrXjmF/DBGXW+0KPRWpNAIJ5u8RJhQBCg5F2aW8E9z85L/nL1+QN1tjD
7ejebh1sZipw4hxdXI9Ne6iISddNpUZc5iJvafBkdgi3mBZj1O1ENLBTes1VtVE5/GR/O8o1UxID
xrICfoFH0BPOMznDNgtdxGqFOOJmLREJPzTKn2PbyS8TCToeKVW2825Ou4QR2O3FOq+gS3hOmf1m
p0epl5gitfpZmJKL/xbQnJvpEcOcJUOjAaS9BTlFbuN6h/MnSlObnfKL38plGAM7oT1dsr0XVk64
jg2RijbB4/NdHTjJAD3i/kz26jDBqlLWqjPeBdGbINCrHbZQFuPPIlE/XLJDOwekxGbL5txFobvN
S1Bp282JfFdwdjafmbGCQlNTyLQsUksDrSJzm/VDC/V0rKrEOezPKkFniw/gloyKMwHV6qpnQyhP
HvPKb2VT3I+we4N458DG9KLvTzZgcq5Clkf/04KPXkQG6Xh+LiJ1/7/Z0pwRGsRDm/wQO7h1Ny6p
tzQf/9BkVwzGEzJTOCqk4Y6vy82I8NWz9LaIVFUAEhyAZBoh+KnCVAPEnnLT4RjwxnjhsDEq1jZb
a8Ij5M7yf5FgwWT1JdY5FB8IOXO6Wg1uExZOE1vThSbZP5DGDdFRBucDyT4p20AaKSvzRN4E5M2W
TEAutEkKua1py6LnuiEBS5yRV6EA2IytIG8U6xcwgIGnJVgDaXAeW1VHt3vxveUXY5sWKXqez22j
rFviI8/iByoDUgvyBkp2vKQq2YdLitWuH2R0pt8LG/8QUCoRuI/99MkTD4fgBwvAn8VUop3u0oBv
atEMff30axoYa0tH5eRVVTzpwlYfowZCC8tqy9Q7k71F24sp/LlRm3xeikm/dxpg9Lug+DKzp/rC
RL4topNehBRq5tVXc1exUiMX7GK5JFLkYCGUBgQwe8n7jIMcQU9Drzc+jT9fiUqsoN7yB7ZPTmVO
0oPVZc65RZNOCxAB094A8T6XLqnfrR0jP2XyiNPEAGLbmvM5Y6U8kI3nvWU1L6CYQRNBYwzBOstx
QPkeLgmNFRKHapr1R04SMqhsFwoFQ9ymuC3QJAbcMaFDXKqHvNg6s1Dj9Y5cMo+JTiJeS45eLZvE
3SZmDhLMJ0S2PJuXJZGYnIrwmTgjOGnP86IhJqslklemVfBOksReX+/oEeFomlskl1wlD/aTFGqK
PDrWYlYlIckrvJWICxkb81aVJf3C/A5an3GPQRsKXNbGUsAoeP00NhPL6hXgrZOhw4VsO60+YTXq
PWcZDnvl3YcLjb8Q3syQXTJZBaR2m+kShcgkIZbORpERHD/+nUD7seXkDCp5L+jLY12tLLucBsfs
Zcj1yXbT5aTpNGhRxPwwCDF7pMCH1Dig4nMFb2UnlieXEgVARx811ZK6f4oaYbSUhUYZ9WKOmFMp
Z9SFPULXhHcMQco4npx8k7U3VSMgSlKbJHLLu04vCHN6zU2vWpJoxGJwXOJ6/r+Oj4YXu2BOyvXm
u/zVZ8Jo8Qx6pdww29pd5JIAOGQHj38rFtKWmZYDB1a1FalyqFFuS+dRqrqD65FqMdUtQc47eH7t
IzrVgLJiKc7bAhqWeEULNtfCGpyWX4mphiGJwJyfenv7sLUqiRaKNALtQxeeVqtMDou/6E2fGJkS
pwxEJfQdnSTKB8DU3N00BPjrzyz24pzq3BgHZSpS+QDQu3gcq6I1bqj4Xm+5Aw9mD/Fx/oXjgcLD
eKyb31IU8N30eY2K5ai8Qb3QB+RD5r6KKVe47yZLCouXby9NDD0bYJV8kXMNzWPxUs/lmz/L3VIZ
7jRhqqrk80uA/3hwD2AUBYVxrxEy1O59g1pwyETs8chvdYImfaxI9qJcXQix73JKUV+FRekb1aJD
ndNkwDPOnG3mlqd6Yx+UFMfqSd+MlvgCeV4zUWuKLrDXZEXfGkYdl3r+DzdRkvhoJIiANY4U5DXL
WIOfhtbjRLd53AskuO9mfWTzSt87xS95a3+/GjN89ACxbkDh79Td9U3mezJXC6RJkDaetIecf/p/
FSEcGpZSma71/R17UrmHD487icYPy8AGSz/B89YRIYKI8c7Rnfh9Zpf5nws4G+lO2blRQI7tFwHO
VoHHzf8LIU9OlEiTXwjnIuMEPaLMVBI7KZSATYc3Xd+0lcs0NFa+HlQM2u4ukeLA3Kk7rt1dCPdR
WV9ojW2RHmyTm8M3EtdCLM0Karo57SS1M7bXtDzYXQycEBZMV+8Iiy9PnfAew3nPeMbJVU77gbE8
A0bVvZscs73FJ/IbRRxlc/x16Pz5zrdfiFV9qXaIGpuo+s4BfHuT5Odpw0buc/W2AH0UrvheN6bZ
hKydWwvpUIqp01+T1NlsImAwn63xCf6FqRo9DqN8cN45q+H9O3w1fMt8aGfwnoPelsLqRCnmA4Ro
gg+TwY6nl81bN4p4ijBiazITZWx6vk585nJd54+voqlSQSR1IOOrbIbLCYRJTYdLQWxT61G2kN26
eSjSNOTVO6S8fc2+TJHJElGZls1gVL7oGM/7rXUAmycY1pxNn0w8APG5R6QQX0wc4//g/DxhG/yz
LeGkYp5lfu6IGqs8PTrNeLI/VW2YsJCqgu2ssxlpC1MR3frLjyysk7yeSKWOOBr5J2yhU/ootDzR
388/8GUKdh24tKLmjyyIJzbMm7b0FJYmKAaN9tHPKJL9F9tyMvyhxQpYxrZzviAv9/bnu+FWu9cw
HV+gxsfoy2GOijQb3nfGZSU7NAtyQGyz/jr3+bfMxAsPnuWIwVRxoBPUnsoy2O4DXaYqoAAQ4A3G
gYz9uFOt7jyDR5dABvK2+GPnhW2Ywn5GWSaJHbRxQIsAsKHDPRFzEbqvLl4GaWDblvEsx6UDAQ4V
BPXduxfi3RrjOVXL0RQAYBophlAl0rIaIjxIupoMXa/SB+lVuLEa7/eAvNsrdCYZsc+xDs1Rqjb+
wB/57nSyaEVkZDSdmWmhNxOKgKSM9j+uzgbD3oPxg4TSamkND1Vhdkxg4heYSC4+aWkUyFgsqAVR
qxVpOMQUTUVsWtwaPS9tNPr7LV/tKa3BGpK5hLqk6gflzyYhIle30NdOQQsZ+1pJ+VX50sz4126W
nS9JybleOiOncLg/g+dOnm8Utj5sygUct9cJ98amREbLh5mT0jgvcOz5utFK8KosuTa6qpUIChgp
xiVSZ5thWuZVgjziqN13hue34VVzG74j4xMnPJsz92Q18hGcN7Bi58NLa9OUzBTsV+lu28HD4sub
0PQ9CLrTns1eb1Mqhrnwau4VPnydOqEUG4NwzJuGZ7uR0vFsU0W2sJvEwKnRlpDpYBPbWggcHoSC
q+/pnIAvaxNv3U5EEakt7YMu5tr5mbzut2BQLCiQqdSeUMAj7z5+cwjbPAkTHYBvnzJOhihTJwwk
nZsAERo1bSbRQv8uhb8ZbnKDQPajwYeVku7LdLjoCMIanMyCz7gw1Pm/uIZnSPklniBVCLwnTu2E
YeHIVfq7FLeVJgga9v19DJEMlMjXzXLclWnKt3R0HEn4KJNsCGgbliUec6FiT8M3f/eVVojAVYAY
VNF6dKojSWTkDKy6eabSi87X+7Y3MgODHwuXf1d5+lc9xetPSc/xd87a2ZCJiO8fhV8R1S5DcIKL
pGpSZAl+yKqW/wix0fIeOFul8T/4GMvcWH7DV19qXiR2/eRuCljZ2+bMYuwi6LgOXqfnT/KD3xhm
Yg/T+BVw1afpY6G3ZcEY7xh1lMurTH3UazjjYUvLlqWfATkfvsWSXyS7hUc2UF7Q0ZYpw7fHSV0d
ScuJe36mTIPKa6mHgGum0KdBTJeGO3TBErqdKa5H/8op3ygJYJZpeBzJpUwQamwfuM6ry9abbVZE
ytrpLulHgiNpaU7DsDIqk2XhNDQAGXL9+YWWfWaDx64JQwXFxGc/LTFaK9rcd01HelMCzgF1jtna
uASwk/YA9WBi4uUvw7eLfHkewlWRD8vvQjfpA8VHAeJQhRM3gffnUiADTBm/8casrV/Oq1yeHWSt
r13CTRWmvA7uElITbNGJjAgl9uncISbm4X9N4ikwVEcr6uNF9la0yox/OghH06Mx/UvCYsYTYVLo
B++BU89utxRTLhfwEuxRRPS3i2HRsZh8CVTiOERpDdGt4gYip8nRhE5U3ZDVEt3W3tI0cUdLdFJw
YU5G9W1ojJE3+GtCr7rJ+nkvCOGst4cUPBu3KoHQKIe12PgIUYuDLpFxT4b+Oob1DmtlU115l+xD
4qbAFdNY94zgVkVPkoxwZVTQzcg4r0DNThVK95MDs1vujML4rzwWjxa9ZHP4WXXHy/OWpmlYXVPs
ELJR5G3bk5kGKOhcIzrqC3UMxOvlEJENWbzvUoX0T4uDiPqnOpozzaXKqan8wTRS8VJoDhwhMYFT
NvEpCqX1Ja5K5j6VPh06rtEcnH0bfPyMryio+q5BEE0RnrXQuV8fhOeEGTZLMFq2YhCU+IDfKsUL
dp1gDz74b0tohaEqoT3jPae3pr7ANwgWGuCeRyf4E3QWKt1c9N4e9ukSbRircfngHJNxKBkmTVBL
zj6AW90xEbzYX1eCtZRbgUpZXiPPIrMyfDEGL8XfQofPWdShlW/hLXBueNoFSYtBZpolhMyf2aZK
A77qrVNdfVZJorPtFkIq6tgLLAMjpkwQz6/aSRZjQ7ZBAu5et//ruSHcK/aXY6TVGxGo/g1wibmp
/YLzOK36kIl3DvnwL76z5WhDvhaeedBmOsHPLQTt+qhaVj+c44SS5rGaK7SWBEpdQb8gSbilQHTs
UVoj+iIgh6vFC+dKcas/A1pm89R+MzX8llOO8/YR8eRCsbT8L3VTgsPbXPDxtU3g24/9a0Om7N5X
O+EW353cEOrW8I06c5ee1KCfZhIw7QLXpqXjAki/wTQ4GdY81FemBuQRRKP5/mOFOTkHzdekiykS
Ejdddr9ipPQRXrfNvQ9PHF82Ydpfr73j0Q6ilWyhrOq3UTv7opLU9ksM4Ga1g5ZqdXyKsqqa28qY
C75K8IXfcOdy9dl1VK6rESOKA5zELVETlH2jMxv9xOQu2421BA829PZCk8nj98L4okj7VWVVy64d
fxRgeSptXvx0dMlBs3mHkzIdVF29cSyc4+cqjh/VdKp0iDqHO/eg/BQQPqnjggI6nxkXzZtmlea6
9GG9eKyYtESeqCT5L9YInq2ehxjrvUUMq5Lq06SwcQ1/yZ2RXsD2NEFfTaDzTzdrHnKdFLIyJgkZ
eVlLADmyMCuzfzRgKlFsIIm46jjlMSxQEkf0h5ZKgGS1l6q1xpwCVqKXXVwb0Pu5/xPa0wLFfQoT
djBLpmFONaNEjY2OZtPxAyVWyzFBk46JUduWfTOvrIkhJQgUOhXcvWQhNaziDTjcMLZ9gwCI7IZk
BrrRud6iMreK/dZjJXyKjW9SuCVLsc+qC8TND2k7TFnTuHMWbABUqUhDgOIC/Oo0sXpicEwBtcSX
klpBZhRU6grttRlCuSArm7LeLSYLdjlkhNYBOQK5jP4Mv5wfzTVmFF6jiVE6jm5PhQhPbX8/k4FK
om57lX5uO5yDgjZOkPBd2lH5548AxKMUL6mV3ZJaaCiFhUw4KWkQhc7ydPfhCktDzujTz5r+fyYY
DATjYIaT9O6JEzvkEl3ID5gNlTX9hLzW3f6ySSFt0b8SvnGvCeEfUqx7TQRPCg/YGlcdXUrwGiG4
TelgItsdvj4/PwExlubIVVaphFfkm4/hp5CwvPV2g8uLvYAa7iWOtNZFyv1HiSYwETdwOIjMjOrC
GW9nJaxQDgg3Ja+ofZSA5J6v+ydmWrSW1ZcO7XMFUTmlJYi2Hz5rGaD0KdY8exVsswvyTlOV42Qt
u9bMaHy95Lef6opoD3vqoWsu3L77FXGdO/9aKg+UuLXNaYjgDeuR08p9ItTHpR0XstRUx9sW/qn8
QvfP1xuWJtjEgFE3irigpWFYQ5BhaPmvmw/A4yayyLzKHaSZ7f++y8ErxetJEe0vxhlwwl7rZRko
7F3XTFdEecp39Kh/fuA0wbaYVDJCsRVd0efjCvjONIt315/XI1H8WHcB8BddgGCECdbOrUy495ww
5MfxWcdy3f83uUB1JJ7xG6XZ9JLDZ7dUmfHjir6xLGIG4Ae6uB1BQ53pLXSQ3nyJf/rx/kc0Rx4Z
ybLOyNPO/n13ZxHSWqC0bLZxGf4l1jP4vw04X7tzVIuKZBr7iddBvSUVY3za7wcqqJuaI9CntkVb
IbXg4WVaT2lDPsKzHp64nQlHU2C9UGtoUdwvUX6+mJfzjXQfhkQapJmmODjZ7G3Jjy0mNnju6i0D
EQdB2pdz7Et6PzKX23gPV75y72F/3u9aUJwOBoaVL/Pl7isF5SrYdDVbO/TgdC/ipjF3gtJoyECK
pza5pn5Y9pUXTTf3vVjmzLKdThpyj+oXMAFqBO1rRT/wU4DOVBErVhUQUlrslf634/j55Kq0rP51
AY97+HFlkv3xF9w+Lkv/HypwcWstl1brd3vCKs7VZ1dJtaqa5KFrcuT1JXIvxyL9k95aJXy9v+W9
AKXwMjWYD4hHYeAzfCLokatI1IQ7wq5/hDDvFa4YOO/Lwfp8S47Vcnmljm8NqrUJeNf7monlp6tD
K4rj0QodFC9hthlMZS1mSfTq1zqdBm+6w2S1cIWZGEnIP8zh6zMPKaX0AuaFaCoFoC/6oXqqho7y
rYMyjZTGjPiGQWwbXoNE5EnHxlefvwG3bZfx4sTbv7cR2EUnRwF3gsDkv8OvWZRPFau3M8V6TYMn
50SNxpahST3TZ02qLxmhq2gw1mL+w4P+bbl3ZpH1U+IG8IGfKY/pv6mFLRMm4j/rsFJcLwgZOymq
6ed/caH7lQZY1+Y2pqORKKrhpcKOdR+0F6sbFakJOkfC4Z6jFyryx+i7V67PCsNEUpIFBileFHkY
b5giXtW4ahHMMO2EVTSSTj/8CmWUNLD3JhLN9mY3aK6LWl2XYQcio0Z+MoAhiaDvxomZvnxjMzNM
bLmwddJFsRp/SAK5rnWFJBbKFxQlhIEYwiIGXw1zi7iimtKOgemOd2m1WsQMhn993tc9FvX7PyXx
rvHbWsEhLRKUNz2X6j3k19JRuNzBNBRB6heOaD+ww+eAlo7iZ1n/ZLyrX6Me9gdLk14KKSAflpmH
jnMrmSk6GbvJR9eFmQwvj/8eBLCIuFFj3M397+YfYgMX3lfgzCe6/10BpV/IuK2Hh1dbzg3ROBtB
dZ0ZHZZdItk4UNewYXiVpmDUtjfI+Z+4xh0wYMYEJyxB8HxdscJKL515WwnVj4t/WZ1Mq99Wpztk
+gtoRYTPrcZbzTJaU9mWJZfdFabxSCEOwSVWP1rGHEQZ+S2nQGDWm1t6UNPuHk6cybIRSMXzRtkj
5O1kvHA9RnGBmPmHIeECQWL1IV8cT1E4k6l96g9nMKfs8TW0e9gdc6YTmIKXhPYwd/X59F7ATa9m
SbY9VCjoB4hIXKqID4Y2tiTM6E5HmHjI6pl6tz/Fu0sWfb3nvhBIZuZ+fM/z8ctsky6JFwhCrfSv
Red7IFmdDmAcb0luZGW2BknV92kfpH6h3I4A64aPA8SBrOeICg5JxlFDlty621ouTPGkOYb1wrRG
kdOUUe4hv5SMVzOpURI/J+/CQ7NBRU0YV92QhVqifY0TsSgj2LThQzDjfyB2WVwu4/ocAQZmpPlk
FCoVrvOCfydx8Z1nwSi8cwLI776C9qoY0dxccMEy7C9eQjxdLhntyGloCReGXkey9mZ5iwIgyNwb
fvE2XK6941RFzFSJjHxKw9dftLj6AxHBxlLyC/uVJYen8kv+qGcsmpcgAGGbqHIvscXI2kw/wnkH
WJphibb4OASkXj205bMgzfQid1sOVkvBUBXvf1PAzWHTaRHDuQIcPKKV4mvP5IOIX+XE75tah9Wr
rFoWnuw7X6N14gjdy4pkJtl9i8aFpOcKQxiAZjASDu14hB5HfuKrwzhnByWL1ZaEtat8zNKMJzHc
Ry6r2BOFMSf6krgXtmXTM5jV0JPUmLqOOwaGBiV3cZKvugjYWRegQsr2vd60KUbzd4YPbRYzBDqY
7INJpqG8xlU0vRf9kr6n9X/nFdTnlgFmJsn8Suz3UVYRNMslOJMHaNx39679mxyAd9FUIC90qGnR
PUimTBkgefgNDr+v5gM751bXmHThWERNnrWNoELgVCch3d4bomrGd2q3rEMBmlYUT81Jycz2ibtR
vyIS0AkcI6Q8JsPvVoZzCLcTwpX26JedaFomK48U0mQlUC+3QKXPbRL0Qu+8B+FtDSnCdzDBfZe8
RRPMzJcD+YV6+GzRcPVkrPua99LnuNZHjZZqHJtHqn+0aAFg3XoJhxv36WLU4OhkVOMgEGaQlWwO
PARPFnBQ7DZFw1GeydnhQQDIo2L1M1+k1HCCY02u6xdspRQ+cUWYURoM75n1N50FZH5pcxqyLoBi
tBxLmr2Zz0I3Sal4XW+p7+SFrh0I0sUDlaMta+Tc7NZnPMa/faP+2sHthU/x+YFtgkKbXpQd4mcm
keagK6CncZ3Mwk/132Y2nysQyl+AbAxIwjyJ1BDOEuupEQua/vRiGyo/X1r8/BCIhJIlsf4KzPnp
31Ss1IhP5BHcTmNTSfPqNOdoietqrUcJUaG/FMlaUUdxUmlok9VjPfs7a1ygo5/v41aGBllu1LUo
svLUYNU4QlrsPKv+1Q2oPtqyD+ZR/Xz/bUUV0SwVaaIBF37Kzo5+cEnuWFnqKHsLUj7jYF4VOZRF
mVD/qaIjffl1GndBsHLG42n1hrSeAic3GBNZnTTH9JVwy2TMHg6ynlrjkOK1csFl9lCbda6b599K
yKGz8InL+shFUiHKrXZEm+e19A2JgIzglVrfS0K+D5wETjqv35t72k8qoZ398zDjv+1RmA9gE/O8
HbndEGRwhft9f7kZrnC2dL/qUdQLMGTRhJ5d7aYYDXU4ZU3gyifnzahFstfZu8IvDgbWMFyFzTZx
xvzmAlU5pjbCrMw5X1SymoGQ/zieQdkjN03xNvAzEnnhHrkiUP4W3KR+KfYIrHHtMhCoUW4QjIRn
HiBfWxqAkeUWuokwTlVKkpbi75LLoXWhb5q0loe9+z/XUwZe+alITUIdyMoHLWomlL9QxbE1NFDZ
j7S9fQoV0bdQuiuajdldcvS95F9+vgxURHkYe8vlLqBTN0/MjTSbasF2WhDlwc/IHZz/euHIMpqy
rdRNh8J6Z4Fk4H2+iv6F0c/IqGBRUoeRBnVahKNnwnFfNytPBhjBh7Ebv7b85jLNaynODvNq5e/b
jQIWjGMYHrkKpPD3mi3znW0qYh0I2f5nAfhMrZlUJ983Qcpxk/FRkYqGcodLWsx8zugbHrjgGWg+
3UZ+JF/2lzY0ZLa23+RMG5UPZ6g86AIcuc2nqUeq0KntieWhuNV6g3EHNFnBYJamlDTHMm5URbyQ
KW6dlfAW84+q7JB8HlXS5UJUvDzDwCebIko8go9O2kpr4uWrH/Koyrx1Cmv4UFnopdyIpUMGapDH
eJ7gZqnNvPonKMWUnd4HT/25qQo4YWXnqbD8EwreiGgp1zXXOBHrFYLpFMmRbO07im3ye9/L+hZP
6mCI+/K4KsVgeu7pQtyMvBVAsY4Vnvn9+GsKl430bBi7gK3aEkzuUeFaQ8CLMnbNT97FrHVeJRDb
oybf8VS3p/1XdWuCeYIo9PhQQ7xxacJTlRL5+PJ0G+7VltdiMCGct5Bfdmyhqh1zLJuAPU+jVuAW
ffda/xijGcrfWiBZfiuYKGCsyaVtY+MRShhWRWHz5cUWUfSLGLjZfqLkM2EbrQr4xAhmYaNbQQd/
EbeIC8+rKE3gvH0JWf+ARRpYSOkOINUPvHDDvMhVDIP06FUXFODYZ6VR8fOpW4R7aINZIVyY8mdh
tE41xfctVJYpbwe/Gx5HaPsXjq3ldOW26eafWrEO9AE/JYz4xH9M4AjOxwLHa75Me3bFk7D2zNLL
nO+Wdnvh6vBMRE5A2rEJeVAUdnD6Y9j3VU3Wq488mD1oxYM8q8Y5wWGORMuuimVctHK/IjyG3SFw
8SUgkTHgOY5r17lqbAqwu7e+AA33mNMEvRzFepMCd9dbFOJJC/rKmxOE+b+5qpfO2bdQljEN23YR
GM27Q7Q5lmVh6nQOj6vAMX+t9FqbH8I9jjy/n6yRVTS9d7O8pKgj7kNbf7laE1BaYGaJg+mMfuj9
uDc5fIPT6heS0BaD5kT/+9wsS4rYU5fR4DFYkMaiuOx/Q6dXpnTDBUbj+bjjqZbagVP+av5OYjj5
Q3Nyqvq0y0ynmTsqEs7SwlUlj0eeJCv16+jktQUSIG1CBD4OhHgXxLcMsZFRmlRfPVNx5hETgFuW
Xmd23Zt9zrFVeyltN6vHI4fby6gwy6vOyVIiKHt/tVkgm4avIbGylXgatYjqImEo2eRBUIepUgv/
qS5i4sTMizaBjeq+mHZvKpKSXPbuSmIsjFaYayWIfhtkBnj2OB1+EnflSX6MsLk6jCP8pSGuPaT9
XjQogYVEyEiHGQOFTe3T6p6grydCY7Hg7soy3C8IjO149XOH9gSLQtL85VRSo9JVm6fvLAD4+IHu
VPL6FDY3csCe2nK2V9gbpHen+f9HBECmy3P9ylITo7PFuhyhdAv7bM3W4Xih8w/Qq9N/r7NAN0R+
VfDQmxFR6rHHD4M2KLUEa6ePTsmqXDMxJJAduEb4Qtv2wQ2mJyrEEV8wgJaqOMc4ach32La3pfIw
92QmnrpdX+y1D4TA2bkj0Pp+ZX80LAY9U4sHpStZuJ5RdgBcs0c+ougRKJe/s70FVUIGHLsba8Sz
hWYzDm8Ecas6x+50GdlzK8MiOL3rjOpLylUa1Y507ypnvrlnqjjfqUbUII698zu2XGsFWJPeym0z
xpcB0C6isC359SODamL2sFELo5RnHJrK77GB5E2pAqBTzE9382fyT24Cv9V8QOHYsaEDoieot1Pt
jj9LMXwppQUYRZ40w+LHrtQLtlMbI049g3yOBJgh1QfWOO+ECRjPIyYah6/DOZBBcLqW4EdmJ88P
PJOyrgQTVHx5J477vihIJ8PQ0MofU3/F0Te8VMSh252Y/moWt2JmYePhl8oU95uTXsDgXRk+WQFH
3I0Pm8J1A69golVTQTuhWhLNYXVc9wC3d5JHlOKem1KVd5K4Iw4bR28WA0A9W4FJHG2Z7vecoamT
as+RiK8BaIIFDN1YcheuNzuJ+bFY6GMEQfQQGqYWONBPilW1pX0YbYsLwwBPExQh6E6NICoJKimW
z5GGm02fkHbmR+aJAvZzRWB3kevgvQUqEvSDc+wYZh1X+Cf6eYjCoTo9lRBvHn+yN3Ent4tTuslw
aiGayqgjhZeJSz6Gj64MJS1TNDtKE3cZPrHyrKT8/80QEgMGvjhuuIkhUNKEyBBQUnn9IoMHysCD
Svw09T2L6/rkne1mRdlOGhvM1e4SpCDJ7n36O4DJP7U9LPwGKNoTpY9a/DVBJapoPg0AbQYHnkdJ
pWVSz8KQcnxUF56GGOc52mdWP+40CzZYqtKl48LJQCxDcPag6v8uWwcyKLJu5CwjerL/wCpNIU0/
Ya2YgcBQUuqYBFgsBFGqxdFMD+R5ViW+TojIKI4bIKLIHOGiWZn/6CLYs39nSM2ogUA2e3X2q3sy
zQAFmOOpFhVGoZTXbcWVag91WweX1W81jwfKP2H9ewPCQE8veuSjtQ2GfJrOOgyc2WelVmDybZTz
36ROZ+z/a+wIjh1oGCm5XLN5yNL/4ZgXAHq0/f4wGiOQXG6dZ+WBMX0cMRFQU/mqdPFaTjN1RtpX
aoHzoN9PzXa/DHphOPuFUFQHk7KM4J60yVi003szTJ1HPDISLfha1y9v/BZqBfRq+AIfRH7Fzj2q
dnoOHvDqOcA225YWZuCl91n+3QKPZaUrGFFwaVflYFI+2lUHlfAIcwKYDupCN/7XNVe0fwgkH7G8
LudCxahRsi6xDwbHGl/L3md8xdZ5IqCt9sKAx+NvX2EZFuOVMqszX9vD+gGsiKatRjM15mPkxZ34
koFjVvT6u2FsHPSyd2QbdCicjDaR1bDqJhnzDOFb4GPnxAeRhclskJ8e9AvXIVqH63aTY1oBeKuM
7HGXYQQWuUffY2sU6WfZxETn6qCXhbFZUlly8VUssHGTauYiuuDN/noIiw6G662A16sJrLHGZqfX
OL8frpqmrXCh6UnUufrQpLA8MZTLEz9TGzHPJx6xU0sM1APqTFTkmaTu5K8YJr77hrGX2LlYBX1S
oK2bBHQTTp0nA3LvD1NTzf/GxsIWZXI77xs9BxxkA+NkjzPi4YSeVNXFtlEaWnie7fDBWAQrVnR5
YRknU+WuNUGl8ho8kIWgdtVvVS9RT6cXNLmitdUOn7MgtvNy291aylswzNrHOOIT58UfMTrG2oFn
R5TPgUihcUP9wx0JDe9FHp6/QNg04DERi2PZUQhPO2Uc3lO9Wtc4enHuHkF5FM8T3XgULN1h32Q6
ny8LNa//uxcwnykBH53+0/mw1mjbYjqpFqVEBbtWZo/aRAwOXxzFbQ5WffIGFCOkcrlDpQtLMaWs
MjP6VGUWLY3OKOtMbN49aXBjyDwDjywawozzZ7ZViuy7WG/SJmrG+HSHkg51I4iatBZsdRxQoFu4
CeVsHaYLjo8M4oWsFOkICsPmZKods7eHsy7tiUtkwrTcuok5hbjeg9RpU2lu816lpJw6p7sbN7Z6
X3ajm7zBKGMuMcr3LXvlBldJlo6dI+yNc2kBOLduE0F64uXBzEhPk2BgSpKiakQR1Szu3gqOUx+2
BVh6b62e3OpqCZiHimaBPa0Qd4e8TJ1u+kbgWWyp9KFJob9gLGq/WDuSkZlo4FY7dQC14A2F0utK
iyhXhlnfOO/LWY/03lPKcB2hw52MFotz5VMB3k0FxwnrywF9xANVVpjCL+2KQV0mpWBNzW7uws7W
Vel3WDwXe1QdZ2JjN/lavX0O6F+Q6Q/SWoO/w+iTMV9OLt2tDrY0bGrMDUdjg1ID6SX0pXoY5AFH
DTESdDFiRcqNTbBnLa6kDEuLZqurwCrJDQuT08WBBOMiexQjxq+SLSbb04BKv8Uc2EN83kWikkra
xBoEoWUjZbc39RL+cY37J6TT25P71WXCXAa0TRO1axyMC2kQHPYHDBZKVaFlvzVdmc377c/zCbRm
/LFYKFpLvoaC9AjwgshZtlXbt1ISpffdrDYPrT7QwlOg4db9mKRwiFCvht6o3mdw3mxlF5+7tLLd
Q2lUxYkEXbWbqRBunzxlEau0K8BlXtKHqmcbKvUvPYD1VhePd0B703J3sVYrMTx11RRGQwMZkr+h
8EgksrnT0P4/7bIjGIeZWnBq4lFrwSsOiTwi5fYTFX+CdKJJxsi2H4jL1/KqcJVUkzGydCfT5TvV
4bARnIZf54jDmCJuk/24xTIBiLZgAIUv/S1dDqs6itJT1daeZb7S+0a12dUiTC57zQN8rumwrpM+
z7LDJ+TVJuRXcIK+ildbM7iNOMcR8s0gJHftDE7MXO+h6+CEk/ApphRPyiUrjaY+bxGbtTcw9bAs
YFKZYXByLFOra1RUHIQ6WFs5IBatl7MH9LF43bdOgIB8zNfeBdawW4VbUoWro0vyTEPrOInQTcxz
Dxp0slMhtAJSWEvPldZMwXVc3HDy75nKWrFUZWedDAAYSyMy2XL98xwKMeciv8UiwFNSUcrgN3tC
ZCe4wpJd68gqeESrgcrfHDjNytDF8UgeG6wCUu0MQa4He3KoMfRwGbimpT+pBCPh8n3icfhfkZ02
tHZiNzHmTNBJUk7JX68QCiXLghWy7z+ngKdqyepJ4KjE6QOJqJ2Gi1/wK1Tf1UZMx8FqWXHDIEUs
4UgQb17jZSJfFtVIbzZCcie+4q0zUk0r2tGa72DUDzLMVOdIELwNNNjYBIVg10vFe4oPkTengtEk
s8A6gGpmZu1QlGaDgLEkdLaHk+uON9/XWL5JnU6cUpgFoUVp9AW36GKNCLLQxcR89CCzn6tPzG40
BVENSrvkkSN9ZnUPVYvQ5jKrwp8MZ7WcSEtCI9YxUb22sJd43NAee3lFSBLHeiYPLYuoImAx0nwt
8i8JS4LW+ROjMwFkk0HioV5hmiqBgK9PGOOCfoqzm/CMpeFFd00ZPtTm3EuAQGBZE8nvrgdJQ1lK
qsyy/AgQCWstSkPbrtvHSj9B6x4+7TmkB5wA1zRNHHH44skq42kTOW5h4UOxo4mYrHzvKOf8ia7i
46Nm8ED35dDtAQSYM8B4Y+hNg8arPpLwI55BIVSZsjnQ4S+DvD6UMPeaIRWfrgjNAEh8fxujQ9Uy
AQd6q0cRiCyI4KnrRMq/e3ifUVDzDWjXHMzYcqI5/aBI/09mrra3NOXmOkEKgnj4gIxc2Z7rLgXP
kCtm1E6C1W5TydABe8SwfAkLrHLpFGSCp2mU9jl4ePU0e3QeE/f0sR7d8stuEEMNdCaBOro5i+G3
bkXlNJiF+guJn5ec4L4iC1Bw3uNAMVI9b0oHabaM/ruU9oSdbj5n4l5N1DdytKHF4KSVAsxbQaKy
eH9GcDBVOPkN++QrR7GeY3dEZcD15gTwaGxFskThUGZrlbG215NOMPjF4Q89mmPnEFTPxKPbyF0U
kf/TYtvwYcfX/GiouX8h9lEExYG3syPbcaymxC0FwNO0RvotAAb2Bgc2E80hOnxzN9rtpAJY+1du
SRPwNfxnbNeFORdlAn3Wg1yrU3AqC7UtHAYvz0r0B5oAND1edMb0zOKo9StpMIhIVO2C3vDTTQWd
qMIJ/mm56CJXCMEXKAWuv8WROgP5N7UHGl3ZygeKPPRCtow3pBgxCnIN3C4TQgNpgyAiDeiSwm9G
pUlk0f6u3mRL8yPxnISooyLyNC4eGXCe4omDVxah8mJ9QCoX9DuBY37SGsz6dc2w/+UgVdb0glLh
ZboxQD1qPJK555C/SqeT+sIxwLfDcc5Q5sGBH7KrEW9tKrLuG8LgeBgD7gwG6kGs97lGfonUGzmw
wnZT+TNkWkte8fNdR1tI5JuA5N8AVYVNhCw7Zn9YCdn5rSb+BEikhn+QrF/83VVqwdQO/EOThUQU
zfufhNwdxkuqBH+Z52emc//eqBnzSO9drxZSGtdNWBsqZgcvtCrIfpIEKFbtExHO8Xkbp6uJ9c2u
MvtDOgbCp7wXkc2Luhc+0mOGAw40G3JG0Lg/2ssZrhhq/YoSWUdYnHCT3ycsiYn5ZZlhqL3xLLVs
RuIo9+QJv4f9+81xO1OXsOd736QCke5C8VrE/yRS5by8rAF8YNO6h0eg04AW31YdZBl5L5CetZNh
elWsRZRBSKhWAdW1sSVTMFJ0GiWx+JxjmlHUm9BAM2gwh/wHNRzx1b3hYt1v1FhdwrrZS/i7Qfj9
uh/VinAzoC77FDttN4qJbFDuwH6WQGmASgjyYlKci6/HLsu1vPWqEhVtJxkAde7CS8EFuOTaZS9V
98pCTXkwyhkdzLDDJCN6xNOso5AoycKvLRIApJX1iNBazn9trqgUdn8elE9V/LF8FV8LiW04zKag
YU1N0AwuL6wlZEwwkjrL1ukK/ZKL1te6QTU3oQN4qE1YIi87vusdttY3zIWAdjAPiaWTLa78IdDB
afL44Qrwz/DbGjrMcoVZxprTKNO8fjCJOUkMEL2YdM1szKf7leizy1jCTHgUj1WS4eQK6rWKU2b7
sa6qmOeXmv1+SDs4fuR3dEtg0ou4GtFPpIN7lLNZOOpHvkAWAEebn6/OVUpecr3ZdjzI2Ighgq6L
bED3jLUcVL5z3E6Z3MwHIrEGSWyKc2a5Kw9AAtAjlJQvIl12KIus/Wl7LWB8iJBeJacMgGb2wdKt
C2F01z2OB0XgvyObZKOJpgXVjhjWkTh82CaCET1Um2XWXEoUM9KLU5wf6R/J+w2vMLIDUHIuvHSm
gvIka4PU4QnRXcmZFnd+ukNf1UCc49ooqMTRIBNqKgBdm9D9EAX4ct3VQjBrx1KC4fcfcHfFILMe
WXaWxSt54oGdl7rsRYURHerMIOb4BcZqX+nmc58QWl50BPqYfdrHOtgORRmtS2ldUPbhZ3O+EQKV
SqeickmAyCXdt1Y0GV8VO/qmhf90/28auuSX7kuyDcf/GxsO7Zlwv7xwITORx79bCZN7T/Hyazop
/dPiCCP0JcSjkuD2yzu5SGtlmhEhwISroyHJdB8Dq61lv+ul6kcTruQ2fKLaMz/fFSq5fwCDcD6d
8HD/LIugz96lOs75q40mYCl7g29CzNoEXw/AD90bHDJyy+oBJxIqkfsQ24fnIUH1h9KU0kEGaQB1
mk9ctFHl9MrBaKLtoinzgeYeqTlCMmvsvT7xG6Rqmt1kGbnn++g0CDxsEfZ9G2o9zTHbTgEYuRm0
ZbGOL0GYZwKHKYxoDclW+0+ttLJ4uuXwwYL7lYTHmDMjihX4E/YWIbCrWG3mWtgKSiCC864V/Nri
djBzq8JiqwLOsogWt6c77F+hEUYRP6dnDjIWOUyGkNxK5P/RSMmdRYfR+Hw8vddkYE6yuQfx13Gf
7hLtNgXVLMyEod7k+CXrhRkpZfJsulkPznZPeyZLmjShGfrWgT1y2yCRndvul4hN/gzSP+MWiGI4
LKsMbnsJewg6Ke+Nj4eg7vOW1Jte7XueAmzMokGVCi/Nygj9XlLZRogqy6VK4/tF+JjwydCgfpYM
OSj4FwA+446uxog7Djke0kzzbwrmGosFjUBg/f704exGrTT+gmVKHmkHUydoFjbUOy1L2XkxV27v
eTh9yiA6eMm820rRWG7QnLXkrPj1Vu3TY2v9F85dJJVYeJarV8mnYMLMTgVW5B2VxyG8st3SDHtE
+3PKz23EtaTpKosGM31a4IyJR4Gu0VBQdDCJNTipaWYU8qhYxq4CGr07kOAQth/mGjcbIRPfKLbD
5ZEki2QNPNPSbK+n1Wk9hbS7mIPqMSCcZsXnyaZD+LkruJt5a3LnmylMwQQr074EApl4qpkiZWYG
r3iztoC4RkaWBe3IYQXg3iubX6yVic0X5p/5TrVunYoTRrBz8o2N3CPR8MoXV/EnATE1CAhTvF6E
a6YKYdKriY2mAIkbVmZ1ytTovdvLcGGCKb9Mu+PkJT4/Zqlyh3VPWljsX5tspSI8uPWJfNBk4h4F
1hvwq6rIw3VXQEg6Eu0ICR25rXxAhHPsn5ip3WGexnFhxrY3nK9LPOgW/miRtkjZLc8BdvnFIDH1
VnEwThStxvPUVpDL2UD2fqGMtvi3SF/9BElYmJCb/jo4jAhn0l0DHue3TYBOAQZCn9+9XMEzqfrg
YooLGJrOtQLUAaqvpOz7e4hZ7hKOBb28eGHiSl0mzvwCEFVvMeYTb9Ov8FpMVw0RewGo0r2IjtpW
kH6ZgxxNmzufY/Ztf3cu8AZE/KCK2CW0jMVvrvlMxwtI5kzVMQLhagqitBa8NlVKMtEdnTBccln3
4sk45WasaioKr+gqEecYXBhc+PTjIOMYR82KfsAmcgeNMp1biJfyz1M+Dib5OxdHrrZERgKPEcVJ
8Wq2WBVFD0RTv/XmRt1V2o6YCiozpx9oT2k7ljGta0x1JUCsnOIQiGP4asHikjjo6kwqgcgqjma3
ZxX73lGXq3ENIiXN9n9PM7H2ZOzm3nrfx819vQwAGTKCLvlnIhszPblNaesYQoNq53EhQbVJ93oe
iKdSEbmjDOdzDVWkHLzjicVSVfJqzICzGUYthwHMMjLlL/8iy8vzRNeJkHUcSKKIuTZParIxJKxt
w78x+aiY3vv6EFVv+FttmB9+vuWAJavbChbsOHPhFpRKFTNMWyUuaCDBY/QJwKa14g7aPykyOFL6
jhsvoE9yAyFBA+ZjZrJk8W66eu1Z3svP+GbtZkOaNvthXL4DVGSJVfa6aFsVKfZ1CanIQDgf1OpJ
0nUZvgzxfXPgvllFiIFbqABMpTnc6f/gf2vh/U5NXSPTnN/ksEmTRlGVH6obFlcmiY8SXNp4fVyU
GtDW4HMrjU1ZV0R1iFKGBZPY4YHe5K9PoTsO5wrSnPBoNau7xjJ4yeE7/FGt/aERK67nzFxFG4CQ
TBf2QzGD8lpnSDIef0NblkpE8nXxXIn2tVp9K+nxJhFnSUAqpkgmCJwGlzu9UqR/haBXJ3WZFo/f
SvXCaFx1cJFvu9aPkLbdt6PdQhD20xob5QKA5YK0uU4T8IPETe2H2kFLwwQzKU3EiuY4iRTgK5+g
MvUKtluRYkeZmZwiaHgjIcDtVv65xR28xoPD6bMhD84oOlm1xgPAp+Dz8jPw00TQEwM3f+d1dImG
xTsKqXP8V1tCeqEOO6Ix9hgqePvTiEVkpL8SqwWnVYHtdsZE1WXo4ezl/Q+uJFCJM2lS2QJjCeYY
OXm9bCRJGqJ/uWb6RUxeOFt7bF1GjcG7DkNHS05p9YFWBCe4mwgeG/U/39suDhrAC+LHDKX/y2Ea
m9heuo4RCJdm/++dtNMrodgJFBX6hggNeisECsicDyHTqfXRce/xseQKWzuNUMaeiNG/OB3bpNup
f7gFhlE1xmvMMNQ7LpGwXxMAB0wFNFhn4hlLkNMHuBQAi2zJTLHSLAYdfGt0fyJXGKJILyb/AG7Q
heTAizkMk9ueCLXGJ2tG9+YXmQ+QazYeUpYxF3jFHKJNJYTy9Vriz0I6LP8gbDvhOpusVovKTRT7
koGbt3zh3AGNCvSAtxK2vbmOjxFy/DSpW74hcoBGY9H5lqOyJdRjv7F4YQX07Tshri2O3O8CtJQO
CjMYP25sMU2fzhwuJuqb8hksH5CZEh/Ph6iK8JUQykOne+lrOqFGF7gHbiIZ9/3C6i1MBcFFW2Hk
cZx6KDp4ZGwZQm5FLKcZ2OAWWQdOUrTNw5XUUaLIkYreXt+1oK83T88XnwwgTSO2GJqaMKrzobSV
FKryKNdCOx/DUvgRacMFsfmTOBlda8SToyZxwCQWEK5WYXKQcfVFPx74g/635LkeaRPxytaXcTKV
eNaTSm+st81e98WvfQPEEL94bhfRaizgq9f+rIOQ/XxjeAZoX1HWgsieoBW2UFz7czr+oq37NbiM
vyn0N4Ks0gQyeFZBk1/niKVkTJyHz7j9Zn3JfU/zf79/s+EQUYy73ZPH4lpuYdbhbntJzEkT9+u3
ltolbMD78alA2imOEeUQWSH2jrKUiFEbJ4vLzrMZddYwC2A8HIwAE1tQVcf6JX7D/laSxkta3U7q
yFA18UPQwdz7VAvaAfPIBMb1Wr0aW2C7v4gKh7TTnGQ3VP4Na/j4xhjpnZR9cF22lRKL9InAuHBs
uLbEuiAQdXpUXCmehlExq+ECAGFF/ScXXO8VeJKOpkk/GCXg1AMxiGMLXoOhKjmAJ9+7RBEAI3V3
QoRInEIQSC2p1xlyvfzVgxQ6ji7gFQ4Ohnz5kru6amPpnSmabTvrp+XMgbzRAKq7twiJR+5DAuhQ
HwZyBd2Y02h9uQ/oaIciDBdZ6O5W/KV/lpN2PKKCCm2Nm/vAllpuApE6SlYgcGpOmu1rpKwSFJRK
LuiATiG4KW9tSV6qLIa/n4MX6TSQfhfO0BN1Q1aAb0y3HWfWYNNpJTZm8qVZzmXw/w9QHXwYUrzt
CvrsCI5/P78Oan2h0sVCC8rCmnU9jWJnNI++QTIiO5GChHi1S331xrUJdEGBUbeStHv4Vj6niAMn
7xPedaCjnTQKCq10zHpAeHcRWy3hzC4EtvYgxcRJeuAsFrMM+aaSaLX2hCm1NCRhXIiY7n78VPnu
RgfmKLlS/qRWUWdIjqnKuyL6N3SNEiWKxhPg6w9c0UU5T6++zDx+m0cztdpcdbkNySZRuaEhNo7G
7GpNTTMLL3yzMjZw7XXPobdwkFa2L+DHE1CwgWZHNt/USpUI7ZJ2KuN3t73Y6L2+5eAHzAn3FW0f
1FFhA9fgY6o0hzTDwCKwVoeC9zHQ9+woDWSZt4nxhmgH838sNMVqfpUFRY3hO61wCvDh7SRxHgNd
PuzcVDfzQBq/lxDAR3P3I5bgOEmvk27MSN1BAmjoSRgxlSw1mRAgVlUmii9aHE89Sq3wKORHvKWg
SAnwFhNjZFN9oLhfgy47E8xB6oILITaTZE2Lxs0O/yMDaJGN56UXGxPcZQqkKYDZCCyYJVy2NHaK
koi1hZxyVIxk+2VwwZF62r9Cj7oLhiHUi5HN1Gl8JIaiKjh5LHx1pQx2BcXT5MgdyTLfZW+Q7dJZ
6ZAko3oTYMo/OEXdGTLZ2Xd1b+NWiR2PQ87ECfi8DzR+fea9bjuyHqVuDsYd4UotK0THxJT68Imx
pmItmqXxYGp1kDtDp7r+Tkq8Bmf9R+egJ62dlQGb0+D26FQHEkAq6TAJlqoJnDlZO/LyZ1Xy7BD8
KgxChj1nLrE2A4YErqH9LS4RBMWvFRxIQbTwDzvdgr+70iiWmLd3S+BMEXxbPvl7hLqBGfNb4KyQ
KQ6Suqkj5OuJy7+CKCBLEGmHETNbW+hK/9MJJeuinzsSQjqjXxQk9NSHZOtNvugqIyjs2xmgp9Ve
5/Tkj5/LnXLj918DEqbQTG3Mr8rFsRzJDcfjlDkXTA5AvcUs8ELFD82NMbZPRVtmAFFlVA/NdRgb
ZvJAIoOs5qeiQVE88nBNJ2yCHithVi4HDSmAAvY4SrI+3rEOOlkFaMcNTeGOVmDRm5No7sfbMz3W
zlx8p+NxmGwJF8zDvDKHSMiLWWOKEncUyLWUdRjgJYz8kWX0x9qNJRjPtFrIbUzqd+OUwRnyNgyO
SeRCG7ovjV7FRHomAyzc6irf7JZOgEitmjbaGIfbis1MSLNXR92KK3NVlPnehyCEfJQVOXa8pN2o
6DK91sX/zhUi7tgDTnNBWIp4gFXMdtb/7ryHD37di6gDvccErtJiSHYkzdvg/jvll04152pWK6rv
DZ3hmRxYwMeN0tKhJRSYwje4bbwlkci6U0onHR/+AbBw1buaX/uHsVzGRuMaEbnC57oBWwXTw7Ej
Znu15ZiubkoXNrJkQl+fbRy/NOuvbepYqQO5YQPN9n8QJP7hvn2YxWr3EeDK7QIqf7G93k8b2yZa
+EsDkKHX9N2fi9aKHhCr6Q+ClY4gr1H9tt4veNoxE8zg6JrFMOrO46FMcoel+5TblXfj7O3pM2eI
Kj98OXGg1loCxpgpNuZEMa3FquijV2OkipmvDwuzXxUjddjLmV4YTUWmc3THoOV8uJjfKk8OLPRn
xzzN3uGyDi9brbUSJWsVw+6U/7ar8ONEkOiWy37yosPlsQVEXhpLwcqS0nlWULEmcMF6yic7OXBY
kFAbH4oPV3WLWBi2ruCg/25G8v7ps1p49SE5T6WHM5p4pcCEWCH7vKLkKySSyVlSeGF9Df/u39Pc
2dVHU399ZfN7meJnQz/LH8xgyCHdp9YB7w/jqraWPs9c1s87xDsruRdYri30WrOBbstFKl3BWif1
21DSkw1svX1A/FUXTM1Th51GSHU7TkbsKxg86xEdzMCr6inSILQqCu0AVjsqiF2dBVMIKcZ62Pt7
kMndji0q0ZxpiLNgJLVnLVh5scc6hiIOztEsS+h+jkbYKCrUNDlhVk0Z5nK+iONnj3C7eT1B4FtJ
nfixSOZkU2ifCbzxdywA+3tOlnH2dFJ3qK0/REU2rRdr9eOceU9leafGyQgdNZxYAGMsdlu+4bbD
baLG8TiIN6TVsUrB45r6WE1Wac60oajtb1pHxZ1dJNh0CI5V9MkHHDDmVC1NJphmOb2xJ5uCbEi8
sto5j78hJtU/5xLk9Xv9bcsJuO2Hxwf8/Nu10WKldhxJE22c3wu4vHYWZd6Gm29p4djXXE/dncde
qO47/XSFV6ZBhvlwktrCai90CFM8HkDL7SDraNUi900lFW4D87jD9yGgoFQltvR7vqOL5+Ca+T04
HMYCvs1foKkTn3/NDD5FFdaOCgEDAhY3tNdmU4le2IDRiUDNKAnQO42t1XYJWAwba/t4083pVJ+z
jUNySwcTPXUWLQ9+RtbqHwl0i4W7s6lijDoZcmUVsZWX647gCHwjhvnrcTrf3JvjMabMxLKLO6YJ
+3uI4QgltHmE8MCZVUGDEm6MIp11wg5gizwiatMUT944GpNh/Qo4N18YKCyQECYfrEp8oL8MjyT2
BXdRVtS1Yguy4hcVv1V90hLCRURuKBCDJ07q98bDyYbEnX9p2GgWzI2Mm1xE1vCfnSZFqTfgqRIu
nbUGY+01VaVXs5h/8vceOUHPDkl29pmG1uIfPtQRKUKu81j4ha+oMsFG0hBHrRSt6ipdSQphWxV+
qAlkUpQAcqBzz4vs8idLEnUQhaP7vA/xK3HKppTQHbQbY4jIuTnuc9HJp/5qP9OQuUkydv6j1NBu
9cU6Z/F2BdjGUIxLRdZzde89Q8boxSPJk4rlhc/RQSFucjMkx3A/hrrClt67IvoGdGGcyDqeVh+v
fk6AGESanjKPMMhpxoqw2I0FL8nUf6M9kw24nVl0K1X515cwCHYvET5JEYggT0c49fEybaOv0qGf
GEHe3cHDDoe8cQl76xLG6IkCLuX49GzwI4Ph++/7EzvW4TRkEhNhZLuppleMiVNQjb5Litz3Ds+/
l4ho3dy9+BZ08gOnjNh/2uMBSDLhJEn6qyHT9+ZfKOFiGd2pUY90VVjC1xpnUve+VWyHUWJpXdHN
jmPBNwixYz6EFJY3PQWvPXVOqiC4vA/daWaV2GdXKb06F4ea2V/IyVzSZGX1yg3js5e1LSJrvgwt
u8XgC9APdo/+UBKwADyDlf81A0d9pOlhrzXiA9OcuEdYAPXG+z+fH6UPTSXS4G5qN1Xqf/tj/Bxf
wvZ4tOBwJmThkL+myTVfvNtED7J/7vyrxePHd4fGWYwXxZNm/brqMClZNLyEE/4p69YAMW5zQ2Ou
Tx/0/M9MH0fHUnlfwbLwuko32uAzWi26epvWkOPjGrzqSe2Vf864RjlHkrzsfNoDiF9lKHNnCilw
ieRWfDEul2cDOvs2JAmpX9bGTHL0XGN1tEMgm5kApRJEI318D/w73DMErc4sUvw2yC3Oto3r3gnY
9XltJ1JzP52f+KZRjbH7isZqw/zlZ96WGWzGlzV0hkDaWwbNBJd38dmSKJDWbJVMwiLaOu/eEmqs
SmJYL8MVvfd9a+J5MNGmMSyf8cjKI+wEVoLfYRL45kDCsyjg9idv3MS7E3sk15nnT6257F4YJ59R
Pw+WAvgg3QP7QnPKf8l0bIvo3YouTeM9d20f/lObFWE5LzZ4PgPvAtJuhI8qrjkSAq8Nc3xy564M
uNlg63pMwWNEqlmoYsvi6nCIuhNnGbSPN3s0cz73MKMMU5YVYC/aDV/gsLFrXwc8OpNcg/KsZz5n
qbDMCdFqqRkqEYx3rp65+Gk15xL4o3qeZ9HXSPf79+uHY1/W1LMkESPoy0GVYKVPdwbfkQeA5xp5
EPNF7LGxJ8MEPMV/ejRFRbdeQBIlQJjommCEpQJUwnMNj1weX5m88iAVBNFFYQZSrglV5tcHuEzM
34EoeEh3ygt5NhHxraRGi2ULLmaNsZOwa2pr6Ha18ptNr9gD9pGdYObCJDUlVK3cloXqtsm5XI9f
YgnnL6uzOhbeqZX6ZOXmr0UIgKSGqLCwiK/8PDC/C6ze2+O4Kk+CMI2aB7eF8FVu+tGKbHeW8QIA
iy3S8SmDzMCwjQalrIpKhxPJAJPCAeIi6C4uVNtuOLNysuNfF4WKhl4nqqPW77Z2FIoq9AO80cZr
Z+AE8W8dfkyCYk0E2jSDoV7xasEIc15eLiI33/1YsT/tHfmQhSoY+87L3G6AblLfgnMdpLbd8vuO
/SQmlCXSZQJ/lORVkpSfGjzlOKYnoKdQ7oKtw4TkkJx/rqucSaygMkzThPNNOQbjIrfkm0Yjmu5Q
kkf79DdqrtLoIg0nfS8aUef9IflktiBWF4BdZ9aikizYksjbX39dacFdzsgEsGyyVNXkYxZdmZkx
AhK3EG7oYl9gSuzVFIeuruFwY4Mgs5qZJNM73yP6tbVRbWBn5+BHYS6HVXdANPM5qbXJYrVl6pRJ
boXCcG1R0qRyrUl2N8KSGy9PA+UTLc2W1hV3wr2vO5XHbZSW8n0AIe2QfqoArvZ4pz6V/xThSId9
NHs2qCM/fmIeC7rBMlpNcRS17A8lCt2EMem1HlBQQz3L6G02IyWlF/SWzzTqaMEJkK9xDk/+e/Bi
zt+SqpbHYR6hoX8pvDPPrh6H5PYpPBYDq8Ds946EN3QsyS/qwA1pQQV5vqTGsKpDPRqHS3nYSZxE
Xk3mVZm7LBGsdqXalMidReVeEvkmLc0KMHqItz3ft+qggh1EtKnKV+AvrRk6pzqBaGd1DpGE6tTW
sTzYRxMVPamAEOogWwO8HGnfukdobV7xgBd2BL4lY8S/DXezKTm3EeLuRkX/v39rh12tYYFDnP2Z
A6Xwn0Sfl26YRrco4MeVfhB0po9r1R5zj8mbwAZ6SjIpdR2ypu+HQialhD2yRQeNpFmV17Iq2JsA
kcbGBy7secDqIbAoz3x61ps9kzdJw1Tm4ss4HHAimzm66pcP8pSTGTEgdS7bKL3ayYXpx5HAyG1Q
1J9Sq39Uo5pc1LEHbSQ45jNJ4OEwIqO/gjs6KL5wt1aWyrik77poGrCfIyR/P8Si1LEvM5f821HO
4+jorv02shdp3VgZBxU5m5mijl0bgXAJ1zz+fzDxSbDW2U5EVVlDkJDxhvMTxEm2tSdUxeV3bHIb
0yDyxQHdJtGZhzITgG1tmZ3YcMGYLGmU4NsN8zcvUvqQ2Qowyuji6nXn1qlmMAfWTFGkRO9XJgvf
RKu8VuIBjveUmQiu2lH8NogQ8Opc0eG9yvSqdbhBp+TA9Lst7VAwWbPat9IbJTUpIMxRtOM1vpGP
aE0Qu4wa9xoGmJIa2Kl7YrtEjYJIh03YM3FibwQXYuvzlDdbY6uplB/IE5XN3ogkoiLbtsaL4xIp
HyDPGjL5l9WqoYNOvI6sNbrVLu4ULpxxabUwghnQk23WlXAvPNiWWx8OYFOhm/SM1vI5eZDGN2md
xDfMLHDV4QlXW2yTmM1jmYYZjGSVU5JICKPjXI711LId5tLjeGtFcF9rCA9J83rf3s1hhfn982Ip
A6FslxVsdSQztzuOCMLJ0dVmr0kp7yYWMUihDuu9rYaItIfyEyj9fSdfJHPU7m46aPNhmoUDW0ZZ
ziepfo6ayT7s6gJ/pKLvvswTY5UPD5uVIEMhJFtHU7oK3uH6J65AjsYL5wLYl2fnbZaMb3YNDC++
nBKTq9EPCiBr8wAAOmER4YXZy62AzIiyPAVjjy+CIwyw6eN4WPqjZHefGrVz7hKSnP9NnD+pcibV
cppAUmaxPfyNEqZQXoH5lAT8Cw1E7vB5k6vACBN0ltUgso/qcq0ZAqbaWM2niAmWmisLHCkcnwDt
A4TnwBREkNFjtRp0lwOmr4JMtf89ibraXlMOllnRpaE01sZIao7jiR4Z0BHrWE24fw/0WjkMXGWs
EsqooZQogLNvhJX/1QmZEzC8a7WSINczevF4gINvmB1+TXk1v2+WeAczRL6qve/C8H7e0XY3lc7a
bZGTcvrs69/s/xGugXXIt3MXUOsmoLQ21NRrUzowwG7oZFlxRBcRb3oHIP0vKgiT+1EuaoMABYKj
79UJUS2FDTCS+S8BUzR80P8o2M+rRJnnQm2FH2ehriHjypJWAsRuxwA/K7nSCEWqZS2eKPpTm/G7
MP+6JWB/txZfK4s+L3k1WtsQHy8ACtBZPbhqIgUZoEbSinB3H1LmYbQA0HZg73obtRcQaMRe8y3e
0KH1z6am8fQJw1D5t2cBzU2pFWgUu9pMMDDdTcnFN7qn7cISz8+knnCiREoOXZR8OALZrPH7q251
7ERckHLDdQRLZtia7pwQrYgwzf/D7Vl5Bm+ngy2no84f/7yMRPNEIlaH8RnN/nnlqUkI163XyZPX
iYcrGFLvVuIY8RkhJ6hlHuX0zIEyqYD4222CzyfpjLxPm0PSmGgAJEUriJLRn+dA5JNHowZpmNME
g7EF/m3XCwWkyC77FcFcALY5sWJ/mJWheDqkX4RBkRco+TJh7MILbku3jc9JqdS79ax68SiAfq36
wqy5EsHCIf87x99rR307Q9/HVQmwxD0jC3vux67vQZAdDX5SvZfQNownvxvua6dWTjhjmKlGuZkm
wFIptogJAouIMQ1DtjKkw9G+UAYqyP3JdErWI+t+tll0t7PsglvTI1MLYw3L37ogcpfJX2ne+BVF
M0cq3AMOV6Y9RWXbyLgQB3WAYkjAWeANFc00jmeWz3w2kWtnEBJBOx02p8WNXf1qBoPaHPegStWc
9adzP9hNNeRGUP+3SlvMoN9idu4xngwb+Mu1JkKkbqg2Fm6jccxVGst2AwlI0JCt8am5AnOqLo+3
87QZcyeXekq9wiS1uQKHc5rfP/9EksQULVonOSGS/n5L6Z3UZXIc5RMe8NOV1hSmjG8q3gKFlh7Z
WThjhZN6XYV9f8GCCfNeR/C4oOFeUL05a6fksn4JIq+zBnQoHYebFv69FZ5ddm5eogrVjQddODH1
tlEpgChcVsHYE1BPz7qcH36tKRWq0pIz8P49iu0tyaZTwAMfKezH2OIr5Fp2lETtFC92sgtyrf8V
Rb0P2tw6M3wDyQcqoTuRrJvMsKSbPkfAiWguvCMvyIGvt5dT1vfW2+tNknZRHyeJt/usYOaTTIM7
+Rc1LNcrGIuSCWoOzmtXKmtViVP7b1idcxKbJzWbbNWmHkLt1c2OI4CwwmInfb9VcMaXYHVt2L7z
dsg7zqPUMdmfBJaZzFit3kePP40ouoC7rfFEhFSgudj0JupuAunwE8DzRtoyD8OXVp8bpXZyclCp
QvhAlMkGOCZGEpn+hSVYwTlFS9gg+vXl7kOYzuaMcfYGKKZS3ZjTSHUV7JsrAp5pKJTMQfjDleX1
c6BiLk0fLoXjB5/yR+CyU4Gcjgz62sB1n/hrRm4bgxTbmNWO3ip7osOcaF31rTGaR15OQyD9+K5W
Yv7mlJFXGc0clnVB73AKvxf0Y+JhX8mlWDf7N/eIB3o7/VIlCLlbFuBwc8hLS32XrdScnzSzHEdL
gkX1WlgpJtw5V/XmVKD27fMOTREIjC59wFQ1cZlKuUtL1+nhBSW8uW3CUgsNpqTT/VC8YGV4s+EP
FybxYceeS4teimxU95IurZ8wkkwRts5azHjICypQuX0Ahy3t5I1Qkl16To5jp+WJ96gcJNF3xSPI
CK+SW8ljy+WI5BSfMEpCym5mRlyn86V3XbohipcR5OFzK45FXFroZ54CW+tYGqLOUNd39S6zC811
bUDf8pFLqsDVfsrfbp1Sd5Q6UIAr8NKVpfKGrJjM94/c9p7ShCd+jY9CX1fczY4ARNGiagC9PX/k
2HAavDXpLGb09u3b2WwCXRCSKZmAP5ckl08gDOvgAH/9n30OXrz4BSsIOa9gxaPS/4d3Ar5bt+z5
tIRtJGuIsh9AQi1pELoD+GmOG6Ierz2g5cGjOOCO5C5VxEESlX0jJhQZwp0nExp888Hb1s6gFA2y
Hzr7EKBoAOYnyhYpTRcVLwdH6F4tuQbmW6HZXktJxnJkWf7mpZK0J1a+XdWkZf9dBTud0KIqovay
RRiEQWozQb/IPXeO55Hqah11bT2ebcrKWGCNSZukZxiW95dJ4kTweb0jwSU9dfWQJVbNcf/Ouz9I
J4qVn6T/KvZ92QZ3elaiN61TaHOuNVZpsEKFvntu+Vo3BQ0l8tWZ5dh3fptWWrUls7LFRSD9rM+W
RD7NGwGaJXKXb1h5QBdTo+HwpODQ5OO652vNPqfFLMNPgQPnsTV0IcEPkwbO/yhLlWGLTMUTux7a
6cS21AuOAUC2yQjWu07TZy+EnnaSvDT7/az7RmMXfNJYBpTCXsqrmCeoU+MmnngMW2aGpHFJirzd
4d0hZsbT0km5UijEvRyB8kHaz3EGDO1gwt4L/gUygxMlDAGYSZIeZh6Y4o9tMF2VmYrY0f9huHb6
77diHUQfIP7gtboNBrjoKKOazPdJo2JmxiB0G4nhXZJhpXyWgu4FjL5yXcn6gVVVSqVHqGMFxnNs
uJczUIy+2UMSHLViWMEddsvHGj/uI/QqjDS0M0HyyItuu3sTQE72vfsdMgn9sg1QATOAwWC3KDWu
2Ynpnl6OrGvx5STIfYG4IBlbpaGFIOTSW7JSzcDaj1pltOUlB2av1mkznLhlo+cAlK/4fejDQBE1
z7EvywOBhEVMKE6VEl9OnY4vbi8Iu0Nr6iHNMSjf10ug1KU8rd+4Q36Ki6JIFBP0+iz8WlLdNZ5m
AVs1rfwMseudj7ohrbDUft99wqLiwOalZz5owwnwdSQIKcR43OpspcskU2AwTy/ywPF4RTNV3S/g
65p+fqQzPe0z7G+ldv5bGKpzYvFSsYXk5zFHlF9ObfB5E5WoEUQ5lnC75h54lAl4FkwoLJ508mB/
CPF4W3E2WkapA9idPDJh1UmA9FEiScvDrd8tCERlhqNRA2Hi5FGgeg43ZlUXE9h36QpwqJDKu1np
qA0X+Goef1iUWo0y79+HN74Wsqw5Mr2sGm75Ws7lU52FMBZYc+P1fYnUf1Ks6pDb8avUkoi5pNB/
4ueTWKC3V8T4Qu5ijZlOAY7Mpn1qi0UX/FgzVb4Gbq+QGuVKsUHO/OvHkDKShOxIHNvINFrtxMp4
JUTihJlQIDnU9E7qtcvkBqkN0HNkDWQQjP2ZI8BXPxjUq96gJR++arn5fQTR3qrid4uTYozGudql
Ye0ZKJ90itBPD5tvykcCzVC6+Q/EeHqHQgDc+ZdG7YBJIN9iFoe2wlKkLj7FpRZUIus3Fi0hqSpY
Gu2u9h91UaFj9gDvhpI0Qbjb1XAdPF6SkdYx+rjw5uOdoxEtGbcfeTJyn1Dc4ZWjrtcc6hwyiD58
ZYVMkww+w9nUw7DkqpIxiWXv3oKxXtiAzyCveOGs9fwcwGQjC0PpHkb3j3DjeNtF1ntVQJXxSajt
ZVt0s6OPZfNsArNBGtgqMXHE3pQKkbpzwLdj7MOPbY9qU8wEuvFBwIW04+MURiIZPDpJtMvxCknj
RRjE/BmcW/8RSzqGu20jUSlTgQ7eeuaIwqGypnOWwhQy/TNUe9j3YdoxhA7jNk6wmIjN1Wez7UwP
uVPGj/Mil5ipb7MPiFeROO2herJ/XNBiNVmSZh9NdugDYsC8m9pZ5T9sfnCoL4ThoCsNv0e8V//j
nRL0Q3hOXqX3MaT7WOZjmxmQg5iS3XbOgT1fOEVpRKTVO5t1TxDHtT7rlSXz3WCiQr8eNDTYEFqZ
l2o1jfln/VMujcgHjbNm3ZIIcCdMrt0iTf/8+BovwMJnbNErAYJW6maNjyCaINkfd5ihyV1Sdice
Ae1KgwC985JuuuEXxedMrEfifP8A45YSr+7fIMIgOGk6fCACsMVogxKZXRIhfgyQaPIPZK0kcjhB
Ju6FeS3s7/2ueYtmYP0N57NGT2GN/070UQ19Ya8/EtW5rdgbOvUFxdQr5W/U2XTkRm3UZ8++FvrA
VvvbCE3hGP9t2SHSOizqTUdsgNTEu4UaMt4YSojkQiMm9LFEJytzowbLQOxUAgcUa6hP6/dB4OML
PtwvV235NXnu7ApGVmODmXLM6P/6w4TVSzSMu562K+m3WO0NPpHhdRIwZYDBWdJ16M1QlAOaPFap
Jk13iiDKEdQYoH8VGzzllWC02XBUTAytg7dQyO/ExLjXliLHeZz68DP/gfISN1vsrsL5DrQBpMuf
ufKfOeAbJDwuCDB0SVeomzRI2+t5lC3Ros4Q1m/H1dpq9iWoD3fgQ4GAmGTm+EseLZvGrRASV4Sn
ooh7KQZ/M6na0eUuVxfXcXB+Y1LT3NLSGVoNFCACj0nN3mnUhrEBet6nI9SS0JVuNyospkO6w7YU
HtRArS2tO4kEuqVDH96YU3pQALbtyJSkFF60/3k1Yfz6ksjQTxYB6HJCZnbims12th6eHXYpDbGe
RJZs32OEZ/FQXPujPU5X89o4LiBEEnxpYgTF9pfw4WB56eUUH0HI9OhSMKn4fh0oeqB+1n3D2Net
sxjQ/taUCrMWX7FWN4NFTzkpflDL4SncUVn8RXYrgIXzMHUwcr1//C/mtotOiP23Lf9bv3NVC2U+
4AFEcqdmFqyBhSify2mVMrwvDw6Peg+wK2YVO7FcKxcLdi9jhJ8R6GGpHI+gOZGQbJk0fbU3OsYn
j8u/PQUw4hlg+cgYxvPwP8URcJRKazd6MGwPrwfrZ1qaXbIl/zV/63j9vupFSnA/k+drU2Cy/Epz
BshA1H/sGg4+/gZMjMyJa+E9B5Ez7vkRH0RiIENICHYgUUfosbz5vHXpfq91bdFbiUpHiBTZWsBt
PTCjdTId2C0MWZdIflcwd8uWOHKRopU7vl0ZK0OgbRgmgaDiDhZpe/2MT59+oE6BMYLCsU9JV5We
oNeSOWMxOC+hg/Cl4MHFVadMf5xHXKmtsBTXygCebEzbRd7bS7g3kqebKrNyO+X96wlboqVY27nB
DjEpLoBFpkS3o8CZK+i823ZYrJ3wuVoRg0G0xTvWRa6cAxaDhe6e4DG+yhwaljvmXkkT8BukH2k0
46ul0vAtNeXPf8hpMUG6o2WEWrqQ0jxvBLcF95G78VaUKHm03xIacS0YGxFDNFk9oCMU9xr5yQ9l
4kWumN1avSld0cXcLXTU6S8+EDr1s0A79aqUlngOdvi47fz6YgKmPJ28AzhyTMsf3v0+I2s9Ahzf
Pn3OfJdys3PY03EpRVqUHsHkt16KvfgaBotRrTUES4978MWQ2vT4Vm6aRN6m13oSQAcKIVC6sDc8
1tlg14J2HobQQvPoSlJ6JToybQORX95G1LEGOhftGgTSfujJ983kYQxsPQO3JjId7UvUcUNllUX2
8PkXylLhw8z4ksWvEnAHg5VV+y7MC25VKXyQHYgFIZEZO97JXyJWZchBV0SlJQ25th6nAd/+NZu0
0Y1Id0VmRiXy21hYz8aiEwh/1n6DnHeOb1bquFN2FX5pH48SqwmipMI3RMUiP5qlN+l2Jxt48c6i
CmtdsNwRb8aPf1s135qEN0nwL0kKLmGy1gQLmOIa2qM+cSSUMduTN4W0SAaNIS5MwVWAEpBP2Fm9
J7YD/5EhnTr7ptArFn8LrwPuUS4EfER4VRDex0MAGg7zbybBWSNDRcR7xoD8uZP2jQJgsQv+KZVU
xTq02T1CDYjdzmRDh9jDL9B+fom/yPpNhuMs5mAx3JGPU6lXS/1eXToTL91/tumYWIzygE7SZawq
yWh0O0BD8tJzYFAWsYfLRAKemhOCKylgPdej+YIW87Kfq0uaE9nSrR1Fzn5p0o07EW2WWpR0z/Je
SV6sfFjK4UpeoQZ8S3Yq+bxzcKKgWmfPWOtFTldV4/sjBNdyPKZXYsGmU10ny7KsvehgWjp2tXB/
mBbkzv1+zsIQdP5Z5cTt5hpBtKXVx8d/xGB1zMcgET3K1GMVn9hxD1oKkx2+/+vMk8Px/luW2jj/
yrM/rREkCJGQTL9ZQtY4cwGDsMBJe0zxWVn/0hWc177pVI7lW8jxvwW0UPekfJ1nsBjkTj+FLl9Q
e1RZPi/LdNbeGgPlHOkyZa3GLT+6dTRMZOjiDTuQIpdjg4MHVWKhKJ5oweJutpAkPoiCiSdbwFqR
qv8yJvdNBlu2Q6kKSUqR9H26hM4ApCW9NRq5ZDcmeToSIYEN6gAmqP4Y8QvNoRFUVKS9Gjve7Lt7
XYP4E1JkZ2isW77axz+83q6cVwvRepuGfY8kYQvBRWKSBIAFRKr6+Go+wqBU4+1/7whgibqJeo3M
vkX9WuJAGqNCnvzrerRjtEUsRGlGs+lC2VTKrVTurvTkq2gQCcLO5xBTJAMPugFYee0Uc1uyHXCd
hzPqP7wHS0zQHIGzRpfp1Zgn7q7u1MijjctADt/8AxP31MOHBgB6dgVNTUCQ090IqHX49+P7SXaF
ZM3xNl0voSTgCVWNaobzLFrJCPjkpCgXJze6CojjWaqqLvxmDo1aXKqHdhzt6Fbv89FJdO29l2ir
beMGo7QawhjBcS6M+E96X2VLDb0fj1sWvG5JxroqLNpwU4PwYIYqBuoKtvDV2QGrr5QwNtjG6My8
q6LeJj1Kq6RHuEUAVpwu5emBoDoqsC/uNgoHmi/Jm3LkuonirKg9Y7ZfNsVIctDCaz9XEEqAzLaH
5OTVqSm+3JndiC7cpkujqNnx6pc4ozmdm80mgSHHqnrvAwzq+nFXxkNNCSWYc2VXDxvg98rWOLgW
m++b1aqau0jQ9KuXnvjN9VR58GP6fVxG2D7qAS1gI9dL/hLyIRa+az4hlEmMeSry1qSKOsTu1WNf
QrPr46+yZFUz+4iLLI2+5tJZYIk3XloxIpvQOUDau3XpXDO4U3KYHoMGDnkeD1hLAMuFbVBn/QXm
QA5EWhGiWRv7ys7Se3Y0GiKumLgljg6DppiMXJK0rb4ebsynTIbiYG369YvWzU6373N/z4Y/Q6/r
DUIN0rrwJHdBfVjEU2xQe+V7W4t0OdSEUlbl2MDXdGIcoCgRL6rDSYLpIKMJsxY9HgP1fgrJ1pCo
ncUPEA4Oa7NuABh/J7mKUINXbUBmGuDPwlWLECcR2/+VM1u1ZxExvkft8vvv/ACVgBDp3o83ne7c
aCVl+TwoDt7XcLsshy3A9UxSw7OG9H7epzZey+w9gKdM8eDv7nXa0gIT+U35VzXyxhqRAq6zFKew
APIxwhepfb2v+OebZ4jRE3qMYrcTUeFtyAVHtv0IzIhlV8l4/ZwVODPxHDB1c/b9VWcq6ug6ZFFq
vio/qXRJ12bRuSBCk3Nu1IlPb+qA66kGS2bfZzcCBf9bu35IR1WNfPZYG6MMiTuOO+t2coXsYE7+
TOdH4MKIy9I5AJ8S/xvmvpAW44MdSoO1QNrkT8JkIil3PSjrWSz2CeTkX00/rDuvZdwIGm5kbCTU
AuEnL9rbaDSI6/YxmPvs5XdTS2zi1i0LOJISmPaIdcMiZoYvxcBgGFVh5JKXhYOx0wIaCIXKn7L5
cxSXgkUYn+eGrSFWKysgzx0kziyOH5n1i5Iw7vNgFtjYbHI+GQDFD6gyIu/azb+bTBXhC44ouIgY
9KztHzx6Qjj6qevaqSAeE2eJ71ihSQRw79wgt5cLrXz3q92QoFBnZ85E0H09XbNPlvHrFQ/fBQK4
lLqDAOBlbhFc2mtNyWIYJuTkN05jSAr+b2Z8x08JscRP8xfnC0zVXiRIdGFC5KVBMZazJEIdbyaM
iG1uF+iB0ROq++FRX6n17qzMFFFkz4m7w9dHcCwQb0CF+yE+WCwRtDBksBUzI2BNRxDtqyz1X8JH
lbFHQXDqF4Go3PtovrQp04bOqrdTLFBN3TaMxwNLy1tb4Cg4f6+QLq/Ba1g0GQfZwOFE72AvvF7i
vTuGUhHx6+6KfWOi8eQGt8ABaHnZUpp1+i1qA+vXjbxcQoohyRKRuj+f+Cyw9G7GI+CLHePgR31m
XdIMbfK2s5VqjJwmOL5ui2OHY/r1vMEVFBDopCbn9NBUUw+vvZM+7eqP6Yp7qX6gD4x2VsaUrSrh
Cwe4gU39PtXSjBi4Ja/5jMJ6f4Q+yySioQy9YwZozOWMj1X4dEy940LCzgenc+b4iz6JpaRwYGn1
bbyo4ZuM1N0VG7v1yW8lDThMBmxW4JVjBssuRkwGwVjmxBnqb3DBI8IweMpk4MK08w79VSAij47+
DW2KW1kU1OPeLrQnqKLwlknrSjDlIcctMU14+7lIXtC5TbGzW5WAXn0fhaFRgUgBjR/Dd/wbwZOm
Aqbd8D/RRwyEeZWQL9Cd3xQG208cxs3D9QxElEQHCF89pxZxhJU2BZAkPR6Sj/YUTzqCvrmUYX+n
qr59VK3X0Sag18G7I9D/bVYyBxwICifJN7Q//7/RkRVrJVRKnTkSpag4lke2roNAP3HzlbnxryBR
38N08Jb2Il/dqYIXOfVO0G1zucpE/CkOuBvZdga+UqS9t4CBbB/KPQ+y1ErC6s7sfj3cOfgvHt73
2KLHMSLiclje+1uNW5LmxA6S5/ecqw4aitAq8IwlZM/vZ7PNUjA1HWwONxvZvvQQy8dWtQEZtAdO
mXsweuq4US1sgwq4ovO4pvQClRQ2SXnym2VkYOBiW2VH+KRa/bQLWXCuv4RkAU9wBZnSZq69uB3b
7+8eKXRe3ovom5LTRAASc/fzsjSi8W8/H3gPuP0QqNX+Ej6x1L3GnAH+A2xiBO622XWddFWOrghz
UpcaR8juD10CG+E00kK64ktLSnamPrBZ/5Yvmi7dPbfG2JDA8xS58kkY766btUOJ5Vv/ezYig/xJ
5a783MzrdGNNnjzcaNpcyi+0vjxv15PiTw4wL+y9SyzPftpCIMogix8Lt5FqFOIHM1ruT+zb+62S
Zm5kwR0fWlTicAVuZ5K/GBrnvsuWhwxWVBec5RcoMXgfCSHN6dB1verRXzOS0tE1LHtpX6J3NWNG
GKTjL2mo1V80ILBPmwOJhOCGvs4SZKfegnPbQRacmqApT0nrRAcmFZOepHbu5OoaLbTFMXDqSMUj
p5hVdU3g3kYFfhp3dnHq2MLXujGmXkanng+uCNtENY+XdGlc9dD1Sj6EhIL/MdiyT1v8Gsu1DvQ6
d7UV1uVQpzFgMofm+gJmjmB+DWaD95rdjE3Zn8opzB8upIZcyU+kaXnN+mnmsIBpB8bd11qPgFGs
0aSqoqDApRNDNKw0bW/ZTdKntkXg7s401dz3Zh6b+TmTiuizJw/aFRL2YZ6Y3evwe+IMEo3YNLSq
3543jcEuIDpjw2nZMP8bW1+0f+ok+ft8I0crkuMUhbZKbMQjiwqh+JyjqAoPf8zhSeTpNEF2cE7F
z5VvjsnZp6vYowy/q/4w55xaJuspWgiask9ZsptyCJKUnCMxJAKXiEOnQnvCI4j5KgEYl4M48JWA
SkevaYEkCxXha8Ok6Bs6W4aECwFF9bp/yc6Os9hHZgogRM89jrHi8uiKQuO5j7OaUfSEqzpxEgbX
ovgSAlBw+Ulo+yAbXeX8BncFWtlIGprOZ1hEpGY9GuvRMAxtOPNq9AhJNGDzlH0DKB0xKqs6C+ej
2F9MZpkdcBe4dAA/7T87fsifARtVW9zgM0dV4yl1AmvAdKwDGBuDtAjjUsr0bHIy/gdGYvgabIJJ
Xeau8POy+ZfZdeC8FcF81xnpRAdUN7090YZvhLeJQjTQEpqs9JocMQKvp3UcHIVo7EIHHLdcEz+G
L0Ha4CLrHYITOU4pTaFa8IXhr3w/wQ9VBJci5Z9s7nWBvZ+2kksFIBQx6C3SCCuhjkwzEnzfFRkG
ZRHj/7iE/EBMNjTb4Vlig1vki+0z1BvpieX4atxmgKme9xItXcV1/f7gfajvup+KqVwEyu0hjkT0
NXRcyvc0sIEgPN/hdqldcUKNX23t0u89BuU5WN5oTXDPFnA7vXN8Hn4bgOnkM9FFAukWGTxLxBWu
rfmMK3Yy2ei1l6CVMGnvxOZeaX5d7RyZNVx/KimlAqS62bYSbvHqJOCxHOeNncz1ceZ7h1xVbGuc
g39SiYk8v898q6tHkTlQe4BQA+V23bPoCeM3JzOE2mOD6V6460AXG46XWGW5bIgfdBndD66KqkZa
qKOO7NKUKfq9fkf00fWwiQcrWBdcy2W0tcMUgZExLrOY6zlYVUaNLZzMB559rdJtHoaq/zJgl8ei
E3VqKpTQl8x7Bx33Ws0vu+zj/vEq4Q2syJx+PhhslGzgOQX+fcYFBt6JgWS15SdictaobuAV90jl
kJ8Cib/mnV1N8Y8biHUMZXs8/5UxPHadVbZLeYs1EjEurnxobiBOkv8ZSxomKqSH6eK+70pi1L66
GDZWmD+XjEPp80wff3+wjYhndyECYFooWRmGt3TZde25Qd5aPeCwV4BxlVFDSCeUKVPkzqYUfom8
PKDSlGeu4tlXDgTqo15aauRLEC2WMj3XamCBqlt2mSsSF3gk7tWyi6/V58S8UdgiK/Nobe+3klyw
GuYjTtTOgWR1xAYqIRH2lUOKO7xEAPc2BHtszUnF84p/CLDOpykEPuVNOyJQSMbtyebgH5fU7F0z
OBQy4lVHDBNtDhcOmg8w/4nRhNYX2bM54CIcDrjeMIgNSOMCTqgTGrFQaRyP+XlbeaisEpCLi5oh
9k4+GNEGWKfMYYvKHYpUPR3wuOeeIEbXfPLmWVmb0I1RmXJ5MeddJ2TgS4K0FyJGEMnmjn6LFuID
PGpbiEApeAVPSp0g2CVzVtGvIRc93FqsFSqbnxUW9IXCKJwLXRd35I/LHwxsJtekqWG3hNc/RJKE
yHcj5sBop6CYG/eUOrtg6bTB31lydirBBEItkY0mvGW5SkSplKt2/qTE4pvQEs2xaUDZWya+UWpr
lXgsFQKXB4CV2zLvXh9KZITtMfFBryh41E8rcE0APsw4gBP5vziz6ffTWOZNwgPv7kCXR9u6MKoN
99nntZ/XEaA9tFi7Feq/9hLwdGKjFHI+MMFFjr/i4r2eXUhuvnyVZqEaZL9qlHKGoKjLsCfjQcPx
e6Q3bRcA1lxaliRlenpAhWPiDeCdizFgpJx4glQ+qy+xDXuru91LuL7Vv1Q8do+hOgIqRhRJPH+O
FdrEAk7Gu6MjUrxzN1xum7aAglDDjhnSLriZvHf/8QzO9kdbdBgUIsx/JZnjGlKZ6O7vcUF6Wrp9
T8/BCBWomGFU7nhdV75HqB9SHOa/BcJCev1fhiCTrfidD23mTg1VxqubO9ewnzZAsgEiE3YmA1Qa
WMkZXfEXRFHLbOMoT6eiwZ4XvRdUg0ueAMqkKSDFkPcfYdpuF20iu/ijKR8jau9JBZ7VmiSZHDP3
WjwXfHjY0gqWy9f59eYQKkp66yTMV+1nFbbL6ZX6g3dD/x+RvMOuYPmGLXE+fPYGBC/tObvj0e/a
u952p7y8U5pQeeLbhrRqZPrUpbgWUgwwXGcq22iOmoPCcomTcJRMC+g5YU1ywGVsxN3Ojb9fMtKZ
pPrKkRMC7ZPkpYMru4cf98r73vdswrcQQQ80p+agnlq2sVYh/oHDlZXc0uzNUSx9bQWIo9cEGuzU
hYanZDwAJ3Ih+hZHQsxt5LdMc1njLRKcMc2XeJb2qnCeUPahl3YEDeXMmluUtYI+WQIQoA5tvv8/
0twhFFclV894yz8+iUGkXzXQ0o5XT8ZfG2bwKLa8Chk8TSJIDNbPKB2A4upmcwlP1UaD9el9xejK
DFP8ei5h+e8DJD0ajMFFarKO7W4B9Mc6dKXWceGmv5dkJIsGMUCVVZajnGVbIyaf8Wsq/q1CGug9
qPY5roQCoI9SHZ+dEbAlcc698rGGvFAoOXFgwWHqgPD7Wwz1rYJfHN3RR0zHCAScwFtxuM4jVcwJ
kwGEEer2RT7t/1ADkZmz5G/XnBc1KXY5nmQFBOAokfgu06EhJaYqrCWF1xgjoIuEPKnBMzDdr6nT
yJ8lgh4LGmzqdmQd3UQfJR7WttjXQ2wKVkJy6C9yBMDfzlSgUA4DdTUWjf82ScdpLAxRo5TZZBoM
QYamR/mqctOy3zPBKuuOHXR9XN64WVoL/ctE6r4GmMwItMDBfkDazksT+b2Ll4+XYbnIof62Jpa6
pdaBBSWXULCf8eyWGGZh4vMlXItARTkF+Vf2NZVuPSTZxZxtihUiQFHJifZmMbEWlNkf8ZLtBvb5
M6nkp0CXt3yUJplLHjAfbVwY+WpDHibIZeB7PoCOg1+FlUPKILbEN3dnA2z05eDIIfD8mo5TyG+Y
dioo3yzSyMRci3srhLW0EU+9zOC+o+gzNdmI4Zbn1fHTyajJrL4/G8DTyaz0YRl0Q0xbx9qEzzPi
iLryqQc6CLgyBKkVNDRBcxKRjAKOOGkBCQcoGZ2wOSLZtze0rHNg/7LoLrlO0ES+bT8ZxAUnP2tb
0Ar5ROCxcSmlI8uc2qFZWo+DlijTkBlkld+hgZeRw1FSJweV0lFWc67EgoWp6n56mjcoEyKM0UcB
DFuiNCaa6AVpCAEQYbsXV9eNoYS8Cq+DbWZuIXNNF+YeFoA/tx8ce2/LvmGuZ6comBKnlADKjgdD
TR/COgIhlfrfD1EkqhqvNXLgxpi2vbU6gl5c9XDGzcqI0eXq3I1qjP2w/4yZcpBjJhbG/NbgiVkH
pEvkHCJlBEfG37M2h9Fiw0mTW36fvCKb2l4HmsTVm5K4AzNzpKWOQ1dAdWQsXr4VUtb5X91cTcbf
q3VlujzVlBAv4yWmEf5BA97FKX/76vFUgoRJJe5Kh0RtBu+EYxEGpY1x7edTytWQ8A+kvmR6qN17
8JC+vz9gmwvEV78U2Gn4VBaT2LsnN4OkEHHYWJSnBWbW2mPtcsfHIaXgYzxhPTuPsN82Knse1I2U
jkAKVMW6DlWaVdI53KjNIptjHk2r3i+r1pXE0JRMlXK5b4BwIcac/wiqHBq45Q4KldhYi5jF3qKf
rjKHCFY11R6HPI7geSg7hHHRvRR3CCxK2dkTaxcRegkR1y3vMHtPWph2LxgwRKdPb4bZ5UnpIa9s
V3jhGbCYpo+1TwAiyMXrXLB3hass4AxLO4kzdeIer4rGZjVtLNGaF+hjf+rNlMWhAiJKnrplf4RQ
P76zBOEmUHacxXCOwJJO7rva90dGLASip3von6rxE0LbT4v3fSPSw0TW6SDVCSr3D3eSJ5zNTENm
GC1Doby6bNaBJLuLorudEK4k6fs5Uob/zr29g80GZS/HfPQs5qbaRStICzWJMU+Cma1uOCVSQvm3
jlksWB7c0Aj5e91xYBMg1w8xGNUHDVHoCe+UFt1VHKmlyzDqxLf9nTh+DSlz6gKemvcWvCieKM7z
wfA2aWqmQ5l5qwA2YLraD0kE2CU/+KZlODiMGkVboLTNkoTvPwH+rAR2tFgc94PHIti2DvxDdkqi
W1QprR4JrtHLCBl27hw1Y0xabjwZ5D6RpWa0ddeJbNHTTIr+jVnO/z9lQv0cLeNGCE8NQnEehO2u
dIlPtxJBg/OPTYR+AKAOVVS+m6P63lOou+7aI8CnBCaBMEf/V04Fd7gd2mOJEbFZCIgovmlWW/v2
CdkWeib4k19hh/cOGkA+QwpEQqnVczM+iIiNqiBKxFx1c/PjcYLVhFk6fTyebgjEQqgCwqflv8rx
VxGmZHjjtrUmeq2C7IfLiWYN8WdHBg/5DwVv3mKtgFEjbqo5L9HS5tVXjg5GH3Q2yppxWIJTuIl+
aHittwG5CkrnegpydLrwCL/lEQOXt+7cmchqzYqwAe/lb5jSew27eW3CVhIsB1aJ4eTGW4IwTTLP
lHSyF0p6BSHgOExzlai6LmyqUXbas48QFVafTCPWtqi8q+WCGPcmvq70IjnpfMxWuxorLTg97r+I
SZKLijQ1NTKzEl7Ak09Fa0qI+WSlyOc3k+ZfoomFBM+8kJRWsGqc2HmCcj2ijv9veL4qPqceOb5D
gZtOcNsD7BZT3vnr3VIzcIe1TdhtH2t15yQOPPTaCKTwhGMqnxaJU/Wki5ygHV5JMDXRFRxc5xsf
30xiMNW6erwgyzitPBl22DJoWDHTGnOJUVcJSe/4qZdep8XNzOA3vtbrYVGeNRIwJbjgYnnLO+Gz
q7Pb0A0tqzxQPCID2E2Giyc2Nl0KsdB0cqhdqviSDqzKJw6HsiBNJ4Qswa29XGQAKCT7s84zzzXi
QRxSzaYPt06agekS/jKGqc8PWs+Asj3MuRHD6iO1ZwjZCfpahzt6E4vdCxciAGGFx5CR6X16vEqn
Rtxt7sDbBUST5V2CsNTZrRrNVjgeLuoIvK+XADrYvMwcYx8SZKLkHO3duDmPqfyIf5xbHujI93+v
goHZV4gGKC9ddEiqVUqmriUdfYV+Z4/LOl+Rl8eGQ3KDYJxDkS2N7LxqrR9bqFOqS0ZTECl2T6Yr
asX0D/Otc/KEU+IoOzK7/tUmUNdlgNOLkXomYLlvA/pSSFcCim8wQsknRxLpff78QkFl83jRWGIV
HmCXqfap/WLHCm9Y+WsWWPuz0gZfrNfBwWgS5QwdWNWTVOx9nWOZGlBhYr7eQUgySkOGnSaWNegh
OiIbBCYvAky68WJnARUwX6/BpWQ5QJkeMLaCqUOsiz2ZpO1iKVzKpyQoTYPMjB6d/ovAyCR9LZYb
lI0oyzCGm/6LGQE21dX+vW1sA9op5M1qFGzQJD8iVQhUPnPXZOt/g9MgKIhMV0Rb2wJ4EttVnK2/
V2dO4vsSoUwDar6AiJA+ycsCspgqKRVySUm73yHRdi1W2NPLgWGRH0881fX6+h8nAwuCj6IazSYd
HEduu+XiaQbHg+6FFg/INvgUDKmL6iQRdvkgmsh8oDdJktXB56vStidxcfy/BaHOkIe8aZUoNhqi
N/m2beiPvNZXjHAwJD1YoJUlqJf1+tGMjUwLMODk4f1f8JbLHpK90zf7FYczeWgAcKWloICDfeGS
J9BgDMiBi0ED3AyljSUOsl9NSZbt4NbbaCUzXTrIz9GFxKE5RGMFYh+KmbOIfMdELMozvUV9Rhya
FLNQj5ozS/6jngHoAD7fSCD5jlNV0+Jo2qZHACgavxQDR3DW8bjb0OY6y4GsL5k31WMg+MR1TMfK
5TMfzRldEYn8Kb1v6JYNUK8wkR6hyjxbGmzZ1NqUvq3s22PfVFXLacOzoEVEg+MKBNRhS/w0nEQH
IJU55q56qQl7p/Ho9hcjx00XE/gcAV8otV3+86AVRfmae9qBJdc9M4ahY2Az1vcbnW4eN+lasjXA
m56d0mteqNXwu1iCFw53UAwsz+jLEHKOLHE6dS7OLwsxuwfjvUhFJDiGtb3q267SAraDl2QFghdn
si2RyIJbJcJhzyVQco9fQLgZZxAZr1e4vNeYY0fHecl7aoAf9Dqla+wcfImYd7Ab4AsVIxGJ8+L3
Jqj0iHHQa+EA3fz1A8V7LIsSfoUXHoJPgXoQKndriu/6XMnjHqRoszgIfdVcA8oBi/0ubOZG5rZ2
5vx3AIJWjlRp51tPPb8UwYdRSWBvA9SCAOdIqYFJIFF2nV3vmVvnuuvOzqZwp0gAe3My03uJazvp
hc5BoYy2S/eCmBxSI/YDloZBlS0yEoTrpW4PF7v0ZJNdX3U2mcuG5YaOdSYc8rAE4tgnN310cGjM
vN+Yr9Lrkjg5+1/QkUE2kqDEom9CWjC+jIbdvwEyNy3LBPbkzof3SBkIoIPu9fXsUhmSOzmZQeU1
AGyp1YDqTiQt3ACJtZBDn/+nDWqf5fN40REcQ2yDcNW/EDmgi5g9Z1glbG82mRqZZP9M/SWSILL0
4QFhGx2loN8e2trxxNdCY3YXvMP/QAsd5iLK1BnBvnicXCwm1S4h6sOycK5wHkz7EnveI/DlqGHa
NtA9SiXcVkBMsCjBLyWV8tGQr7Anjp7vWxuQJTUPDy8ddR7AeJEm+intpusqbHRqdppBz9nW/8YD
Q2qMMTidWQD1Rjutu0S323J9d6RcI7sbh0BN5OW4erGxOqL7paR8qrV+AP/GrZwCSx454UANQrbD
meuLMlsFWbghuzcUr3Z1XHqu4V8ULdcM0l2YN60WbdmZlSwcC6Xz8TioJ2fqzP68Nuqwj5GGN7tk
MuCqfIe8ZX4zblr0Z16NPhAhlrmxpdAc5bcCb7ovc/HNxdXzIk2656tjTMgZpOFPdAcWqCFkeMNG
nq0RPlZzfo2AoXkhE0b+aG3QfvYUwJmXqaU2V3V7Bc2EM5xEhP6d8wF4+0j2u2AhZ+elJSVBr+rS
De84gcvpszY8GNdfdN8O/m/U8pJN/m6+VpNVtFj8qGqnLL4/bSrxRFRxP/6epGXPVJXj7UnLhpaT
CNyDdVafArNIKvKPI4wrNN43L9xeW+H0QovBWq8zzJ8QFM+lFa+y3B5oI3072TRPGV+6ncxChwA1
mN+xdIIw7t8SjuF+epVE1uvmyd2FDq54ulzyFm+XmcTfDHhFUIXrz3WyEByGyzi/DXVzr3mUoff3
L5TS8tPgVV/b5OwczAzL25HPhwA71ABIdYpQftxXhxTS3fvH/qOx3SF9eaBSFoR2CYhkLjzQinDK
oYtwxDWPyfIJFRYj8kzbyu6Wp35F/oVIlTaZeowKYpSqZcwLV9Y8XoXJEB6GICHpITlEe1WFwoYU
8V02tn95WWBIPRrKy1hHqqUqPx7cNm+JbCcj5iRa7efiALKoY2BE840CHGL7gIkuTZbjkUygwR8T
DzCgZmbKTR7G7kpYCcOc9/zFJ9eni7GXLtDSfp1CUc0OpUZRPTKj5Vf45nmHs/neEhvqA3doYlGx
boya4uEWYV84mQzhRDjd1HtSFS1toZ1rtjyfr0isACFOa1Yrai3bV+DpGEBMV56dZZSe7HuO7EeE
1P4xpteR9nGvCRRsE7mzx3PblXRETgrr31Wu4OPcAdloED2k2p1KzlSCt/ChIPD4Kz0Ma4oYVM1h
l7HwSaQdUEMTSItuxDD/cfIoD+Poq9DiQFpAO95ayyIXDmGSkF9JgcLMlRgGoOmkcVo0mHAzy9o4
TJsOTl5s9rRBf+tmFaHzbpQ9YotycNs02EhDM79U2/egwRLeqcLEsuGWg9iv8eV+ccSNuemP7siX
Dv2M6p2IP8JF3pwcEU4B4CNPsqy1f2cT+epygF9xeN9N0s+OU2Gm87iIBkH8y3xMwZSoNORbH2ld
tMY0RGAS/7xEE6htbCbf22QNDuCuA8LbZTw25DT9h/wgkyO17PUY6Kc+u7f3+vFCtuTcBiPkG4AV
JGVU8q0gt18BNGQiMBKw86BckqA2OJibhHN7/mEbCgazJFSImRwV+ZDIjdnXVGaorcFxwswmkpnv
YejJb/7UaFRBzq70oFCK7O7DEBt+bNtiLVe+awv42Bc6v6sl6cTG/sPtPhcvWyQLpzqqpT7Wawu/
yYDdHNvce09lHkLzzSK6U3d6TyDXVec0iWF62XHdBYMZoYi2X4LXZ1YQytPtvNVw7m+1qRT6mwMy
3Lt2VwMNGjQSqw3oNdI+LVQq+eCY8mTS33UgQWlp38Py7v03m3q8YVrAGU2BMLPsiVldCCN4A4bl
KtL/8lgLefeC2Syr6klLV+dU09GzhJgkuqfNfS2Rm1BD58jLwuzD0Zwi0zKYKleyR6ndwFqehZ0p
B3zOMKxuRQZuMf6DpWKMBbJGl8+VnTq67XpPdj1psl63V9WvWS4tRorDjPndrIPbjCNY4JIjfju7
0210ey7mziy/UStkk07IBaGSLRRxtHJJl2wiIoxU9pfHSsfuy/u4XRC7nvJeePc6SShx5ZtW4513
Ht+ERYuQu/wqnNIAN7yjQYsQmPUAAmvg1FxLo6r2KFpFU3zFpStuiRggoprwensFtIfE4CGlNIN+
TRU2SI68SKalUiQLOI1vj6RjgmcIwUIIWP1E/rDH7W9zVgJLvQzbRoyAyreULfaaKzz5hGkilWK8
mgwp+ci6wwN3ookuAoVOCtO38Cpy3wWjshy1uQWzpI+N+zEZBMcIR5vFki5bK3qCrJR/o04MC8C7
ewAnGCwyYKRLBRBDWJo16tnmb2fugiWtlZjgmQ/fmr5dvnS31WH4TUnhnh6zhJT8L849MJ0Ou2Ui
A6SpVjn+F54gOLfZbi4PI3FLOCsFrPDxnsLU4VLlry+pTiBopf+2rr3XHY9kikCJartpmfXhAs76
achbbuG2EV7RcJNShCYbrd0ozwRj8EFpp8bHdymQqQ92V5iuFx9v3Li8bqXvqESGZV98Xd6bGyIJ
KCTsoz5XPRn8z/46pyeIgz+BTkLwIze6f1IQakMmMtr86oHkAcnweuEd8UFDtKlt19c1mP/pdo/j
/ldb0YZ9gPaY63zg5uC/3Mnl1fBk3VVtYuVQp7Wnevk8SFw/54YQs9yMxJPJklaPcMvdV03x4f2S
DUErO60NNzJnIrPhcUZlnTq8Qnz66lnh3yOcRMj0dsPIB16etkf6LqfY2V4mdcnpsfiRRv59p5sA
PXeISDqsBPwErrZjezEtmnTlqr2NsF7bsEhIuR/Un8gpp146d2qfb8ph6GnDLiZbcKtANudFhu8L
qyVvIfQvsg4xEGQWqAakjNOFmAWddktEqheaay2n2eo3qEkPSAtqoi7vdNExTKWaebbtEvoZyVM2
2HYfMUUrCMFUxHXXDBbQn8fl1W2Nm21/X3cBdqvj778VKWZI+qRjP7BN7WT0dIIJvNEXQ8pwucJs
nDSpsD+vAo5d00rXXfIwWZxB+rKnr+4ZZ1fwvSXMl13a4FY0+jDAfZ0DrvdVM6c3eOhA+KZ2roHa
h0e1qqw7xEarCCiHWUy/cXVPgKREsCxhAmpFPxHd1/9BlHj7ITFJT0S+Ej7xlqzhnF/jTpVzfuIX
NVyEfPQmaGv8Kr81NnWQG1FuKyVK2jBIXSh6NT++DrwJe1omyUoJK5YSqk5l2V1T41Q/PMkXhaaG
hyGGsq7RxUGqDKo4Pxb7AwKMAFUCAn9UqfI0qeGt8V1S2zxrYLOVTyqQyBXlJpdZl4jZXTcOJOET
Fgd0KYS7fDqzBvsEVvXRzk7RWLOzYCZQuB6SO7x9zIr7RTf1UfD6sdZ9G1i8UNOVm3KifyGwqevx
ufOUfWJz36yKsJjhxB/RS4aZJODmzWx1lw+muhthN2GnOJ2b9qaCqXvwLo2+vH9s8oLsqtto3Wuv
Y+jUaBSKU3dl+N2JE11F3IJXvgtVPk5xPnIz/MB2/QoXZWUD0cRlVNeTWCEQloC79uDYbcKUwQ4t
xaBVPTFqgOZ3jALhvlaDzVDEokqIo1hm+6Ebe8QfPsuKlOS3lWoDgQtFhFDmR0e8FNe5ZgEHdtRU
f664mkdZGu8WFCgGXFBkDqjE2Dg0sfhwE2fWuTZ10sBSwec/1y6jyJRkXJdtjTbsCTz1tEZwnmYh
DHvPqq5FNdApqBZIEl5O+L6yFKea1gxVQo5w+JD7MV0idDK3QG3MQUSx/nSqUsX7/l7t1wUuoPQA
5j6R5pibCwZI13VuplkttR6UQ5VijFiGKcvKvP0L9GZgnHmWXGp53eILm/8TC4hvhMpVRkNFZopR
HBjuBcYFM2h6RTWRVmCEXu0s/5gPwbl+qtazjUDMOCD9vFfQsDArzh1M+CbBrfQ6+ESXu3ApgM2A
q0dqjyM2kdzwzdAq5h5DY6v+D39U7OQ98fh1/pQzga2HeN8VByKr7d4j8og2CfB2MvNOzt83r5B3
q6xRPtKuA56OgVzcYh+VVTBUY/d0BtaQ+9qXM4ojP23/uOMsSCW9nTcxGK1KV7UJR7F2ZvK7KPa7
ZTGDHi/4iQGEgB22A6AsEPSLLtqlKEGWEizWXUTeTrxja6/LNQD7V2ZzOtHICdcO0sStRwXuXRks
Im+afqGKkca95Xpy4iDuYBzRDHlNGVgvhpN77C4uBwXfDhDbJQ/xVuxT0lwyVQd1TuktLCZn9kYu
XaSAKbbBITBrOCZMH2z2+hbN48jxo28yKoi1uoK+U6Nr2t7hxzmF5EkEQSEax21nRsDWSIkADU4F
KCmRTw+g6Jc7sj8W2tGA20igNoiXOsvxVn8NionWCIQcF9Geo+FB9my5TLjp4CwqTyJdV+Fr1GmI
/9htd0lIAKxewQcKW2fqgMMt/qEHGXpfLsDkjkKoy1Sq4w6EnpLAcpNrnS/V++EUde4STGv633TB
JEmvXy9+cfvsy2QxogtQ6xLzZGguZ5uBEiNxFBwrSHXivpcLMAMmsHwUrwgYMu0foquA8eS4fnNw
jMe5o3CVPmFuMlgcOv0Ew4WzgC9c4OCkLztiu5R4SpH+zn4oyAfp+4lRN7tAlKQMEuv798DJGRru
m7K4b03cQDBr0gbVsnGwIJ9ftbDnFr0M1nAp7QLAZlAVN3ZZubM3AublKs15ip5H3XKF+DrUiXke
AJhPheVlrtTrQ7UD8lpccYMTIERhNPJFHrv/c2k+P5MUkA+5cYm/CUk8IY4OgADPzX6h/dQo24tQ
/l6CNlPFo4+RtesmQQPNyA2uXvg6SjE8D6KRr4oTJFc5Bl9Eq7Za60lRlho6EOv+SkqyV0xLe6yn
YQkprEhQ/N1TiR3XiDoL+jnh/OEpnBMa07HLVnMqJC0buFLYd0yx9KilaB4B6EdoXEGuPSH/qSBT
NGWwof5aUfyS7tcH/D2umcUVkIEYpKMNU+Z2sLtvZvb2qstFDQffUVOFZbL7qIu1O7JMadxzqpne
guTEEDSJyevyzNeWGNyzyViB6Y0QML3pv4o9kjRxGUP0og66dfg0P2yO2brHfGD5es7aHTxm+W84
3OG4XQxKIS/sO4m1OQYGnLA7YcjAibaWe0ivSoRpagFoL3Va0ky2tJpJZStaHHiUNUnLCjMjpRJZ
94bBXzOAEqyJ1/ohTAP7ydamh6JN+chZaaP5T3UQRBiid50coPJ/LHNZ3FRZE4opq3qHGb9R2Op6
tcXAPw0RAau9roSiwczJCQQUvJIjRE3KRwbojitCjYqSvxbxx2bFKSjK6kFMoq+UTdig71XimI4X
UkOQ3cHD9JNFnzxw+6PmgbwEi7xfPVg98/LABf+rXpSJ7HXz+VkbKh+jNxxfhY7NPhKC0ygRXlHC
pYWdNcVECFdFL1EYwq+ipXpyZuBjd0/rrEUSPYNN0vWxcW6RhcRCbOPZOTVcF8cXgUZ5e7lNcko+
AAAz3sFj0yYbKzfTvEA6tw0XEDkm2fDX7CMIl2vjrUUw029mluRTq39Ay11Cky0AAYjl5DCIU7rD
S4hzORzpXTF2NR8ScTy5AlrLGiMhkEMhxBO4RameqIcum3FeM1xD3p7O/da2Xq8eddYWTlQXXRfr
S3xS3IJZuqte0ja8/dOn8lKGeCbvwm9Ne8rTedl1Pfn+JUasRf9CLHCFBRg1zjQzI0msq6r0UTpS
dZApasJuBZ/3bFwqpPg5WH7itsTSPD3Cg2IcJ/n1NHQAiZXTsuY3//pfPUcNnW13h2zQtzCzsVOd
ucU3U1wMhCwcDhDJfK8mt82UPoIJU6dGDsjNhUjrSRiWSHppuqFVYqjHLTQJIQFaWGFQLAPLDHqL
qsatc8vn3UWG1JfUoUXdwHfaHwWXNYU/aqglq6cPMvFft1GMcGqczw89VpZbFAElJrOUoOLC/l5M
OSc9JBGdpXPUOsLL8FSd01zeMut0ZoGFeL3d+6hbWZsdMxXeWTwbKXhYjsCCF0LnFt9dvL1lOAg3
zdHFUoK07voXJ2pQtrfK5LtWN3nU5353D5YLEVK8rF3zfwl6ArpcC3YcASsKC5fU4GmaD8CL3Qgl
v+AOYnb/tsIdFzeIXFSBGnJ6AEicCAz/hjX1Wxk8hjuPgt+nhpEC4J8VGkFDOKauZHnYo0wewKRr
v3cmmWmEVnHK23qMrW5HVo0UhkimKmgAOQj/slyvVN6LVSQMy2IsSf69sMokFIMLYK+zFWa5LXfd
zdX3C+dfyw8Zg2bhg2h+0h0IJ4TRCpzCFsQaEpEW/sIUq1s1Wl9Zw5WUFvxdDTG16pTdQctHyqvI
m1BnoDjcKXgSQcpUmTBDJQneasPzABsrGtD2LLCEt+VCNAMQfRHm3g7wAHpEyglRDfegkFHvMyZv
0GsJlPsrV2LNcsk8PqwC4FYI2sh6D4q5byFv4iOnLDGvKCvMmYa9n9BmCkf0W6V27iXudhoas/0I
/RM0zDihXCbVltUW+i9fgYw23tSM7Wux8jjxUt4eP/I8pL3SpJfwfQbrTnYlqN9c0bxfNFwy/DId
lNTmybmoOp3B9Dm3gyCPSSxnHGhTl02uGO8BRD8lyD+/jCm6T6bAfG6zW2v4VNz2uP97B5Z1VQqd
llrMC1ko+26d0CxCDeRI0gNGV81UH0XK6qnvRDjRXFvkCAjCGpAqfMSy/oLmk/IDT8s+BayJrUU3
lgvQNmcbThIVt2hAXJtBI12IdI22UFPvFGUHdz0EYGkYri6Ku332mdgaPdww3uHJpCLxCqqOR85o
HgGYPfo5I7sBhmCS4q5KGDRLnsGLJ51oB7wSZtJSsiX027vZ2hl8Ty1VRiBamoWv137XL87IrZmY
oCuEpRfs6lr7CD/CF+tIPziQJPRBGbRmKroUVeukqT3sPiPrSG7lu5YVZjzSKV95g3UR91VVOAP/
LEwZOkPQ2p5z7nZWDAA0fK3dgmhATNof1dtfR90fKwjZkcTYJCOLTQEIAFgnU5vsCylWjTea08zI
eYXOVahFHRuta/JM2S4c0XQtTWqHuStCoggP7GlCQ9GMzhAtl7kxhgY5LIKmxPEkv+tdrUujE5hA
Po5x5uS0tXAvFZCN7ckd2rjiSw16Ccqgw38pnqXDuzV4rfL6QWNMzhtUjJaPLscpTrGQFugt+iNK
5zilWaWp1ctNcOjJQSpClMe0VlWgH3TQBEo6qWQdDmtNN0MO4R0DoVFE/QrVDFKtEV1avubFqBpK
YVVZznCfO30ZIBg9UUDRpyVVR+mToz+ilSH5g5W0O3TD2fgEzUeuVYG6zrw/UKCCOc43PRYOvkWB
kZUbRgkmfAzZ67jaTBAiFDI5T8HPNzdASUYjps6qf1cSWhxk5O1ZyCVe/mzkcCQcMLx+foJrrnZj
XLlJUjDLuFRaY5uR++h7EyBv+dhWH6tHaXPnoZIlbuZvAz7k0SjB/p8ujdq5Kw9gN1uftxeWxk6b
xVyh1Wyu5Eu0Y8XSgIYPLze1bZJkYiHv+3PtwRG9zjcik5FBbEatIes4hgx+w49IcoMNfqQEJBn6
zoGDvoVmHzXemvbgPIF/woyWACaNKDCNwCsXtKWj9UbGSHQ+t4uZ78v7yGXXMo9GPUcnQCfEpAwu
FL8Sx0AooSbG+SmPrj6vDVjwqVcxTCQm7L0mYgqR2AFgbmI0CZRdei5cUhcUU4folsGbsRdV86kG
Gq1uQls1YWX+P1vR2xsZKJOGUm46bMaIn7oXImQwQ5RONAv3FeV9iVNKOfFLFu5IxDd6HUTD1g7g
TzIfAFAllteBePVx3d0GEdfDhma471wJTP+/cOO7mGijKC9BUeGyqEtcMJZQxEe4xaye9sm3UI+A
lqdY8NS5OEZcbz5t0ZjIp798y+agvatiL8TMCCFCnKlpSdHawlF/MvG1Sa8Wq2um9prIsBHh/zb9
fbcTnhmxIsved0UUBqUdfL3Vo5QQmCtV/aIig5/ovzyhiaDq+jfQ63w1bJb+DmqIK9iVl8htoG5N
vYFhVXgW1UTyazwkcPZ4VDcM2AlkulX+UoKRCVU6pHZejVnh/OOIW8yUlJS8hnFAUZaAxm3pkxV0
/uB7dXPyGn9HteGh5ZVbvk4zVRi2Ksx4iSt1A2P2Zvuf5vUPZLMA48Z58yOoE7Zct6BphE1Siydh
5i92uVxYmsptr7HHHm0k3DyPKOBa64xLJWYL1eIKIlOERZLbk1+Ry4v30G9dyxz8n57UxROnNs+f
iHHS0iPqd8MfROt9AAXDjafj6yAU3qxIMc0m9TRbUSkBHseOptqbsvL+UjmMSJ7Bude1FIoi9R2J
7Ism5eliGWYPRasetXabIyyp+YBxPuUAGJVU8thTfaU/ywJjBNdgsh1gL3ZpnzVx6ttGuv0FB7Gf
s5OpngGCnhO+Aymws05er8DYglnso1RedHxU0UDBabYWLoU2nck7t2yGIkQ411X/VAikZquir17O
A3pz/LeBLk10rSsnn0ncXGVqMvMpOhq3C8Qxvs9ZU0PpXdD17jBy6fQWwwuj/g2V12YM/4M+ZCxu
UFnn3HoBxBs/hvV8mCsTffaf5Ia/FFxP/GFEoWueuyrvNo/ausIhZ7svPJXLtGNgSraxIc00/r7p
wjDJBK6Tf3osD53Top1h6qT+057PesKNgW2euee+gMCoGcOWkgffVHD/0BmXsCHwjNkZNSqnHFx6
UW0uZcFZ5/cDQTWtPzg3UFwyrE1at2aifgrp/3EB28JzMBHMesscUccDHo0IAPsbwu5dl/dP8puL
/zWx6UyAablLuiDPPEfQ9e6ppiWbU7MOCBRY/auokAW53kupqVKtqPI6E+dQZuNFbQ0d0D6jkOab
ep3D44r/FsHft0L29nXu9W0tFi2XZbUtOHO6KLRTru4tjvfqq/59Nk1WwAEmAMnyPKNwBH8dCvzg
X7i75I6uwaJvke/m8LkDTDvWwW+Z2jkNbIa0YWVrmTd0aIJSRgcC0m5co6/XxCz4fJVH57lRu73w
R/csxF+MZptpU6mo84N80lBUc/K38qDW+nElSHHIFxFe5ePm8+1XGjuForZT0Qqw7gSHQOP4XNA2
+ULuOJUaUBd6zYCio/sPNQuQrt2iEjfv+1sFs5/jXDXyZCACtFCu8kD+YOTxIca9YyM5Me9+akZS
edBcv8mCe2y1nnbFQBQA79EYsnOLajYtAXMMpNnKZBkpaOT8b9ufk5vNOtt7mKBp75KtOZj3wOU0
T7ofAE3Koskyc2UEccEGYie5O6s4iGbKw8eKxioz9/ORvUob4hWzLC9pfvdB7KmsW4HT6uQKZxLK
Q/f43w1A9wDHJ0aCMlqRwE6cBIj2VC55q2S7A3P8/J/KBYQbijh7dXcB1cOwBV05L+9RZmnhZzWI
+STGXOQ3cl6zsJi7lLbZzI5HP69BtB2MxYqoEe1+eOD2XucRhCf4SDjzFGg+CHy6ZmTphT0XJqvv
ls6MJqr2Cf6s9kJmEMeW3qoWfXEh1gZEoq/duuUo5eyADCNI8SXT59MStU2LqxRnv8enK/7ysHd8
j/5pd5YDEbx8qxZqbWkdFho/ObormqdyAF52Occ3HDlJB5PgnCSHtCaWNpqfSqHA0cjhs7LTPGfy
KrVJKeyzO+s3lB7BAuoHy4dYQMzyaYkpf+njGwM/QRUOeUaFy1LPKWjGnqQEPou8e9KMe2VTyXXG
RdXmLV/vlQgwxwJlcB4egIsxx2RGdayN4k0hdSxA/x/PVnKpQc1dTCNEwLXqiaHhl1NxJRY5nn3K
esrIA6rf2uDpEBldPj2k6ZZOu0sfyNlMIoq+GHfPCga91xfk2rWF8dHjGDQUuVL+GGz5I0LcWvCN
7hs47FkDPxbFo0d+/5I8SMiB5bdUFQSZh/4AfkZfPlFccChR2soZ0t/vMBoFAYOEUiw+f6mBdoCT
4dMro85IwIOPKZxGtV9bMFYrxYduLiKDB0RP3ZyBOrHUMruMjgUZuuNPM4IwoxfWOJFqZ3Ujazlk
CwhKZRLDFpI5cbThmHTR1rOD0JXKR74TBaF4BifG19p4wKDS8iCeW6dS6JejvFw9YefeFrEcZaWR
k1bLH8UTD7xM3LRGjNyUVDo6jzj7q56RfvBxP5qbEy2uYBOSwGEV6N/yrDfc3Q8KCesthj+YoBHv
NPbIOUhzLFIuitL71QsbhiiSqCsepz6vl3nivr7dL6F8INUOgsDtT4MBO6VMd+wVLFDlY4ey9QkI
FWfs2/SvQttuL09lkAidIJlU8toP2vU1yRI0E1EYfacFTGJgroef96EQhfSI4exMAXrJxekTpPeR
WIOgN5yPOaccGxj2DA5Ahvl7RBYWaazUnBaOsKl9qPf8ndRp3V19YtxA/nlt4e1HuwltgrvQPcO9
N4hiaayy2Vj1G75rnsuK+qTtVKnC7eCIuFouZQBcXtHUIhFTf/t5ZGqxZCK4y/5iiBuzMzqQAvZW
pVIUHbBatoD4AqeZmhX/Uu3EdwH+GCq838SjLbzSkamm4bzcuoEi2hHDgQDyzzTqtoU/fFfLSV9C
oUkY3KZBhrRTUK8KmGxvrx5K2cCJOMxzFDO8VQqKRtxwmQyf/hEVeo9tEgIrBpHsXbmyHLg+Ck43
f0gI9+eHWO4TogGSrtrS2BUo2dHw9g5ODah4HtrcIwGRc8CtnGpllynllEJAsXgoXoPvy6LXYPP7
qyUoTPdF+rL8YAOzKDX84eLx4//b1cVkcCJn7GZ444yt+/v57FwALcNMfSJbGAxlx57FCK8SAj6j
9M0UeAE3GstgOA74LMfQcaMGtFC+i308+9CinmRuvInajmBUcfxi536Q6SMp2hVfKyZl6iEa1rym
a/nzwIHDv3S/U4Ay2puXcOIWPzI3dky9lTurjfmkAw8pNoCEFQn5nYRQLX4bX1JFkttUm4iLDoU9
4zvcXcPWCbxVQzcQFPfkXNtYVDzGzrCMwpxljoCu8Z41UCTKH/JFWs2QusIVjJuRAKJu6/wOzeJf
OpeID1UfRoR1xRI9bIR3Y9bWI1TTfkt/5/VBAKB0L2C9Fjzpa/HdhpGYQIvroRHYdEvfzzh1oYmW
xyzIPylZUNfVNECJCZoO9o96YKTrQ/zupiHA1ijV8PAghnFx6oMbzwqGoNKxMO8Kw4lUFy2eII3J
C1shFYvS6joxdthkKiVS+K4QRL93ggBc2GnFBzwwRAaT2h2XaWeBZRnmgU0rI4ST+WC1gv19KIiZ
PYaFq+wsg7PI3yWt04flemQMv6FYBWLKgS8WY+FYFqyfUG3JuGINeEaxsbMq1m15lUtZWdZmXjiD
Ve/BspA+UXPZIV15EpMY7aWf/ZNNMwMyPp8CYZKxYa36Ml3epl09dgobg+i0EY2sk0P9PL1rc71i
k2wY3rofEKAX4mPx+DqGkD2dMbOsHUsH7anVdUWMlEmMLXTwf2e52cPUfrGr2PpiDO6Zk9kEWQDe
IhA7Wleidls+D/tK0gN5I0GGCi3AXWDl4QVK9ZfYi07eOa1PFjjc2rQWdtPMHVlRIf174NB/5iWf
ZoCSgpX04v1CCwPpZEuNyJxKipOI36/gPYWqjFogjzV44P3DTpjNUuuSMag5aL1z5CDkCSXJ1I6L
Wr3Ahc2K+HsXXZoaRRc8bzd0NAiIV30nRD/QXxsBCFYqVRzXN+1BMPzPCac7NtJU+7q/VMKKfz9c
n43u5GKi06IpEMFIbmTlIhxLgiTwLL4dquc4DLdihZyKSEI/Z1Pgo2bdGbu6Obpi/aGFdB5wGgHX
reIaxjx1pHgNNPnOpwZ1HGQsLtpt86UFFhbFtzbt5fNizZHhlPz5WKEnlYlkHs4vbgTmh9T9uCJw
seGBaZrwWuVWcELloTncvnWayIfArVEerKgX6SFdPQEh2mQD0Ir+nXR1uhFI/4xlI5/n6dinS65O
Me1tQZab5QQVqJa+wXGkIfS/SsEpD4ZijLem7dsUUDOz3KD8uDTPZtmyLXrfAi+mIi8RlzWpNOPi
gb5VkrFdhxozplC4TBCERUcc9fshnSBKK8Ncy7hNA11LxswcBjSDMvEGCaj9n0GXgPau9a0l9c4Z
1x9jumyeAxwTZb2ipvYXPwoJyJnDWLwjUqjwE3Q2qcS+TVbSlNJChIoxol6DqxY4xvsmKlmtRQme
d4QGUsrWAWDAuFYf+DiqaeZnM0p7MQ7Jxo3mjS6wkV+4l+iHBa6bKsRL1oUlxJGVDxiHz5cNRWiT
k1Pq+RHjfE12be2xYECjpjnzO2SjkcoXstDFdpQC+MH83qGuVxBhM4o3XBFYFzW3g9paARre4pnf
F/0oLGI1T/IKo4aAyKCBSUiAShQxzyotRLdmwbogDxUCslakIBoLd9P+PP8+9KTomYlDFE4q5edl
bRgEUuYiEMGB5xi2EQkmtEAe2fZEIoLBO7glkmX1s9X7+TrFmZ97BE/uvzdMQ9bePP+AZTsX7y/r
bnzyabiHXnUJ0kKBoNFSxZXOylGJzXIeJPvqxs12DcHV1bL7gKDuTKQ9dI9lhHF92TefWymhlJ6s
tCXaP/TaKsA7s8H6m+mV5CpiEMWtf3gru2on4Fx3BAV31bWHUSRzBRo4oVGBEu4NlVMNP0M9sgIo
6KamqOyDCbnXdELhFH+i1mylC+/3Ly50sLYl8yWBOJ4Pjcfr5SjoJQuLcRWAZ11Ycx9LO64OvW/S
/yWUWWIZZlIcfHaacTXAN6YyPea8ESE9s+ekJlx3gPtNYo55wV12Bhe6qA/7kHVVJN8bnWrNAM63
uyIMmR3cE9Gu+obDsMPU4YQxrdvb7sN0PLxY0Fd14akKTrht0tF9yV9P7tBqr0GcAoeUduhKOmZP
737+lbPc7MFYD17ScxCLmHkIKGY6onQCd7ePaa27cCtc6tIMw3qxnnAaE5jFWLATO4eueD+wrPV1
TGuvQBcprlnqNty4OvOf+9K/JcbKPUfg9iXxMP8DjrqEMAr56rnJndefgTF7m/2zknfStpJeH1GL
BqJaSObU7IoLBOyzu22L59NAbNiKasUrG/310qKVywMmeBeb5f9pt0IREVbWIRW6mcB/+B9vXRvK
qxMiSGLxZeDw5qNL0xftYuETQbzorM+UdYZ61WrNsjgZEdjYR8URGue3rGpnMa5Z6c/Q36Dd5RiA
2SJagqPBH/L1abDtFa7gvzJh3gfZHfmX2eICxNz+/kQAwY2gUT40hAW0PDzmOYgA4uiq44+ip912
NfBYyVQtYv7IbdWOmIhxbpKcN1Uzg3NnTwsjOR7psNIVZOUXBX+F6sSWW7S2ngnfuPewzrB+CLwW
+lj1colnDCJP270RdYEapalY3/ty2Xkp5Msom/xYitrXTb770L6yOlbkbhNJ84kP3uVNyN/R5/ER
bH+BoeLGvWdKzNjMcbwisbD0ZZDle7sS0186NJmHHnQFhaS6dYGQ06KfjTf9ewFRk8aR5TtzuaDq
n6fInN2B/m9LIh0oJ0fsRThAId0673/wO9FuA81g0lwH4gZfV2UPhtggU7581lx6A7bC9DmQqyJ5
s0jLhJHf7ZNrvw136k43wNU2yXGofAz9iyCZQYHQqyZmlulR7l1iuohM+Z7W/o/2iPlyMIg601Th
h0+RGl+kSbmKZAW+3KrHJCNXttPFg3/CRRfvVQBVV7E7zvqKQLB0CISrwrnkA0Rl/RvRYmPEHWhg
HlccouWyC9VFmykpdAcSyLOHbEFw4QexCzTCMCKs0a2inW3JjC7vsVxVTggf/ZMKMKHqlPfKBbMV
Fcj1WgvmQUiIgGOT22Di/80PLecXhWh+x1TjAmr9anEWQm40abCs5/etokvZ6Eo/M1zNLSViZqkn
C4SkDnN4OVmWNbM/JwJ1/hMCWCapRikQXE2kGW+w/AG42hGEdmefmhDTY0J5BLKYNW5xtwTi8QZA
LDPbXrjDdb7mCX5194ZBlakmbEqHiCljY26UlSFJFVxxvQMUcolBX2abxZ4xkdLdzXbzN1Bdyuba
ssJo2WF3rU3mOzgsCPIjlHV1+ltx0AZXklm4H64UdSWpiO5Ttx+LjARqaLSpt3tqweCjMxusdBMO
WuRhx+NooRGCtNL+1lb+vOnREK9Zuyudv2Y7FBGJraYttd7IsB2xLM63ELY61dQwDNYWv7aAY1HC
rGDCv13er0x+c+6evalA4fbtnXzmiLOOYHjb6R0VXpNyNDV62vGCqqucXJ2TUNCa/tWHWv9ezWq4
GZm/FNCpAawAFsCqAQkVcVfStM4U+/d2XTxMVCwFdQa5z9rzhVd8InvBBTCKsHYq17pkb9bmE+4L
QHatIkej6psKHIcxYJEKh+pPOYOgQLbzEvLbZOpAzbGyXXG8mqh6KaBavdMplTWwI3Jc4stq4znN
zkulyWuyH/tGzpyDhKrGwOlQP/LEwTBaCc70ztUqrNGTBjYM6gtZ2/yfFJkXuMfXTs1qFLe3PaVg
Mhjxz4Krg3wbFlXAZ8foxvFqjZ3VGLQUIlRoYLsg+jPMM9zh1UfhW17AxF8OHzkG9seuTTHJYHFb
mLLHXk10e3/rA1bd44ZT/y+rKS71r2jX1QKio9Fs+QoARIYBxxib7qinkfkD99L423fk4Fgh+3H1
4BX600Vw0GSWOaSBi3fKOHx/SSbZq9BEkEhTGRxqkbsnE/yW/elq8AcA9KLJhOekm2U9Abyo/UCO
sQpPM3bVgZztUnsccnjvHpf5dLJwmcM45k3foSEGP9Ki89jN1no3EwYIvAktM/1UgOfudKCu1O1e
UwU7T7/8/yxXtR6slCoqJcRpf7RG+NUGbNEXy9jBXl+7AUt3/XcZRnoITGKdap2MVvVFosIHjTDt
Ba+lJb94AOaCXp9lIIUVuKuJitMlktaUv/xnRhJiX9CqGJCw6v/dp9FuQR/xisej0/n1a6RTuXIy
1vp4yuyTyMOE5AnrNQUcMJ4K0QHqJtq/aArYAhQICrtv8Q4w+ZzWPRNJQm+Ww1zAER86RAKjMayH
DzRGpc3u95x4wdhv0dN3kUK48Velmy7RLjAG/S0VX2dUjpxWw4NHPShn0GWV7NshzaRN2pOXpzA1
UMiCDXJESyCZ4926D025Tc4MueLDmN+st1tP3XqEKmWYnvovX6acAqvYr6Ci5SSKxtXJ7liRBkyo
sJPVWUSKpdKiAKcKYc+JG2iQwlkyGIZfEyDx3sBFksMRhQeJvolN8eZQp8yi2SvLwvmyHlcIA1ay
VlPgbdRL7FZXyuPTVJJ+OCUMATvsO5msf+LG5TKUJ8PxtUgWUw8JLXsJ6y+rS+DoOPO3+stLuZgG
8jcHLN3d+/+CRGcStjbhIddJ+JGXzf/zLS4Yo9zQ9AyWj/gR+VVQdNa32oqRER0rXhSOkgGaOFj5
wUDI9HObfJ0PrwN85stSSZu7i3EeTWtqHmncGB47vxDbq0KKcxrY5WE9PWayehA5RzaoBfCd0Nmz
v0u4KJpGdW3CCO2B1e9O294Hnp8o59H0mEe32nn0Qq52yzlIK4hB3q2rLdo5zS79fYjNgwJJmrgl
jc7A49j33xPoLtlceJVx1gkQsmQXAwDq6V5SWlJuIJ4yERtjn7nACUPj0j5Kat0i9xlo/UdEElRH
MwogfjJiGN8ntYiP/XcasZkgwbhyVE6V7t1PY4/K+McKomeKy+XBBLgk/hzfVmTqOg4QbZKz22dC
ZodjdeQDD+Fpr6tJ+HCoo+bpewjqGbz9ab5ad83h2sBPS+Z7nIro7SsF0XAmsWEoVOJvOye3UqvD
0gEm3yfvqQ+uaaU/GwufSzG9l0u2rFQeq0sSuZ/pp5C66WpcQ0WPT+w4MHLvJBH1AWIKYVpvpiWZ
Q+YfdxUI4uN1Gt1ApBCZE9NTQ/ylHRFgl63WqMlni+YOMnLZz3zw40D/U1CaNO4V5r63zuH2KWFu
cqtyMuMX8VYSUpE5t2J17mpMFxRrXDxHsrlAI9FQ+hk4+gUkfJylK8qHBUV6sIczhoy2d3baYZ2k
+7pKXEnyBSa68YTB+6EphcLg/O8NvH77FNxyzPiBD8eDKyfJ638/R6exRepQZ+jx/YZ2twppDz3M
kgDsjp9hm7tE01tfucqV+UkWaXoJWEHacp1SDICVeGdx1BmtBs/MxWkv5m/qbuJc1DIE6pJ8R5oN
z24kHEx7y1+lsjNg7eUijPdSF9/S6rsbU2k8K1juKUcund/OqAYvsGFU/PscRzJwwqm2fUGnqMIH
WKyfVD2aURRZjbBoBc66cj3kIQuVkuLBdz6nFqi+nJQgWuNJzffS7hzZbznHRaiEWTfrFoodmiQE
nR95bmHq2tA2wJnKEiw1NHNsJGf+axK+t9x50AyRKhfSsVd3vDNKTiIMW4OwDDvwftETFRV9qHsh
xWKgam4I6rrb5exp8lOVzzTEBzBDMmuk13iz88iTqQJ9FHmIsT1UwPOHPFFvfZ3gOFgAq/rVc061
8qeR+lTOdNrXTij+W1f83sSqLavoEF4WIQfF7kI9wSBxUHEyOoJcgH/wUnmDrFUv2iS7gkUPzkQp
0p9AtSzzMGspUeYKlhdQ8iHLq6rhF8gHqXS1UYMtzz0eUu0U9wSVPXnHKcbWRWd6TQZb+EOAEunq
AqJwcb1PUoZUMo2E0theZegJNKxsu0FTvqy91PL3Eep1ai62XrJzJA3o69f49qbGJtlxgA0T7Jts
5iNwCJRhCroutQpohA76HRNhWcDp9wYQxk13dTYi+MjjHnnUmN44l/CCveF6ejwttVV7R3MvZyEG
YMM/v+1aqnwoubGGQsKuIktJY+WAWY0PItyR2nKI9wz/zwvKH/1wUa2aYUrGMZ7W+xdDX9xPKbv3
+XlziofT+Yx7Xd7yo5OYGtuSq93vnBuFJyR62fezR9pXw6WJ/1VusgW26MFjhu8Z0xZho1rmOFtc
zGwAVMJUr8Zuh6XJMLJlE1LqHUI/RDVdzvtne9kjx0uEilSe4eq4DIjuOQ34EU/eMVIt27dBxBEL
Z141X3+PPm6dssC2J/KlT5eN4jMqAQ2wDfpbvMC/cxWd6DlntKcK1H2h7JQAHuLrS57Ptb49w856
pKqCH1qcLt7jHtv9htYV2oVF3VlH0D0ncI9VtyBuQByT0X0YiX+kn8IcAqDz20QLi4ryikeFavrB
siRB/wFT0qrPZYxEtq+WiqtVj8Iigdtgyk4jDqZfHcqYkxFvd5pVfroV2Ldn8WJjwqMQlZsMWDAP
2oVHXtmVUpbLhVe5m7YRx3jgzB/1rF0MCfwoQfBM5JTHASUuN4UzzpHMdqOSsoKE8cTDoOi8+ELx
DQLV3MDYjujf4lnjmcrPe1NyM8XQlQu//2Nsu0AOPsnfDTSUjkc3z30OrUAzhmVTb+52/PoG7xrk
j+3wfXRaUzC+PD0dTXcG7xk+wF9/SLd9Ce5Nj7ZxpI6aBJP97Irzz2ikYs9bRhRRgCcMVtV5A1r8
lY6Xtv6pSQDEmDtdDmqq2cDIRAPV4EH+EZC7xvR63aA0C3jZlEOdBpmKxxvG328on1FyjvC6PfSA
TV93Gj8XX2kP55ih12JGsqWPSAWx+M4EYlRvYEb9/s+1jRPkUTNiMSfvCukwHxPLgswMkphQPiiy
aucbTYpVRYdPQF2kUqQHVtqyNBFcLQ15sKzon2v93Mm6F6Suixo2W/8R7kNnIdXYTBpZ8/nXGedx
kvsFkYaMK4sBTKuS5HvzBL3O+2UkETlfpEEVQUYQS3KVZo7+A47OvK5yy+CjbEBpnmVv5TGzcI+o
qec+WGijXFzKz9SFGQ5s0b1NFqGFNzqek0ow5dECSNRo6bONGDxB16cm9j/9Mnj2eFsLPHgmYuoi
+sPKBflzmF8p8jcc2cKa2/p0wqumk/RyOgmXZoi/XPzWLhsPj+P5KZ6v1xACkth4tg0NCcYjDdk8
4jC1Zu+G5/bYShTAU1mjMUdctplLINiFxrUa6Pk+2WQvLu3U928QY0O5Y28YRyB8tjLIMQvrccdO
OcXMaJgkipFkmaTeCZFecQGf2X0bL8iwC+ut6qiDKuykwQSeUWDzmbaCBBQYb3JlmxLJl8uZ3DO5
05Gu114LVEYBQDZS6wJ8lMY6RSxvy36brJjIUVrPxFa3FURLCcablgettBm1zbBNYIBOeXPlZFtT
hsmEV95rofMLskCbJLaxzINCSvQqgSFZiCAwWhIBVuq4RtLyHecRNU3YfmvEgt1zT2qfW/r86hGS
21ScjGgOreeBatIzVTgDOWkUdavSfwGLP80u44pNVWjieiR+/cZ/pcRuUtqvFFw1mvG9591qLMWd
nifZ/T1FnJmWA+4LP8cpP7RZfZvD6gPJXMTqcTyGSiarklqzGTO9IQ7h96S83Bnc8zN8q45oCvMS
UA6XTsjknjayBlfcYxvaHiboh8rfaMcdhg2qAedTchV4pKXd3s0w6GVn+Hcxmnj7j2joq9ECySGN
rboIcQMoWRlOMsZGTRhbvCwavtGeraQbfAfmE5fmoLP0WwGNLdvdZzTfLTgDyfk9QVAFNCK3dNGy
822+T/fTOAowXyfCxGkg5O95A7VX1KEdnt/nEarBfje9WuoXnwEPph3mGHImt1bwL4tNr6xhUZhQ
pIASGhpiPwKH7AT0ynsVdNpnk5ngt34N3UV9+/QBaQNhknu2/MHnJwrFwAfQZQyhuit8n5kAseky
WzpuPg051++njnZpLTJb2Qgv9vMEah2/zEiiSDauYcLao0J4J+SLZ4xM7QpdoSHP4aRKw0ngw2Y7
/PltxEpRTn1b5xKkcrlzk5mlSWZ6HLx7ToNmpuLVagEzTLQm/kV5JKeZaFFecRmq6IeMpfAUkSjT
jb7FpE+JHPq4ejhdrbI7O8AAExo2xz/nUi24NVx1RQkX4Fsy1UwWQItPBgauBru7c2+pjDPXsKt0
DWbSD/62Je0uqoL65HnxPhmt9C81yNIfrV8f0yvp89oLozhDqQaeiYlB6qdRRjJAiiDm3Snf+isa
Rmi90pmej9EvShm7ydfSonsf6hq2G33hMlWzx6hJsQoPFKNLDN17sbFb8rjKND+3LfLtOs1wnKQN
4EPX8Y7sEscbZS535OZ0BF+YAKkaX7wbe33JCKPNl28fhfhsog5i0k8wPHEufm5kzw9R99W+fWfx
oJpMK9a0FCJFTWs6RHKWQbNpKgOwtLx+I0ORZI2ZV2TgxB4t8EkAgTVAo/tRnl11M8muItarMqzw
1mG8eyIB/3hvylkuBQO09Pbt8irN+BQZZAdRamqX74vyVVC4/b87zDazBikwNfs0lycCWVu8n/pf
fJRWgEvfWhnrI673FI9/e95GzDiEEbJD2I89VQBL27zeov9jx7Fec/xnmeELRSAhakVXr/c5jbTc
40TUQPSduuNaqkpUVWB9yRGHUzZpqGT6fZm1GQMhhfhnbzuAF/nvsRSI1VrN/tSj30IK57d/Gxnb
t9SXjMoxihjXxmBn0v3pWQlwEqg6q9Y8rW4LyqLTyrUxjMkzbIsKW3ZVA0NkHEyQ++OICGJUPJeg
2mo3zPsseEHGPsFySP256Ly7RcCiGtBUdKKm3cdAE41tQuruGH+ms7UdGew10sacBHyOkbqHBRtD
hcTs/rdVoinxl3jEk8u5oVBdGrzUbyb5xgmzhl45I4FZwtX1qWEoZxsn+/ekXhAjC61x0gNHzF+q
65KvIXsAFbdmENQw3PrJw3o13zrkLJDdFva3x4oJg/S7b8X/ZwuwO6YXnllifAJBxPtid0TNhUhQ
VmNaFeN/swmtNcFjMxCZ+6+Ykw0086+dxcQ4f8zvzgxQ6kDz9NiTJpiqg/yU5m22QxpCb1KY6EX/
mF9YYBs/lMnVCv2Yt/6hziMgjcMxRnYvmkwXm5yWIDSxseW3eU5nIrIjV5L/1p/pr8yH8QvzK41b
VgmK4UWURnMwbMwQr9+5tVv2lSUSKZothiZ/uaEDIbbPAfG7ZWIDkRcstvn7qtYpoCSrck/mXdLL
eTpE3Lp8DZQ82aRVElx7bCPM2ruw1sgFGEehot2ifObq2H/QHbjaMc8ix6e6dDRIw2txQKMJi0CY
KRK7aaaDncNoINDug7jR5W6aFQwE17TImr0r+/tNylVfQ3vScFMoEmLkRjtdl4Sz0VA0lw2ufJ9i
pwcEusphfm489QWfOF0Biv+t3LyoNM82rCQMlTYZmxDh6cUbsMb7VVb4AOoBKYi9kur1Ts4fz7FF
maNjotwvTX4ngYlty1InfMAocvXy7fZDmOPwenn0bHGOpVqclLYdksRt6CZVVDGjwFWuk5DV1wSP
avB22OqP62ndGyYS8FcwIkk4dvfcGMVea3pokPRR6ZQVuTAB1HDp6i9+n+O1Lt4ZadAMmmsdPhib
AxrhDKqZ4uyc7Xzl+Gsw9xjneFuyWBpuAER1sMI3+E6n8Fpj6gxkmvotyx+mU4ERnZW1nXu7duuw
jEVnCPDSNrWFMd7TyYNWms8U4lNKyA6a35Rem8an3+nkASYVaaZxHbaVS3QHU6hgKk56kOoUqsf7
G4HAYeRCHhdPUx5iKLO+1AJ+fVALowrLUBHY7FFhITqFZMNA9CKVhYEDMZqE7rr3lN5gmzpIbgrZ
J1HGPl39KBY77LhIdU9k5lWpyit4UWAb/o4M1uxeL9Rv4ZwvPvJJ2mRNQaObJSCi9MkQvVhoqL9T
Wk5GlRuZHfizQ/6sahZDPywqzXpSsPvlOWU2H3dURt0zfp7+nVUbhsucQLpyXfbrTgvZq97gI+Iu
od69P5bmG0GZ9B+dLLgLY6KvS94CrNLwvaM1QmM7KAdjYrY9Ul3s1yskVQxSl/2bIxds1FM3C5u/
bA5JiJos3+AWcbre1z5yzacUXRpS4R/vKl7QcpNSdnKEdaYH1qUWXFgQh89KbmdUBXR/HkHtCLgQ
EIml0QPHBJJZ/JwjIZ0mOB1FRbWy5AQpfhqmL4Gwn+OuU/0JpW+dlHQHgoUmPjwb7XuDs+0+4mjK
CmnVRYdBb6F4BxRA2ffyCnNpWiYaApNx6nLH3PxzHiwfFxGR4royymU9AOqq4qBRWYZCmdOg6+p1
+6DOUjC32J5LYEvt+ajnajNh+qQGdRs8uJCCBmc1YDpAFVHWofdsbad9zJwP8bxkWsjN+7JLNSih
oIK11obnFgkaV0KJERPTjSxa/0A66p3bbWQhsf/mXMEUWOjv5CN++kN0xcNre4JIBhmtXS44EK3R
C2b+28hFCc0q2wX10sfllKpjCOU3JlGixcSiEqn8IORCfc7+U7rThCPROYxxbpb+Xu/rfksCC/1m
2etc7pghiTEkFAEOXRNwbLoquIBlSV5zxfBo/e6s7G31UPDffJTuiAxpk2+oTmsqdkXIlaM6fq8n
/8BpXsMMoJuM5pFMqxARKVtYSfnPkBfixXy9/+fjIszmCXiPr1Lj38PZr4iZzIG5dDu0kQUsLnFb
yh9vjeDzgj7ZT1RfP8olD1Gmcac1YYg8S7L866sCtjQufYsq1r8IsGk5InWKMUdDxA9AiJP9/i1C
GIvS2C2hKeC1h9LktVP3JfS4WGR4bFqWR+DmhWzsIzDo3eknQ0Py12fGVQIx6KN/8U2yCaq6D2ij
T5yOdPQ7XJesRADJ+VxzMV4aYEpZ60a7EAzoO7Wgm/z2+kFZ67vfMYUjFD2aZMg41e/XTr3D3Ym+
aNpAJlyisrFiZEYKXHLWHA1h7bCp7HQrJvc+0rVp5Gvn/Tsuz1C1Ki8xJMpbG2IX8yy8dCSQxKiY
HiYsHjgapZQPpo+dsubH5IAib5Rb3ZVJdjqqWLwfGKi6n/YQVOEjZVaetGq9zfMZdzECT/cYYWcz
zs6UjzFkrgQ/UXjvywt44m3ZNP4LKzlZGcp2tAz6DUhXtGPCX5wUcBeEx7H8sXod+5QL6m0DPwEb
KmOCd/4J54/SdmqklN9iDlRFV9cY6C/lhE2h+9jE04JKPMIs3Uj0VtTl9pC0RlaaGzaGfy7PUS5n
t3uTYnXyigTL5H+8FUXQfwyXYptFgvpdxDLtnlnsaa8JTZCD1RoLpI7qV9dbsIS/ccl31OeoYHW/
p1/NFyCXNlhfhI4Q2mgR0TbkeJySP/Z2uIZ4QxYt3rCayDDIWd5ySWlQ0OwEydAPsdkTQsIbWziN
9CftXYp6rj4hvAAQ41YkPepN4KBLdH8F1OJWKd67qzJjD32jd6kkKkFZR8KArlmhtYH7xuuM2wmG
FxrKoFszn0GPM0RS/UvHn0EXDQ7ZVlV/zznJbaj/ZLTd0UN14StZ7ZkfGAiduHYNFEcgBP2g26oO
HcCSvl1hxijdOMyfPGssBZuYRUN5H6bK+07B6/zvnqFbfLI+pP4HYrEPKCxhjMVF+a3Cn8Ntfw2A
Mka2lC2RzsKOlX80uj1KRWoVPG9WtTQ51h543i3nECfm7mdySQeQ2ebuZ9J96VrQj9X0aDjpqa55
iSrx1h6HD9zf6pV40EPYZol2kg4f8770BfKLhwBmzVb2D2sLYQN50UId6EbFJ90QYqJWVbHDkR/X
ax/oV8r54P/VGuek2K0wdb9EW/bqcP87/dojcwXY4ddPLrh7Pg53oNt7J3InvBFsy6vONQPAzHfr
ekrQVQ2+7oQ7Q6DNy4NHOhrhHNGc7q6uHMcXKcmJIemIb0XxOrPM6IhxgwKEWehc4A9oNIdmDFCk
16ENfK/GVXY4dWPPkOSfqqC5HhEK0L4if0FkrmQFu74AcnbdvxrKIAbTz3LeUk/wTmqWWqheMsy4
N3yoWCekpoMfTseTgyNnsjGFTw1flin9cOqXI4Xu5z/2+sIrm13RBQzbE1ywr15qxSajb9bf4aLI
xGPvnPbsph+EkAfhL9egLAh9anW1Wq8bjmHC4PHNWMsuXNNzRtDAoKwR/x5w/cc0R/DhbSpzypzC
vQqqbWzLqOXw2nkxlLWNFRYJvrT8XWmng5vhZd4I70cly4b/0xJ4pvvHJLe0aR7uVJbno81PL4Zm
xcYBMFT87cZWHAeEYPajnT+c20OSFEugqKPFHkTShAhcIMXyBBeqrCVUw5r2m9EFvvJt9XTTnOda
2C5a2Qycna1PyRIZbJ7ohbWkAGV3pW3ppKVsLGylVRQG/+21MCh35Ts//jj9G2r9RisOjB8f0AC7
EqNedfrkcca2clfs4rObr0FAC+DxLsvblSQBESmPMo4oRbc3uH8osJ0F3jeCVUm/cjhJ2hiytgP7
dVRZ5Odbw3e9G1TCKfI7HSivM07KaJELJltUGfC931U21s7oiR+POiAaXT+WYV0iilbdkbuHS8Km
niDvxfk39EurJIsIKY8AAf9AwB2HvIwnj++uso7kOzGuRckmJYr89ThPhLrhtZQHZ9s4RhSnwlzm
ZuPGwb5QGa4ke53290MLh0EG6s7yKJ9PpcEqVFf9aIEFhfH/Z2xNqAr7yoclgIKiEjwiSzfmw0Wx
jV4ofXD/Igs2SagVkALb4KgYpCGopK3dwyTqU+cS5kntwjfZVI/ikIA8YTNzj+5EPPy+wJmxyyBj
kbKTQstD+fWoBaKa5wUfh3DfIDlr9XlyM5209IhqlxLG3BrDkRhxEdAyj0Qq8vck6oFD1D0Xby0F
ptlSIB6Lk8IbUIEmK54SC3hYhBaMoIXB1tr0jZRSneHT6vmoN2kX7xEtmXKRTorik6G7bjRfNoUZ
GPnVhZeUSomExf3HXzUqc0su5Sm3v8F5H4IRQB+Sk10/xCgSYy0lU/PQM3xpZ6//c+qutVLKwQKt
pQopppUZBLfdDFIS4vOrbMoDJmxSoS/4O/EKi11d9Wh7/H/enXLqjdUZu1ubf2R78aFXxX6nOWn6
wleeb+OMXR5tJLUfBv5ClqmBCNJTywgtCEmpd3jMKavZ24hbgmEEKMR+F+rTHDgb1vUkz4wMDzsO
E+E6gg3KhbNtG316Ej+J/kVkvDH+lQMztCDlxeSCk39Hkfw9WIja88sYL8mhGkIz72r/2a1vOkwW
xt51PjJFY7BvwDuNaMFUpkdeehsoxb8d2avndnkNzF4ZhESD656L/+1+JCR0aqetAB1/7Q/SsaGK
tRFzQ080joKkU2hKkMkB7+C4eDBzwEbipyc54tw4YP8R5Ht2vio7M2onBy1bqYrpHEAoqE5Y1VTi
vlcCFN67o18fZDGMmYzKbApKxsCh9YJ0Gsvn+ALl9IGqPNqAg1mH/V2G2QKLayvqsxRwKTh8L4/X
u5/BM1myVmJQcRlUmguEBoKjiAXS/ZJm0U7t3xqj3szMe3Jcxtv7On5Sg+gVnI21QtomHCWqcG/s
zDegZhMgmuILL0KZ/HB9raxPHqQWU0BwVu4ePP07SEeG80ny5MxN1jT2hvgggIzYHD45y/I9VXwF
vNagY5EVwyKQfQyid4cfhlzBV26cYcgQ8yp629VJG3M4hG5tpoQ/+gdxkfz6d4Turt32uI+ESjSm
aXVRz7VjutdE5+JLrxNJsQr0u4yjm9actBQcnI2j6tqkphY+eRDgWXDKCVZHtkw5sTKByzaY/BRd
xKLY9QmHPHutTF4cHhcXdb721b4tkZHQqZFt9PfM3o2+SttOJCMnvwxYn9OPBrB8tnEE/Fuqqk57
e5O9GKD8TEacruhCawf0EAVws410Oh5BZH/eM3lIsuBYWBSo56IMSSJXksE+gmKeksU9WBIm9gUL
wOMEccR2aGlhYu819Ehpy7h2YHk8v2eYrFrxgh6eaI7EkoI/0vQmgG4rYK6tlDfI5is97Dc2ag+Q
OdP3x3r9bu8kwyAlegEmgwLYrTuhgZ15gGCDZKlpPt9obU+FWfh1BBYhgklx2b11yHeLnEr3j6tp
ApRseFOlmVdHpb3+8SdZ6Kl5JdTN/X76AYr6hy0hm/ds91qxu/vOavosMvMssy3i/8/SzzbMp4B3
L3pO4djrZljcmemu4tvZuVk4aXU2oP5ngeUOJ41WVu+cbPbvB9u1z5A6w+8WycCEI7yEHkCMqjdZ
dhh9HZlP4O5BXeS7eNdfLshGavB9RLxjEhJdRMRpgyJjdflIZ2R1AD31fFtNEtGj01HZFvqXpoVy
xHtKSRmrFl91JgqpS3j2kOy3Cs0iYalWwEejzgf/2MonFbYKN/6KzesE6v1AIPorOlxJa9RsGLga
WcCUzaj73cC9i08S2zYbcWodNnzGoohGLDS1yTSHju6DmqH/+UEKEPb001BxhJ28gyEMbtw8HVvR
dsg6L+d7xLEHFaoiAf41fhLPEy00sFHLdzecMMykGMKPeEYj/0PyWijLu3/UhrV8hwOPoYWqWDTa
Hcnp2oWN6vpatzudVtjjJUBMYKs0jxzOxaTiEZtiLstq6oxyVI3uZ5cRPZYwEjXexAYdpmgkoTxf
UHizV0FBAP89E/i+lraHlZOBJHNzBBxqmJKve4t06/bmthMakwqaFJb8mZ9K7LPQnk83HUi87FHY
rG4sEl+j7bIxRbt9mF0hdL9ECvgGtFoMpa3cjE8qfZBjqNEEeMb39m63OqiXJ4wk2MeiLeBYMAU9
p5QN7nx1l0XP+P4BegaKNELkAACyxFYKqcBcDHoi2V8dTOWswIiUgF9vY1IQGfPkuxLGAoaUQaDz
xUqppt7ll/AxzZnT25/poCvxL3JCDTJ1BnfjeTq5p0CuoOhFD5W5H52uRSHczAozrvk6sc640E8u
b9HUnN6qOnXY4DrPT6+XMFAZs7jvuNq/ArIR+OpyUZmiRelj3n962pukTy4nR2qBo1HEMVCoVV9P
gvxo1gEjdApQheG1kqsTSBo6tWvvLdepW4z2efv6vhVVs9RmtkoREZLw8ZC/sVA+uf1arx3k4V6t
9dG1c2AheXzJs8/SkYnlzdwEqJP6S3nHz068qVPk8N+ciiV8U7HDrvnKQZt97mrevfZQ9HcYiPMA
tG8uWAH1Wu1QoR5dezYpN2MGw/VCx8L6boWLVZEfFCjYobYIhghBKe+WNZ5IMFKZNj8gUeX9gZwc
oNeUKHRsgCyso0Q6VRZP5yAcaebjyzLXkBf89XWXR9zP17PbGSEO0jy8L2TCRNVwDTL2+wTC1dM6
cNkryKbTO4F8CG1vQyOlMEc5fkMYGncZS6qmYdbcbeTCxzNQYxRzFiv4lboZ0sDWg0ua15aZ2JY7
QrV8GQ3bZqeZnuJI4myqM+rfrGnpZL4pxxIyPtGqBAfDiFhHGTEyG7fJlLeI7Bddj31gTJYaliWx
yZQ/uiVtksTnt5fNCjwLH1kF0y/AQq2/UI/keu+HoSkJg7fC9xKCeSWvHc841IkynWRpBZqH5tj7
aE+TeI8P07jneZwtSuuNoR9R4W0h462GESXJHjxHTKfTckobZOWesxTaxVoJTtpr4iJZu09Kr2ro
5icFd8s3/NMLz0sSKUxvq1NNyU2bkLBLSyTjy6sLP4JOjdM7L4LmXGwrWN9Q3gPHkEQSm0r073Sk
M5yC4DetZE4HW7+tEoMjyRYnBRwHQ5i2+0FAFN6Axeo5GXPOA6oeePppld0AYccL5be55NAH4kpH
aCtjUZrXtoiNhA1trn26kmeZQFqAXfk9AZBuYeIZRQoWcM3uNZO1iDk4YWLqrZoT436bzdsRWxHk
uQ6DqfQ7/SMfE/plpre7+fjRYSboORdFh5qdw0fOCwzNH0GbRKGrYYW/QjNS6FXEko1a4/0VIdBk
ZLnPOC/mpjc0FwO9b3UHaoao9dJop++VwnnmMX6POJuIGpkOkcDoHo3bshLaUOYeitkHxwjqzYdv
qypiJg5X9aFd7DDqn/+SlVJUoRZxOG/NN56uiIul5IBhhERxlx/f0fsm4g65ORvTGIEj2C9hkNzS
GvMPcHPhZzHzrtKjPgLGQUB2INwnsY/8ZY4Y0u9z0hyEXLCj10GtSoOZx09fbreePhI4tMWqk5DM
NCD3PbbsGljkxHGxnlXsXvXMFcjn69+7BPdymLHAH65pthN+Mt548PHbsOSMQ90x4n8sWevo4TBr
1Tc0B0QVRcqkvSjt+liyFGiLy2o7mGoS7LoXCc6trjy4ec2Siammik/pH1Hx5OLJkNqDSUnuwq4f
mNWDgboGBMqfXuv/8wacljxa2MQFeYuoc+2n4arHNENPgePVImHUHt4KJopFJmJUhg9d/EntjusV
N0diPqKPSBchnCaGbGKeyDEo9ECP/HRi0+VKDK+9rZ/hiEGD+ZNtSuq5EQWJw0XP9KQu7wWWaW0g
SWMYppALUwyu8OGgSjFg0Uji7p527Ixwbkk7xLTDx6igg4IUmvuYTXfiRLJLIjgmbtCZww2+JJ89
gzykKXC+Ua0YuX3141W77hwpuzII+I0VSxrHVm8oNa8Ir/WmemrLVBuzYJUv2Pth7zDpOQHdCuqA
lYjvHIUFvj+QU6AAT4z1DwFnuWDODqfj9I95TGNKX3ai0JrUIfmAtYSGo7LupQf3CROC1tmWB3qs
A1ZV2dDhQY9A5juvJ3XLUYS0/hKtasc/8GB2JUfTUBf8SsuYvzDCwQFzvu/rbd1nKd8h238ArpZz
Re9XVNRVDXKCvkQhWH8RWtoiAb72kar4t2gPWUYLJ5GdzRqt7JsQCYl4wGzbwChQOBLmsKGho6SI
3+lwFHPVKJFFEbNO1TbN3P4nBS5Jh7yl9zjTf+BB0THzZx6K7BxdjHriaob5SjB8kHzwmeWbMFXG
aPQsBI+vW4YNwGIeNZhDjTc2pZzGE7Tmrgf2kejdb4UD+k3cDgruA6otVK4WRrmSK6Vrsr1HZ83x
LPpQMNaHsiZSpMQ15or9wXz656tmZUYGPczz577hb8RIdqle2sK6FcAGu9CtP4uR6IKlCnQeQQLL
wf7UOSlxlzXUa/g6ScoPv9+5v/vFoPA37uvLiHRp9Ymd2sk9G+LQ1e4nodtkk3qYlOg6fDEdumCp
IbacowyQVilqV6iB+6JPmB7EtruaT2SpN+7KXSoV2xHY8W2D2luiC3QWD6FApa3c8PxJxXufmyI2
EbCW6ZvOt8bSyO3Xe7/j9+/3p1SzrZe/p7AofN/PTkVM/lqA/6Q9a8vV/3Nh2URZPqv1Q/iahXzv
PeC95YmNNxUbvBwdUlqdBq55/mv1eA6MlI4x0MYruBCnFSM5ZwlTyIN6GTl7NzGpyYxnvtINiGgw
pUY1/lxz2mQ41C19XC/Udpa6FPBff9OcmrmFE5JuSQmlnSo2wFq16s2RVIQafr7PYKNX+Hwo9QMp
u+qvk5rFT3Q9owuCF0Fp21gZD6k85nbSGGLKOv+S1OVRa34WEFKhS1ZnzNFpI/LNoxX1a9/ZC9Z4
/fQYEzB9GiQpkPL5q99j+PIRbijdAZVU8sNLIqBO77KHbwOu4FZs5LoVToVAmRgrU1X2hnb8vjYY
82wG92tLZEabfcYK2WKJIXwTZYhH5TjTF2u1NkPKshIQyHOqIkOwoJ9tON9jKd1NTRcgLPKKeOuP
zBzKZsvCwSkK7cbTcnEA7HpV1g118UiQATpZYnSTHouqQTv80wNoCxCB3Vwls5T4u90g5QB2uUnY
1qzgDTQZ+MxvDWGFPw3Q7SNSfNKHocgzTCnUuiEUMTP8PdqhYk7kA11ml2hyVlm7/Ivlx0fNsRoQ
6Mc9sZJ3AK3erWdHE19Zc4zujIDD20yCXjOn8yPdOWcXlPVZqiMLjlb66mQYIAiN/HpOm5mrpXgs
3PSj3BdL3PncxcEkf0BnsqrT8r+VAZzKmzjFDO+lJDVO9DrhppIKP52MHzeQ+FH4+G+NTgVecLIh
NxnY/Id0GlvPq54V20Pf2YEKp60bcKefELJuf+LNabJEbKxBULXkkrswBCj7S+7x4aL5Um/iyeOk
0s9LQHqbs0/WRibNGUEK/5D69oURHIsQGWzOEvLIrz8Dkp9v1A/2/bMewnMX72w68XSGL6GX9HZy
wd0B4Dj2apQkI17QUKdvK/o2Oh15bs4/07kV5Fd0fIFo+s7ca70aYXGSlVsRDhSN6Pqnt0mM+Pec
ouatBj8VAI9ewFYS1FCeHqHAFIsjDGyR0QxLj0UYyahIcza9AUyvoNkP27D3sepWANkcI4SOFbRf
0Jm459+UT48tN4RvXDNQFzV0Ykz/hu254V5Cy56PJz/zgEYibxse5mjrKbxDW8ea1FqEm2N21Aww
Hl7cKb+2olFE/aQDl4H+5LKBjwYX1ejuzYRlPuG/vg8hMCQxCnJfglPPHyWepmT3uX2yfHJ/pxDP
tg+GM/vvuoAlJXXvuu2O1g3qxyKpiIcyPpVfnQg/gFyyGQ771OQgJbcN9D7D4llRfhCspLmbH21z
fryyHkH04zH+2SSBtCe5pUqAb/Vh3Y1hOJyKJciHcL3Y7dXp10Zy4CGr7sB5alll0ASDaOeoi+IF
oU8hRsGk5bRJwj2qGGJUdE5wLXwix5YiyMIwr+blaDdnaf5ci3+Cc+YfRToK6Nf/N3OyN1SMwsKW
vV8dgASQQ8NXWvxpmLL7c8aI3dsB1ztREg1f1Ok6jCnc20YYYivyB3RJzVAu1g5c9p3iCwWdufoO
5GQG0XyKtXsJxtEqpkyCmUCudGlgZWTAZvKui8Q1OScL62BbfhRwq1lJlgWL1P1Z3yJxpUActjF/
7ge3cOGiDGid0e52Bo8PsAiHiBob+2wJ+6hFokKN/l/vHd56MoN1t7wv1gx3xDo/ZLtWPVvuC3xO
Pxe0C2yndPOKxlljAoulXG2MhGiApGHiGof5pwGzFL9K57fJ76jCX8kDbEiB3V2Hgi3WrG2gk11j
eSlLN31kh433r1qSMmmrI3yQu0t1CfwM373Z7rNnCePx/tt4B/LJgYrZZVbU1B+yyuDrCshJVmrY
KUB/KTOEa3v9ut4R3yhLGOS0d97/pw3oe7WppahbAk5t3JW41Vmvafpo52L0u321L1YWCPdmBRKf
U2R4XKyAPK12nVAw9TmwW/fdlNfXUB2Y7/3roeg+nBBx/o1y7W3mLyZEvdWtIaaJyJS0amFO7giN
IFNQUKEoY3xUWWNGzouFFWby6PKeOJzO2fnDSoSUFWVZEa/EyNLhQhyFdfqPlV9d+X2PR67nu0+Y
619IjBAkrNFqdLdXo1NhNVaUiFZkk3pWeNzj69caydwmzFlD+0x/klk9UkLNQn6ZYTPA/UI/d01i
G2BrWYEaJ4OOIzmCc1u1R1WKsV5OCxSpfRmuQddi5xVV0OocDHNgCGlhnkTLfwrPPhYOIzch4gfZ
T+KB6SlVY12SeaaNGGHrZhjyohYn5QvrwXUouagGxV5TOB2MPSSeIQ5mxI0LE1BY8ROaZuBEmIB7
9RZ8BmxBJJUoAs2U98FN1kHu4nwBZ7K9qKAwPaXPvFf2Bk2r12d51NrXnmaFdE6AZ5diwpYzapR4
qqlvsc8T2ReDXqj1gZVJqTJi11clNg7YmzlISuQv8es521htGTIsUD2oE+ckyJO/uwmyKmcK6SLn
8PGWzAkGtkFLB1Uf02GMXN0gUCdW2rERBjlpHiznQrQPRVlbSUGgwnuAlhn8rcLKeU1snwwhfFW0
bsz698Kpnv6X0WdrgcFKEMh0mqQ/W9pQgvWScttr0Xat9Yh2BKYyFC4OBn+igu6q1OxxfaxvpZP8
6G0lmO1L3Y0ozUbdglRi8Kfh4fyxJEo8xzPoH5/SIocwsTmTD2icfzbLYxLQAtZU37EXG7v5xOXS
ZFDdvn6wOqxe5em2CF2mboSabuUEsAdhXQQuOBbJstVFsxWXLsRe7U5W9uU1qgEyrj2iRoQ+OITw
nAdIHUwj4U7Px/OJfuB/jBlfHbaTFEAZ3Q6HTIeimAHZzEyiv7v4eRu36m4KMpYMcuwGYgm47s9j
AY0s5zQFO3g8nogH7pcxrZJ7P26lAA736KkgWgVu456tgS41t6QTt3TH7Khj3fdqGRp5jRGYFSL8
6CNuZRn4RYfbWmBsELEzOEVFy6hGx4iTkgY4dP66NpY1j3X3x2hf50xl36Xoxn7/zquTFjNIN8a5
Hb+0Lt+NXC0VeG3/eq8u6kxyrvkSTxpUyZJ3Y2QSDQ8zN6Dc4f/Vnu2VYa/SwexcDBhB0s6md6c8
4IW/nDnOMgKomO3dwgFkV2dqgqv1jZJRaKWiTg6h4R0Rp+Uot90o/L+n76pEoIWEivsHZr8IZppo
4jVYZ2s7+Y0bHBD/vqDCGvomeYaCkY/I9V30PRLG081KqQso3VPr7r0kv6ukX48BGEtuajRkmfb/
D5fw6hGqaldtJ68v98/0gqFcWIesoQ/IU2/XhhQSzRIfO/UVRq8hnsn6Nl92tv5Jq5zxNVyjz2kg
B0eTqJgR7GtHh1g8gS2JyADgHRhc0nhDJwYVuYp8Gi2K8LJL/heEXjWHSpO1Shv//vZSk38VsjDi
XnF4l0n4wqQ857Bei6LFp0sLsZ4Lw/S2EkcZ8La7v5hRF8sv4p5SJIfixY+rB6FwpM+ggo3d/Tmi
I/1ltanxtf2XdtKAbWB4GLepd4OXJO2+xeGqMwr3wRjw8PGuXrb1rpZdYtVzeqfvJ/skyLX5/8pD
Xy5TtYCS4svhmPal3b5zxgvzNSeNPcYLRw3S7UuqcMiVD/oj03kSrnl+zOHGchLBplP6Wo61mWOt
GKPL/MrlJD5z+AOldeoNnNrxCOxtxGftANy5AjbR/5tcvlnNspT7ZzAw3A1sgFZHo88Y3yjMjnxW
SfmaR0LzU7wBzcUlPN498Vb+IJidMhtJqEI8OtGA/LZIxWEwEgl9gHGdahJKql/c1VxT8OTjautX
uc61qOBYp7ijkaNraDYLc3ROE4Lk4zWg3xEsk4bXOXymmYwufDPHqt3EuxcJ92VmKIQXQaOEKM6w
ispSOgyy5KSpFieE3A86GCjeiXTfxnLVb9T28TG7X31Sb+d8F7y4pnlLFHUWSX04BPRfiOXOi9EA
4TIwSH0DlNAs2bS+h+hK2sLq/SjOO5eJjG4vQDHwOMJJUCa6QnmYjNmqdoeyMw3v5s+HFHj1ZfuJ
JCn5lY/1a1xUARI4EgR7UvrxwgxByDRUodKW0WttmVnbabDtlsJ87ctwbcVlGm2evlnBHAJyyBIQ
R6yiYTRVTI3XA24qwTZwl35fY3QOUvI4G97s+n3b2wmVMgtiIRhW1TsphI+vixeTSRKgaj8YEacP
yMcK+PlxrsEKCSNfmiCe2gurcKlagn78prt/wt46XxJJK1WkbNn9rw1e25ba96oDS8gXKuBMb2HD
rnpUd8XAKdlc1OiuehjTi/97v29v11b8rVJwII4uT/RVEebsNTTUrpsolEB4KeFeKSuY5xyroeg4
WuQ7IN7qLrnCsO1taXYS8lkc3VJzP0jptHDLZil5qzyI4bSnaCMf5ynMB158+V2KrrhEfnAmQH64
o/4wUfrcYnpV3qXZW9Hq+uE9hZJafWqbAMapL+44Gbf1Iu8t86nhZwAr7Uqn0HYH3iYLrrZI0pi5
yj3chS7GtzKI9QFcLrRoA95XV57qHn6Z9kb1HFVE5vRqarxIHwTmisQSDzp+4CALut9IyV2r1RCp
CLawHJRgLz+E9x1szJ/hRmg4O5DPlhOyQFhavgAxWh1PPl5vZa54Cq1+UgJM6srfFN1Mo2m18CfP
iCA35/I2uMu4XhFWbwjf3X0p1AUaqnF+DcNWcJwOOJkoMqzYgQMVcuu58lkU6L42W1rykKORPwFm
v9ZTLh1em39LjhgrxTEl5hecfbMiCqzuRvs3i7T7T/RKT31/FpProl5E7HKEmXfOmJkfJfiRw4Eh
XgTCmnbcbsCfWNddmu3miS2GKjGgH7RTHscOapku8monYsdPryS2yqf2SDrI+LiJ49Uz/vx0cZog
9yQsh9pE4o4b2ijWGEhL9rTLssCVDNQslbxJ9BlTNtvakY2nK0tpGb5OU4Q3DPo5A2QmfL4X0/iO
U3qVBqf5VBasjbfrDkp8mp0fxaOC+hLjwp870LKfIE6z+7qli5jyrADggjEYHi3B/4Y5H+FqOlD2
zWxeZxIk5XYa3g7ktaMEW/HMpLXcdyhlLoqu+bqz6dM5zM/CYV4J12GuG8JvrvvZ9X7T0sJDyFYf
Fxlxt/uzFfzS7AIdlSTWBBqWXAzIPPFCu4he1uOqlzsVc0YxyOxPprjfbV5JIcuoVSs/7LDIhqc/
YPmEhTfUTgrnIhp7NW1pFMfffsoaDbwS8tpZF+s9XNhOv6HJsSLBVrkqskKgFdvCqbLcIV+JEpx8
q8VGfx8uFTzu6/40PCtgPAjOEk3nIuTUJBhDpgCyelWuhufpvMwrxXH34SW7UiQuwzKe69THrb7B
KvpwYKhpK0e/lUuMZxlWzFYOyuA/V3hahKcGCuwxWAsl8qVs/pXbnCihW+wr+NvmXAbdeEO2AE0y
ZH89cuolKLxcZC7nt90XXW+LtOsi/MNqhxZyuf+lp26avz7n9r1DoruSHPyXzK7BjhFppPnuXNt1
9yfCxuJg/6fVaWqQpuIqEsfP8VAbvly44dRf23X9Wezr+MIKMzdRcINt72WRR8vYJ8OvbcUEU6zu
Gysbwrg/DbrcewM5kl142/PoXFSF8WoK0Y2buKlWQyxkKwE0qgVPKkH826e0vwfpQxMLdAHE7H0T
xQBfm4TouooEp/MAU/rMJFsd6ObOns8UbS3zfpJgvGVzJDCyGoaJg2tQiRpmHaMJMPcObewvUjU4
2PSnilKv6rW6F+XObi3wiglDhOBOyj4cSWfWUDTOq8+BQ1av5qycjuwF1XRswGBgvthuiHQyRX0a
U4on7GXvoU+1hPRE9PaBDJvI8yrdFUc7xPPpNttKoUrpSA9Y96GBM4f0fQgDEDZh6S47N5EghyN0
Vcj/ld96ZQpr/INSAM94mH8J5/2wtFNaif9Gki0AvoU22csovjW8xARh/J05dV6xVtBTThPYSkwF
ZLCZNa3fYs0MEwTtife7OuW8V+aeJ3sDAWJ4dzhabYg10xsAt1CnB0Mw1Bk8Qi/7NdYSK8njcIdn
SeYhbUXTUqweElNWi09bzizofNVEwShwCWzqBgGkTbBzME7kFk8Mr9tVSyIGcISxMznnz9qRC33k
WRw5Z3QXCZyO4KHcpcaQD3tJgRlMdtXLd5QK7BCPJ546YZ9LpB3rfapFake5nxM71aSMYsrDd9ym
ZqpeezxjQK+fLBWttZPrC7157d54bEtJx4RWeYYeQyzBIC0VwMAzbnTLGB2wt4LCYaxlRI7+2AnV
UUQxJNTV+0iTwn5kykA3pdBXg0NaYBv4cQkOzQjqqIEpGpwa/0IB+X32rvUBCkZnDb4S+wNeh+qR
scYvhmTCW08KtuGXXTEBObev0vokU7Ab30XMfvvO0FyMabzGOAGsVZRtMqFqwjJyK6Ovf0vFcseO
b+OgFEHQHnV2VPQs4A4rAMUvzvneza4LJ2m4hrutAe5hJ+h2OGPV7PFaCmAlILNPKeHju2/+eU+t
nLm1yC0CGXgySNsrj8K/AsL4/f2o0vXgFMePsy/kiBa2QOzUTYp6V/4fFSi5IzUZmKAmDnVzLOKn
6qt8w4qfHkfmrjZSxYdeCn58wKwAXcaBYSXKeJuhnpoAaHSBxlNzONUKMW9e3KOUkln8FO3wK9Qh
zjOWAPiLnhG8yTLp/VFdxkwnrXEAHcrOcSexaBTXiHWcK/vej2U0IxYBms4zJurJZpM8BfMDb5b3
MM41GUTa/oth7NeaDw3FQ51bMwZHWtudqnqetOkJRtWmS/jiKSwaSpGJfFd90O4CjKCwzKYrAeTq
CFogkLEo20KBLZbFVUPGtxHp6HKDJbXvc7kv5fpHcexrvsG1opz9/bO2Aa+l4sZVUPG3IPIlQwGS
tHnSL54jX0LRPI4ap64AE01xsLB3q7uBbkPylqtEsISqYOZR7FGPIdJeAHd9Esb4sesZT1Y9em0W
OrztDCEt+iMxFkSZSnZqvjPc+ybh1tyV15IGC2RGKZtzP/PxdGa2JZa8ybElORol9aDsCsh352kp
+99yWxxZt6ZStwCa090FRxWs6gpfdiA0Rag1V8Vu5ZXNOmFWRQ8ZKPwmo2UwipRJJpi7ZrjPPCuE
3rN0ZK72xMgMWuxEtuNJS6gh2xw7swQp27LmihEsQDYMVHpqzse5D/f4iC5pGeRWLuoYbqq5YRMq
d0rfMnA2LrqbPAD4I/y4liJ4bqdjr8/oGbTwrC+xCNmCCcTrD+g/RlxbGC64P3jdWCCWa7LUdcUJ
eeJebOD2rI9YAlmSXPQp6PUnUa+7JxylCr/rkF7M0wjtED6zatCxpdYEnstj/i2SWs9iQcdCdFCR
aaP/6ItGpwW8XhLTjRka+u44SDZuw0vf5kOA+MwR4xb9x5xPL71rhjUGxeYjEEyjVl0YFIc/3hep
fD33Fd7B+RiVctHCtM5AjBhwB9XEw8exFYBD9CxOo4crYr3kJ90PVepcxxMtopV+oR9qbyYbkwTs
FggX8CnSacuthhC6TLnZxcDeCSI60J7Lx7i6FoSjozrPHWIgAwcYSMQJwgJZUw2D+Ck43sKmQQQR
jTyTyiqOzrr5EkXnxVRu3Bczz/LNb53hgPP33gH675yugPUxpajvIvwY7cPwJnijveuZlztENwC7
0ceMPa6KoPXDoTeNqU3KBt1EtM/juTjlkMnMUwZr88doBd4wuG+IIV+B+PeFtgr5onskO2+HLjgT
uselsyL7VhefSt0P7I6rjDzS2jjMxOvn/56Ta4dJD/Kfbth8ttp010vBon9BRCeZLB8GMM2ALB1N
aDBq3/2Jzn/VXeI2RMU8xMPOYWZ9lwnp0PkBBiUxltpEGjGKywcZS1cLvv0oHB2mcquyFLZ6UTC9
TlLoA8kqCICYRkttDZRQQYY0xIjBAb4Bda3jG0bXVprmVkoINjlAsQJnzIxb2Z+xUzC60X5LrIOj
5J+PlFCo828Y6DH5JyFN7R5gUtu8xokrbmBZqJk+piyj9vrayVk/TxI9s3rVBfYxK58emwDPEB0m
jD4SyF01OYsdUykWD7iE+HJR0U+GYKOEvvFS9J484Ow1qlfZ44KwxP9OgMSPSeg/eWAo9YEML0zD
ThRxAkchW8fqasP2wQFDXVW2ruVAR11ezmM3UWmRD4B743mxxqE0s19Jk+teyHv4I6caPbeGmFdG
QmRFHsNEAPAZ3M53MFxA/HT3DKuDdOAcvuvC8QsbeF06GbaAFyKK1rirEw5H4xNhQBrHWzbp2JsQ
/rpndZ1Ygs6TLuSYmlkHEswmzM69hfq2/hkFQuUYAYaqbGf/xznnYCPGHwCLD7QUghbsGj7xLcBt
oxOloJlJjNY+78cvesW222NzJtaNzko+vjC4dJNtfq2rjIE+ai86dqUGNuGcTxvWQbqe4isbGcvs
0QpOLzkV/5fUVLLXZWC6ismyhFMGtQzQ9s2GqLbFjp/m9H03MFXAqaKYnbTtlBV+TrpQ8re/krIt
/KGzVxe8xcPt9rm6+JSsTKkJ5quDXq5YemGrDDN6m+ycPLb8US2P5pXjmm+RZuMBdGzT3C9OsM3b
RfqQI1qCec5SI6rcSH8JhT10091h17wIngmPdpVbaV7d1KlPukgZejdbcasOxYduia+4FEHNREUl
WcCcU8w189riM62mcutd1xODcnG17e+i8+0ZAvy5Tat0D5Qt0sjIplAkNwGM0hzkS0snDd8/SLbK
i017d/gNNEu9viN/YmKKWUls9xMTPVj6dPTz/hIpE4ilLDtIFeIIUj7Qto9Gx1V67a8+/0zlik92
e5SxclazZ2eKCaPqAlQEA79eVkW7TjDo9E1xFsCYpa6L+675DCXEQnDBW0j2Z3SUsQmwPaR3S90U
7Nut780wkeRunyuptNX8encTEkCrla4Uj5iDNYhhfVhs9SOrWAJ/cC9iLAMTpyQksm8v93wbm2P6
yTWqrb44LTqwFGiW/KJyJye1k10azMHFbHBqj6T32lR4rIQgHYiC1ejb8jAngBy65dvEIq8GRjLK
4yMCM/z70ihZAVOojqbL1uo1ji0C5vJdWjsCAxFRoGwvz+ygmy/Wnf9tjZxVo+J6C9i2xmt1Gd6K
gHuA9TxG24TQsNdFdv2bKCV4KFhsT9bkLQwvLeQpuX5d9tUxDKVBkgx8iQFjyE+VLxwKhlHYAUKl
rqtHPP23iRp/iuRRKmXF+A21HeboCx2SKDJWZ99vHMxGYGOWrApxNYse/v3i1XEIwMcKgkjSQRkj
Mz3eqt0zDLQVP+SOtnVPNMb3lnxZaAfRe/3q4HgVu+g7wWmuhHPOHeJWHSxMnvJ1pNEpE2JzUyOT
I+YWGrfg5ZR9wuuIgRkXWuaKRQpH27sueTqo0jVvVIPMjd8vaaRrkdo2h5YmluDZDnn1t45Ns5/6
M13MQQ+LCmlwUHBTaxZRWQxyZxBSv2qs3pLQyE6P9IMgnTdphfNOpjN7famZhKDKHcZogj5eAFjD
atM7mUV/LTtj4/5wq5qdCsmTx8Ii7IW4hWQU2CzqWnZXQ3xA/rIl4otW2yVvjZOmwKwBm1cojwjV
XLjnjO8X/ZuJFk7nArTo0vyZymm6aXXTDjoTCU9uiHNu41+vqzIdoLPpSPHqiAumVMUuwS1Ji6GV
NZhCmkJtY/Rdt+OMDvEvFO2bfg2cmb3ftGt3NvWX0cBh23lNeOUSS0r+4Q3Ce0lexPziE1IlNrgI
t/gAqzRMw1yAQwUHxiqjqzo45dtrwFrm2zW7jfr/8lFoeWLio5PG3XpQs0656ogZS3jVovR/3Mu5
yhWg3nTCZUSJYDt4upesS5g4H8K8nOH9+n+vhjYeSIM9M/mLomcn0jRoTS6XY3Ejpa0tdTZewJmg
6g99Gh5aGn8IXRZJfiWooopD0qlqEMSglb9YJ5qdY244DRgX/G4QK5U0Faaae2cYFy9X8d57TXcy
K+cW6Kp7c1uScdL0T3yE9KscNa33OVVh6xOtuYaEo9rzTdqk0vqrhWvsqiixl7rvUcWoaHFb5GlK
v9hYDcGeIscGDWsUQI5SyCiYKtjuFgvUGtPH8ijD8c/d5DQotq/WENpmwoZ/qujnZ0thPVgMtttn
ujip+Vie5Z9oMRsZDFNwLhDhYWDxMpCYOQSIGHj3hHW0Z6acFBGI4jWZ9neAkEurFBepxYWQKa0S
EW999pfwvd6aXNlrJ2oeElWaKahOER4BgyUIvP6yAU6i6FlvjsPj2te+xr1Rn+NQ5zDOeGcfCBmH
RnQbuBkuzlKIA+G+AaXV7Rq1c8wfCrP2iyCEb6lzY/VIQluQ30Yi+b9573qRAZNSG+z7LxOfgp/a
nsbqBpjyv+56uQmkeKKdlik9aQY5UO+Is4m8Ax8pefQrWXJx9oEu+engNbwOQSgh2AzOtF0LraST
RHPHVK17GIf0B1+qaAaK8qHzuW/nK3Th9SyfW75DDqIAu2GBTLDfY6bcDS7ijzA6oQhCOpbZV6tC
wYBjzcPPx9Qbf5u/+OwJvn7aKKodf3E1U75w00IhuKXZX9LJpftUhdMZ8iIVv2LCHZJPqlZHww0Z
B+pwy2OwUV2F474i/Ffp6pFwX7vLpr61dtOsTSh4e3BFtHsIduOjN6/LlljxZypZyBS/FOaLoImc
JRtiNApK2eTOa8+D4IiuGL2aKqfM1e5YRs8DWlA2EL3n7vPG1ORGTl+TThqm1hlKfSWjuBwZEsm3
BTnFMwJ2dndwf+4jYWiabXzuk/ow/oWwZwQ8D7jarO4Lub0EFeg94EscjBzpQXhaW6rYm7rBfixB
02q2bajfbcmkiL1CajtI83+BkkKsanCkErS6Sjj1F/UU0i/QN1tBx5jGzPNF+gju7iFecNTWpy6I
cLKWclQ+olkYXRpktRjnClr63GImixGJ0QBCbxIfvkUUsyT+tg3aC9txlIET2K4BiVe+Guii755M
SnyEwscJIxb64zb9hBgM+ItrfHV39REK/WPJSPju9cTFQMPXOqRAWy4cOA4uo15WCIZb85VC1BBT
0heJm/BD7/45JiXVDZfbA/d4SMrBqOqLea+ZUN1sW19CYapyEExCeorpJoL9ip3Ix3u+c9QKIzmf
QF6JSg7BA9Ami0UihK9rGBIVd0LMwcfrxoDIL7170a4onvV4OvrDMQPS9migNtYDtizfbxHUtakh
OHg3B4HCpQ/0DuRnKYm7XCZXYij1MkEHgmBW9DrJO/QcNpuEuu6W/YdnyXdoLvx/rUUBCDC/rOu5
zCybWeyX0cDgn+NROcl+lVf4z5OxaQxc1G5XNUxJR9sCTWVIQEQHYk0QQS61EjxuDs/o+J0UTWoA
kri0MuHsR9gp0nnDL0S86lRcL2fwrXgPzDfTnt6zmUnzDqAzAWk9N2ebpi0Ht4oG+hexlJMDe64m
rFiRagcnqL+nDkdpoXzMErFql9ptI5tbk8YgHdXRA0wNZUqbtcfWYiK/6uL7UEhaEyTezyIWYrnC
ga/WA3rnTDoh38aCisz5CeIgFY0uKQSeVIpNUpIz7uxgoB/i4HjourM6+qp+UeMJcXOfHjWbXAIH
2pxyzW8/IegQZIxqAFOSPFmJUqRqCMVW68gX+erPIf1f59ieb8QOeS+YL7pr97H8AlAY8Fv6uIej
ymMa33tSIP4p6jXLQVB0YT5+yZN61rfPMTDtX13uGMlnU0nekiQD0OT3pnb0BsDEaxgbGadRAgra
gpE12r0jtnPuetvfuKCjtLSh4T+v/ntNRNP7FdlSJx4qZH0Eub5VP6/r7VERcpcL6u/WHGY8Kv5A
7C5ugw8VTTfHaoo+nRc896lsrADlcGcQ2eJh61lsTmlj3MT6iLkIrB7W0VB452m6xunfLjow7Hn9
bwAV6UL0e01+HkJfdmoUmpAYZDv1EoUS53p/w5YsZlSlvuOylIPoP1RDTB8ui9frFdsA9J3UIGsA
Z8dba2NZ4qbNIBwmlf/WQY8qIOnLE0EgppSwXAGZVCdj++LaLIu1GqWZSeG+Q+I4arBec3xXMZ+Q
4nJIgM3W3jYpBNMla20MYrgBno2mr8XeGShZcG8fhHQJvbhurLZaEsbF4h74iX6NabEKoKKRzESY
gU0wpRjVzyiLRo8MMGerxgwNeexxHYb2eBLOEprfQsPn5tBoSFttfFS390B3IwPbupS5ooBGKaZC
tKSMfPfByDufbJsdcHzOZEJh8c01Hoi1P8w6hCuwz+N6hit4GZzWUcEL/RdR1FuUP5b1fE35ity2
lERQapgbocpTsjvTT04uY+nYH/I/JHQTTgC+y5TddRIUoO0V7WZGi4ccSTXEkm2OyTpD5i7Ki/Qg
qXSTg9fa5mLzM6F+Ii1pZUPeSU/tv4TshoU9f++lNwpS446HRgjpH+VOlaAJTbMwTimvLremV42j
8xYLD26hmr9ejmjO0O0mOpoDNAFny4AvTqX8zZ8bfOqOGpaqIorlTZklFZShBErB8s5lm2vgZ6/i
JiCeobv1c2YCxy8JHia8Vk2clsibgjf0NRzkNGi9f54HgnTUawXoVpOr8JxsGWBYSJ29cF4wXHHe
w4TeIzl2Yc/5xBWosP0JkzKgoOvLhSplGg4qZoFyeT0PEqo2+Wyb6qrxh8uRIfc5yuwDf7qoxuJ+
MFcpMSGhUrtS1Ud3D4MaGweD+B40RW7IO4QJNYtiaZcQR7jbRwDze2tfvgYJgnBDCOI2kqZdYJeY
xDPfkrdXOl4wihFPmG4tu6yaCvrty5NlCMHUof2jkz5WEEcC0TKJOTlAw6HCykhfNuiprCFfCXkc
Kjip6wR5pWxrGDa0Inu6UJCKnMXoomNfHrqBvE6bTsofU8gk5CiMcPp8CaYPFFyrArtAzuaByZD7
VHSVt343pnz66QTUDJtvDJ0iRi03naoeZRKDgJUGwH5fRQzGqhVnVTpFA9dpVh4hCRTT5ZXntE6P
iWwcZ9SlzcOExm7T5r7xfuSUrSG39xEJ30MdbKBDcXe5Vu13hKBf4NSdz6YdtkyRgQISdQe8ay8n
S165Blphy7qj9vswd6oFqVI5UXkKDVBcCjltx5Y+N8WB8hBjotkOXVLNGv9stqgx3i0tbPJeFK5U
yfUzCejPdUY//QM6sen8zpyGA+rzbXnTVvtjeROqgPhaIoNi0c6gdRKZ0NEkrikfv8k1E3wFCdaZ
rKoEwX7VLCjeaLMjo2gFZe51q3xqbEAwskjv7IelU8glTh+W8h3775UAKn8WRyzYe6i9GO7h44r/
6TYexo3FO6rX5tmGvLmJBShiZsTX26p+llyLHA83qas8gUX/Q33ElLR0KzaniVrIbEnnmZmI7mYZ
yW8F3YRcT+lIs+J8hOWMdJk1nbYLBTJCbaHUWlNxtSJ1ygiON9Rx2VlOnKpVIIP2F3ZdfpKRHDaC
krEyGR8WYALiMotSqB/jtej9k06Up5/Ug0q5LDn8F2ggwLG1j1jzK6WLZagXm/NQFsAd3dYKNj4T
W37t7t2Pig8EsGKZVVqVSHGVWQ0/BxIIYw9e9DAzWbg6PBrnD3j2Tz8L3Oe551optzKoA3GkPNOj
HWKb+Z3WBrVUnphvUhG7q2EA/oY6IIztjYXvSlq2HxDiWpInRcDi0CZK06Jnw2H1qX33dLY4PDQ8
58h+WuVYLgRjNcRvxc2yT/OdrVFZ8touJ+FIAwkfMQ9bpauXqeum1Q5sQFf/r4/gSObul6LRHEWB
NbtuwSMkaardUj/pUn0tZ7VVB7620PKG1jgZ4nxgvjZsqzPrtBxLHG1CLFAeioUoKPVjeKX3E3zi
P8ECKivfA3SfEg7Qf9bNikNXTcwdBeKmT+oMHHSeEjRmX9yh0bKcPneWLHBw/cvFOPbdrTT0OQF1
8OrRA5uSY6ez+qwJA/7RxtF603lEVWoNiOXO7xjNypsbiZzGpaVrqPsb21tnYNECExEF7s1YQA6P
6cCjV7eLD36a48ZBzj6MtARMsI4PgIybHHPiKfdPx8lFgoWJdHyvr33rOgOGRXrByGpGzy0KYBNH
Jk5BpKdK10xv0glG07NQ2WmXSYWcVWqwvmFdIwygcQht5xfDgWrWk8m8/uNHu0H0Z38+WYTD1L3M
LNKHFN00K6gy2R47lNG9qJj+rx/d3IA1CzVodmxApmbZTw/P7LJFzL/ivi2BwHqjamEm4Al102VR
WrWFdDbGr6I9gXh/bfpsY8zg9TebX9Dm7JGjnZwJmYPQdmtftMzWHkzede5AGEuy4msbxEJQAZ2Z
cIdsQzKBXoTgklEN2csQovDdRKIW3DNd663vFBLbR+e7xP+EgmeAtu/UKAPhxRCtaHscH7fxAlCC
p39QayKiCL0kaY8dnEvcoZ7PJD5N67Zo5xyqjb9RZVkmYTw0VH98aVINeTxO+ndbXX3QhMYL4nx0
st5Hdz6MuhHf5fEyuBfZgMggEPH81spBA6taD1VbFbruEdBzOz1HewM8Rx/cEs/7cuiLH3Q20QVS
QAHT/a2qBeCvqmcaVIono8rAjTflXotE/6ZhvYHmivUdJ0x/i7fAwwhmEvsUAMbiz+2GoQIz70QI
MO57C6iAdSCtyTcl9VqYf57QSREVdHoFHGkiAdNMyxeCMj19dngGNTJdseK6idhxjnHNPmnFU+tU
E+88EV1548LxuZoq5DRR1ranOkQZrGlgWkU/a+DRFtrHwqmk9JvbiGcngOJduFdfZHVibC7j3zAM
t1cOygBWLNy3xYbCWnJMOiFYE8NFU73mLDyzGdTeoHIaI8RtDNFpI2iQthmE4A3C2VP67W34ii+v
pOily30iaF00l5Xt1WfswHOKimrR4GWDFZ9DrOlpl1Phv87nM39ePr6l9dCGbqMvcVCZtJXbx/9s
vLuqOd+h6k2asyxtu6z4Kz3ToNfFvT9XKXbqIjP5LXfcvoGPvgwoLgmUNt4NfJk21ntcQZl2DrKk
tDSJSHdnz97BnzIxq2HYq2Zg4rArkQPNjIXC8WL35kNaHCgKYgJ4VTzclRN+v9m1GsuH/my6IMj9
ZjeDyV4kNWSOtwIIv6/aQqPrf5Ga/DZjgsP/ck2YLQGWKCrrraVDd8YEc0ZECO7kYLuIMCzaGWXC
pyuB7tPTa9Bry/uye48IYogrgmKCWYUkT99mC+iEaM8dIQ8yBgVBh2ukc9FcMx/JpQwtrVFJdz4Q
OB7JkDmgkmn/7i83/uWePg10Rta7iPQk0xbLFd6XBuvBqI87TP8KIRwoP5roc+lww1HnAgPEWcDJ
R0ckrKzENiTwVMs4AQhlvWhixHB+THQPzJfaog7yj5mru4mrFURun21BjPWtIjHkaXHg+paRx+vY
53rfzTRX9ecw8c3/BgjbLwv3kS46Pd/C/aSsOclkYBWoyIdWJ2oAhs/8ktZNnufhlRZIx/hQ7mm2
tPCjdvqYTPVvBJNKGoDS8l6+BxcIaFtsx6gLQb/c33lRHTRBF6h2nKyMPjSuFHTTDyI3EWEnUWWa
/x4rjdRCX/DEbu87YeH5Q+tXE7D5TGcwO2jece6o7PnMqnNqxqkevMwL98rHqO9fF4t6UidzPdSV
waNbl5uag3AlHu4zjYJpMAVDLYqPmRREsDzkIM17b+HyLQgMerQmvUaqgsxO26eQ1WTpjQfcFpOu
IX1J2UYlrjemSty6FyjjP17FKOTrrT+yoEZDbwO/Kj9QGXsPmFwJ5PcX3Fb6NALyYj4hZQ7JrFu9
1FU3WkA/6UPVq0Zretl4TF8HoqLi7+uvfEA76q02jVSth+V7YKq/j7ZSBG19hPShD/mc3GfUL7b8
mteHYkBmWL5FuvGz82vCos5orWx6P7aeRXSstYHVt09kZoaOqQhAYmYwAX9d7TuJS75ZzcU9Oy7u
lK9tX6mqmU2HraYhuzLB9RNB22kayAImmrIyKCpOOiA3wrOr3EnjtC+xrohAinPGBizzV90vh3la
G+QbIPF6UoCTIVcyE+KdkoHkc/Y0TluBQJToi+miEkbSn/psTL3rsWnUNRsMb9cEtVA+vixozQgH
K05IzzmxvPAbxEfMnZXHS3WAmrk5pKJBq2IUjqLYZIKLcy3r88AQ0KIGjsflRNlJHx0uTvYZKx6e
rMEfN1fDwM1lPX4c0358DgWG1JlAG+7KtmrZxXBCTL5iuDJpwStT7sCcI8+IiuMjVy05IjdQFwmC
+GQ+v/itLqaxJNft022si90891ieuIbJQRPPgAFvM52qQH8OblnrFthoQ61RZm12fjAChh2XtBxI
UP3rrAIcP3S3xxb0MPGKUCA9HuKmp5AehjwZWlvVt77phOvkDiNESwwCtrvM0YlVFblGrF08ShjC
NxoZasmPh0WatXq0jglR+lhfQkQmJJf9Ehh4ivMd/R6jAzoWPFiP55XvhbMGj81DUiuwZUsgYM0i
++5s3EHEsDztCcQGqXBDv93wnaOioZTVhYAyuc0iT/yFu5SCxCa3B9iMmubPF8zkKWVN3NawedN7
+IRwlyi+45SiIYY5L5DJMLaGbN+Nu2YW+v72A3Ek5i14Iv0JVzYS3Xi/e/u4xpIJWQdaZGzwXFw1
aHI5ScB0aA9uGzwwWwb0rfSOIfE9q9cpJ3YdoVUcV6DKE+YUG15TW+nLWc5P/VNQKL6gLMkFQeRa
ES6d49OrCQ+utzVhtrsbej7bCy4OinUwzjx4dxvbFS4lwB5CCJVB70dAcwzybOt/Ug62n9IwlO16
c/4VR/vYOav9XcU1COktgS41ZaGCVvRhhnoAukPQXSxXSw5Li8Fx0Adnf7xdiM5DuAZyZ961X4aa
zPTsINxVy9WX/6LedSKblwzz3LFYCh5tsjlYAJmd8j1Mudvsv/SpUo3f+6ZkNGXTgcS4e27pnIqF
jUZBcNeoH9qaeOm4wbmD8lM/GcFyhW9hkl8oVyffo45ZS+HXmiskfY1Ed+Ycz0E5w9LYCugR29py
/OhD5dH/THjUueUx+V5BX3XT7yLnPqx0QOV45So+Sq3F6/QuW7s299ahog9fbFAkDFrt02xcl4dT
bQC/tsWP2UZv3Cz9jXjCTRXMg96fk+zPV0wVg0LYQ7H2sw4hPUVXy4FNUbylp9e0FkvmsjxNqpC+
7wI7W/A76BsO0yIXqJ8qn+IIvvIQFK9awSIAMNSgx1DRoHdeQjyYWCpsGIon/PMEgPHAkcgywWgF
xBVMisn6AjuWlVu0SadIF9cu0tZ5lM2zTyXaiypmMjk10J6KHusvaj7KKQbS4Rry1M+4LXBGeY50
0vcusWhX0MhcqvqZk0z6DNKfk/eNKd2O9Sr6CGtphUbMW3h8LuSmcmSlAVz8QaiRBpHaprkQPWMW
YshHSObXCrLKKFBPNpoHpUA9Gchs1UwYJ9JEAxa0yP+bFeQVnQiS4KqfAgcjZUlr9F17g40XUlvq
RWo5arWS8aLw7ICh2xrKWECqOKui2AeB7gToM3DqJZenQFzvxO58DU5AOqZ8cXPY/7I/ZnXmN7TZ
MC/ureZge/yAv+FkZCPG7EzbJ+E7BHoiLHbFE9aPFDR2CDc3WtjiekPRQP683qQAL1FTSsgX+lrX
J7dIuVle9Egr2osTpcaCyggvwN8fEjAe2z01/6DKUlTuWV/8jITZprg41Nq9gXvHwVoDtVEiddcX
lU9QCggWtlfNbivlbHi+w5O6RHnHE/U34pcgsVLJQopicAynccDjf0d11BIi6leLlpUjyjYojRMD
ch+mYWW+UTtPLG56zId2rt3wT09/Ulnna+nkvspEw5UGG7kP24xyTgrSk2KkLWvtTco06ruXQpr3
ppCMOxMzhDNiWws9gPKLL21P19TLp+40k7YVdp5LNuoYp2XFs82G02HdMNsA/dTJ1nbK9YdZnNfh
Gm5AMDqeaN32M4CvX3UwGHkBszYyMOnEtzybv30WtIWB/ArZFFlMWMBCRSi2QCTbljBEVY0gHJds
oz6whUPiHuTfKk7gwXt29tkTYZlr212jUtiRlBYvK9lFZ6flxOp80FpSgockIqdLOLT0fe1QVk50
5piJjkrEJuvAL7Aelcj4XJoHYnmJvYyEj7j/lSnTKmMc24R5xAOwFuhyuvauAy3S+0jB1IL8uz9p
Vpdt3VHhu8vi0jY8UhctaHdEcNLmQ6qMAwgnfcPc7c2EBnh/SD0ZPKjvvMv6c/eQ5W6MZjAuag+K
SlOL9rGUES86sFFK10+XRfMZYR8giAPTTeYQ82Svls36z28lPP31dzQFrhWDllBSgfjWvchKX24K
kjR/56cHkwC7TLDQEgywpht7kQa6711/UjyF7bn1Z75LE16yUyEqN3bRtf3UAUVvNqs4iHgXry79
jivcbq6AiZOEb4C5ifZ2Oc0hpVbS+uZ9+z8sujOASjnrBkGvlyHUgX2NYYloINWE+zTgi+dURBSQ
YTNKW0ZizkFrixZ4c0L1tWzAnB9gH9i4121Cb7rRYZudp7r/I2xqkcNVNiU54PSNZXfUPuysTF21
BBuuiXOKheUEUCceM0WNdv6dNhfYe4gPLDsqf6KRa/jfmla75owPY7zaPR8IRSty0VRWTwDzHvNC
k2GjzKN9UHJ889S9iZoSxfaIfbrsuBGxjASWVcutLbefKQ/YVH2hAzfkqsBtQKaaE6Br+VlFcKn4
8cZP8act9TO5cR/YAUuxkLsirla2FgLGPdu8n2QMI5erzO5/RvP5C+Ixn2qsBOxKFAJeF1iHSuTu
BVZJj7ebj/jafVPMNRO2uTdv9WX72bd4bsi7u6eswP0lRMJK9SKRwsyFV4fi16ZFLbcdGYh3JIPW
OURCiMnE42IU51KlWXfkDxOrYC5/BM4OjdUECsnlrw2m97tYr5KA9q5MSMxrDCzH+zLmUGUXbiHv
V1xFk9iNjp3d+/blP7mJAPc3/9izAquI2rVHu7doPJc7V7kN3JmwEg9OMvZn5f1VC+snygvG0i9f
revFsq5bPap2pwHfRHC6QhZdcLs3ypBa7g4H3pSudW2IuLeplDlo8q/WxfWtv8ZrBks7zxJiLvm6
joGo33mtAyEdi4A0IHuIdpZDSbWh0qsfZWttUmGt6Bq9+r7tsQuAmUCWC/IG+uyJuWnesObzk/bg
T6s+gBAVmn/joIOid1rLhd7/NzQ1zE9+I9p5ZnQuXy7Ih6hDcfIqZi248RZnVaHrljkaQ8rYH2+o
dSSBWNx9Qqcr8N9o0At/oUzR9Yk4dF93RuC/OxbexOpRPLe+1C/LKYglE2vvjs5Cw81YPfP+Gxbe
iOXJaZ7lCLhXIFIexKqfGgm3F+MFKHchI7YqVyUZAWn+2b5k50vUp6tnejudCItT3pgp5+WoHRWt
SwFH35rOwPXjkJyUAhqcVoRP4P/ubN9Eq7lZ3hKorj9drwqHk1mp4AGe5/iC6labp8BPEbgVYgFS
WBf39ncGTEd0SEffTad8VW8GCza0/p0tG9pou50FHzjXRxNQxE+y6dR1tjpe26A9XigdgEjGVMZp
jFkxDH2zc1h5ML/XgsaEVHhpVbYjWj+oD14rJxbcmjdBYTV6WUSh+ApCV2fh9/lZk2/CObxnYv34
z2XzLC7GivjoiFGxYRS+jtBahNgkVisBnDyav2z2r8OICoYZXFSptjkRm/Zculhiu5aiYAcGgjHN
JZjgE073rpsDwGJJahV+Z3HspBCYGrOkVqaagUc6tW3Mm1HOexmecf913ZtB+7Z675VBQoH4lH1l
gKXyWHkHdnSuRHQqnktmdvKLP92wFHtoA8Siasvu2eOP5ZsCH+iJhQzL1s16UsKgsKkH5ui6Pilf
TF36gU2MCcY2bZYyT4FKDE55GhCOioe+DjUAdLRy4wKO3xYse0eFLkq4WeorPDAZKW7yvuVqnIzT
EoVAglVqIuYQN+dKlrxhMrDIDHi9TXA3Pt+ny0MNWs/EfLHeU+dZ7L25WtChap6kGlo8zxaDHejo
jefyZq5wN4L4JzhE7vbZO2NTqRbjuINjyEpY2YFa+I16MNS8P/Y4BcvlWqzc8tuxp2RVLpmY6n6T
16kVnaauYN5OBontFHToBzPaA4Kwgv1vyppE4uUVBJT95a0TnTZndhRxLiSaV02ZT7u/s54/AHqx
EkGMqtyi08BbX6ohUfEBVS4nGKRv1z4AglM9X8eLRPwXAJxK5r3BQQcQzKlZMcZeN9HtqbmG99aS
Qr0TJ3GHhbAagxeVI4YfgEh+Bngri7a7KK0zijS4Mx7ftI+B/s0tFWsqRv8N9GwP4/xGTGjo/GRT
f4vDEOJnNp2iHX/4DE6jI4zJLk8xgqYx5BPGQG5GfV1idqL+e/UEywzjZi4kysH27ZhSbiQx4BOC
BpxfPRitvtt5FZ3d1F/C+yuWLTIjnmdmrPGfs3LukvjDZ+pFJwu6Nly407Y3otGGS+wRO2najSVT
D96mS1NcK3d/xVVqDEdHwl3EIddsLAiU0Ohy3yVcgLP7MpLP60h4HFXLuCYF/pbTRRHPmZrMVG6x
TLH5SawSdBh4s8rB7U4iK7yl/TdD695IhyVHNuSQUB/aIH/i6fZ/dNX83M2BEnQMcwZ55fuf6WNv
Xi3ho0J+0ReMuFC8VnxOanSyhNcy8Fw4NIEBWaDdVJZtel+NFw/L5UfKB1y46fQajdzBjtl3F204
oUB4zvzi/qRVQGFUCCUWHB+34AdVQUWw64/i6AWROR0oO5OqMjBIYpfWhVwPpMyeD+KWA181I8Cj
XBj8OkbAF7NtzIl25NOrmoYzvNmKIda4tt5cCqhLDDrNg8Y0XAFEXTuHik/Im9AZUkJI7E4+bTHJ
llyYI5p3Fr5KbBjviDTkVF3637c8ose1FelspsAPDYp2ZVyEZYk8CFf6ivCHlXRCKBp1RA4xCu3M
pJXLwcfuMlvskqxNYn1ZEGg8rwFvBIeBQvdCBH2onLIHg7o3c4XCIJBVOnacpXkKjMlPsCFUY+Z2
Ctpp/HV38yxCazZOufWv4FNuAi7+X9oPYBXs/oy28kM79SIwGOeEM6xdoW0nsqkDfbs1p37vsBJA
PQhMLLx7sCnPFVmXyyZnvYEAJS1DKcoT/E6xk/uWcpmXmaLeQZMYe+5HNojVYB/uRLOHGBEffv+f
5gdrWgk8Ak3Lxlu/YFJ9Tcdhn4BnzBUZyFG118kHNNAdpqezyU1PZR50i0hTl4ycOZI1rJLXRbJW
ogLoT7E7tkv+p9YzwbzVu9bdwyDuuALifNV6Bg9aCJApdmIXLPKWZZHVz1et7caut9wAPwhW1/uu
qN9pc0GElxrypKoivzUjl9AjyrCcLmhBrGySXqhMCErGpaTQOBY/1Ha6UX1pjqcMJsAy7zN3YQXH
bC06Vv1H30cDnZotKfCEZdhdvtk6QqMZMicUWCqXYiJx+RlXMmL3kC5rzrV6XGJGFq2pQcJ6Za14
7ajDA2/6PgBArOVF+sZ2gF8O6u8qvj3Cutv99+kJ5n7AxqkSx+Rk/26LDes9M1ebV4ivS1lWIecC
EOjzYvv0+VjVhbMxkUVVtChwSY4+sZShw5bYrAYR3hfCRTW+do1RqkzKZ1WmDU4j64YrSuL39ZWF
bJ2IsTYRICsrmjK3u884utJQPvyvTpm13q5NmtrFzri4bBy9XswmgF4NH6QquFLhPX5tcxAkwB2i
UvTx6ztOcYlkmaKC7jjU0rz60g96fgQK4IGf+7V8h8KGX+7aMtMbnjRkNyXRZDsXcoYi6DXMlnwJ
736CUBQzkzad6bUgRW2r2epieTcez0HLsbm5f0BdyIBDv6PZ61SlhLfQgtRTGzGzEuX6ARhbZ+o7
Vype9XEV+/VncLG30mXH6yF1DkeA/XVnbZWlTP37kZU8EpGBMeaNUzetjEHA7TpqpSQ4cuc4VcNr
uZ3r5LQdOt0tdr8LGRCmN0bWI4rJXCztpoIG+9rKMpZ6eed0Sbx2uGzxvG42GZ+T5QrZMKjKGsca
bA1filzOEoi2y7EbzAIhnXQQVDIWoXUI5cOk5BeWJRp2WSSRFL2Ko2vHCbSK5GyxQl2bXuNwT4Ha
3mGg7VQQALocFhgzGkeRPRXN6QM8NFNj/GpbIxDk0s2Pwi35hkpezbkxF8IIoSBdzVFewerLr8hP
ZbtM/nH55eJ6wkvGxhIaSj/ewCkrD1JKHJZCWWaOPTiawVLvvyJ8Af5ZhIJOjPo4z/gwmZ+CINeu
3F14kQ7/1htz9KajxeldP4N+kDGQwmMjAtHVTBqd1gdW7GaJ7Lo0CKOsqgQBtshIft+poc6tKFqD
vvsSnUAQVd27FC6zqt0eC/UPmZdhaUdC+rM0FKI4YGX8P6GdLy3hfdLxkMr+pJcxOeDnRfSo2Wwg
sh62w9wIZzAo8hh2GZhvyQ/5QwrG+vBY8XAJ0gcX8+aRGHHJ9ZzbSJxvhkPkXX3/5Et7rdvLE8KY
HCgop0U9lq/FPnlGGZP/B4+jAL/hs8Dw3eZa1UMALGyazK/vmt+ibq8zUDfwl7kS4QxwtaG1Hm7l
IXHDcGMohf9+jKU+pqpJw5mxe1LDYOoPBDt+HkI9+k1BOhNmzJMZJYZQ+m0tP4uLcQce7PDZ8YIo
u+9oiVx4DAprOhjBWYb51wrty2RR1P1eZ0bQHx79+ZFEDQbziAa4mD2kQ/8r5M7bGNlCuhpc7SCX
IoGJ90p1R3Siq26G6QEtbywxLxzIMXvPlIh+7vj1g4WHk8rh8jzPRnbgVxN/Zk3u0R6MzPHPrQMt
89tThVHo/ryMeAJvei8cJ3Fic4O+cruwbCypsxcnSJHJmqx3cLOTe2Eh2GN9k/hUW8y6sUMR2tN/
clOZvJZwW+YTp8OkXYjT6PBmIwYBpFVlRZH5Q7cbWJYXDaQ64jsFv8o4+TIG/vMqnkAuwtfp6kci
ml9JEiaTgc4DA0lQZVzJqdfUak2VJlIOgtkuOdLK4D9kxXlLzaqzXjknvdGKXGeTYfyJ+E8W/fhK
FnDymjvCvPo33BMzii2Wo4zd0dzMSxYOv0MB5dE0WYAzoOHSvFgGWLu4k6pwYQsXaHKLDzww6Ug7
9zzJSV/7rdq8iR7uV8A0U1VqeeelfkMdREOCSCZzJ4ZE36srQUPLNIY1dZigs3qSZKsVbEzEZfmn
HSf1RjmJcLvx6za0eSa6EU0uGwudfZ/J00MgKBo4CAVvYk85SAzr6gxnHr0vsPqSvLEwe9xsPWVa
MSyODFmMa06tM9QD7klhTL06D719ojdpMs1PhBgrajgohqAZAFC3y9lAwJVQG22GNmFhJWxidnC/
stf32jBFQZDs0zZH3lnWeCRBQ911OXSB6pXp12wuBL0p1ohNb5zX4OlP33O8dRCC14HHFZFSIQLR
hOOJdGK+peHt3926U/0gWQvMrexObLA9xLQ1UGcAM06QMegMDJQHu1uLJTfnoPDugprk2vnSWM0H
BFm/aj65xjOpgaqjjRQa44u5JYEVGVrwsKjxLB3qzb0T9JOyugs6faLHhiVRnTXLQqKZJLsp6lgj
ZiGAbiMcdCrtIpm7kl04gzMjIBEPUsXGBkV9HZpURNxMbmfBwU05c2knLQDFsALBrhdDuHPENqag
I13BWU4cCxwJm19KiUkpC27ESxYjNb0rxA8uArDSr4ecMRLMBFsgaY55dbPbc7oiqafoDniBbkd7
xPu1Evh9u0GaSq96A9TGR1lcrvKIISqLkIz3EiJ7+rtLuGyGDDpTV2rNAWLw1V/KZhNRK1mFJ79q
rLLbm0KC2Y1G/tXpy9Pw/QlKRNOM7DpmNQSJDt3xfLAIFgzcNcNxpiJk3Al8zJ/r4WqVSYsRnDYW
Hdzjsb7j7qY6fKiuTN6akVlmtKTnFDBieGa3N9X6Lt9uqfOAtubzOWs1Zf1rOwTTTLJ24BSjMrcb
2Avo9Lr+m6B2OWmR3W5acykBf/Q/Xjf7sIr0DTBpA45SmsXcKsprgxXkvGckcFPcefBtrNa0lBed
PTOKEqrvQpTnMcq+WeyRvbIxSGhgIKEDbrQt5x+Lb3ULKRxtM7DA939vMHVNOdK1O/G6upsxFq9f
iYBqtNOc0sCE7k4FWolltQs/uq8fJKoOXVOsUi9NSjfoWZ4gFScLFWD428jkK/zcWSapXH5nadNn
fI7jvQTUrOgmcnMqMhqQgnOVckVAOH1zv2NWiO4pO7uMaQikYGckMJmYPTHoKHR4JjCD3jN1IEjx
6oChJRLWGJls4Ve6Itap30WBk7tIg0kKeZJWa6V3QlQgK/kLNhY+NWt0WhygiLHyjDPEs7ERo9ea
MiAoiQxGZn34NkotfWitK2NR2j2riyPEW+N/FC9/Bl0agrMQTVdveShC8qnSocoVYhkNm0hJh5GB
/MsE8fhYKsLQgBvGD5wqcSsEX95hVB+v6tpriM7q0bkkT/JKW3jZDIDc46auveeEWZPR5Gl8n5dj
tNYzPjI6sh7cHEeanr6ggfitemlOW05P4WkOE8rW3LLKAPONx9X5PSAMvimCsRzmS4tmFHXdF2Yx
LQoJ30BcLiqvTXSbqWcT5tHJBNyKwItQ1lEGTTXSVMhP64ne9ort4SQxecrOHFbs06NXM+Z4RDNM
VAA59sYSce9Womnula4rB9wTY7KWuDkXq6tJmZVnI3VXqbiKSVU6fFZe9bzhbGDIbGZFGRUJo+Ws
cvtWTg+MdxFhSe/YPpXkjg437IHG6lWpmlWQ3PyFx/t4rYPYjEMYheswopzu+8I37J71noz4QMU6
XJAIWJRebdjb4fGDvTGVCjPYL8FnmtfhKrkLz85pUILodIBdUjIfcYTD5J5rFexhUq185iuZ59JJ
S6YMwyiMN07L8crqggasxUMF+1ALBiUcuSQMrxvWPyZQ+NFt2Fuh/rMXKKUBf7ob/jt6petwEmfT
WKLwnozdw//drcQbpLGezq9sKlPAK2pxij8p8QSMV7FTMDrtWK6O/WGyBhetQk52sqtthPjD2OS0
0mCpCyhtDLt3wjDC896UUUlmgyn3IiUl1zWMQPws/HwK+1ZTcS7j10L/B3Cy3nV1Ccp+oVf9X54m
3MvKnhHN3LpNQbho8//FSSiYUQEXEmgCHzzk8Vf8XU111TnXtBiu5ntyMDQLQLgg678YX9eXmjN0
4y04MryEEs3pjEonk84Ip1S9Tp/gVNMuAb879DTRBTLAQ86heOh1JkgoD6EKrVP5W/hvZMdXCH+Q
rxZwMiuPhKHtO2sTOqhRoj2SAgGgnl7OwKnWsrouc+Kpo7nvYOmmCj+LED5fF3w3VlM4VoWQGEK4
g90e9K6A4tD14inW8djx3DUwbKVunIi3vH7r3HX2XhhOwROzvuELiNDseLr5FTJoEzunNHsxaxRC
dFlq+g8WM92soZOlGrcuwleUXvxFRTMwkd8z1lDBOc4UG13RLda1WA6ohbb5WuMaKUhElyqvf/wE
MeavcBaUxeIyjiML/3gSGAy4CJSgK2t7fuNCwtivMHp5vMm5kREhGh5NKdNeYblwwH3hAMw3AVY8
xjEkbS/v87txA0DPbHEsQgop1P/Q56T5wrPUUf33EzBN6JeRLKwkah0U3AklB/RAXxPgcFkRRhzy
C1kjeWQl19EcrUGH+N4/NEfx1w0uJT4FDHplD4TeHbctDrLJphwYsGBsz7IubBIdhjW/72NuqDMV
BchMDgUdNBe/rhQekxleIggxygnBjzbn6mU0g/QZEpYh3Ga+XSkdt020euQsDACTExf1tvl+WI+P
ueBhs8X0ZGN5fKI1sMv8R+29o8xWUlOfFd3fjl+KY4ouHQh4dwcAUQ4+QPH7LDXxXvF7moqKqlMZ
dlfszAaocA08okYuJPJ7GF9SNfyBdnk6mzc5TfdWT8pO6surHo/R42SEVwi/pMLMO/SmpYS74IL9
B7/7HurkpV9eHH24scLtj6ddt/Cpvm+y04Oz/gxt5cTzMlo5iene6fWgsHO+yM5CwQywiUp3c2IX
4VpiiemMaUsDMt1b3Nf2bV70vTIqQF8A1Z3syMI352mx2G1uW2O88nAG9LNHWGqVTOCWDz5YDx53
4XPSeil9+R3JlE3DuyUGni0lmtNRp/2YpP6nCHIkMySjxyGOuwRS0nOnn3Og0kkjkOQwxT9J6m5O
bnF0/LWxZDUz6bbbGcAuWaoGE1Ilxr+gkJ0w0QMBgo+/hh7ADOjXY0+fq/wTVkM0062GjlrRcgZK
VbQaKoFH/EHMr/bBkxiGTb5G8xQ7JW1Pla2U1Mg/YEW2N2jFIC+GNHksq64QnKyfg/1toKNMD5FA
ZrX96w3NzKbD74in5ZoAidh6OQLPKVoZogpZbywE79kZJOVYgXyCwa5t1BqXVU7zU4Lt+C1jb/Y/
/WS2xXbBO2ykomwgki2LZgMWDxuSdPN19jEnksykrORRpLEy9Hvz4J6WQom/8hvmaC6UwEedaMi8
FnIRABx7m6ACwoMvdZmVv9tHmDZaFfYV1VhoGZ5q4Jw+d0//tgZFyQSPAOaYsSJQXCpd6I1/hfBY
jSWPDtUL+ln3ArgXkRAVc455uoqWmV0VdmuwmpqT/ofDmYxhoBjUefkzHu/VYDufpGUZoCfxXXno
INLRlu2XwxSjUsf7sjaRwiNVJAy6gXC67eSPPIoxcQW+qDVhzxS3XkTC4qubtt3hYLvDqC/PBgUO
0AOD1lDeAlNRgHCRzmzfOfXExtY06cGg05b4vicDct24g6GZHpVgjDBO9An0rkH3MDtZfzY9lPy9
ho1V4RjqHGgzITq7VzAd8H7DMJwM8aaxkyqgVQFGwH7wivqtIOfdTwxlzxZTWjVT5+dY4erOntZV
PteplzbSH/4g3NUfP7mFSd5r4nlDUou1Pkcoy/j64RHnbZ4j20z5FzXK67DGj1D2DHXGUTLN7UMf
00sxhfJfWjG2NWEOjVeHWHL21B9Dy6b/N5sb0N2m/Vzrm6rAwBqG3MCchRA46LRZz1lPTsB3ES3s
TIPPm+edUP8JKmemqt2B5GTPgZqC7xDmoZR8UhOVCI7fUyihxEhhEE0VQb9SFr7CFSkdOCEQRzgl
PETk+H6gkzHtRNtUReE2h81CxnG2wcZNAiShC3RS+2RKSJZWNQj+SY891M3T2hkNFHrl62M595Rt
OAqyPCYgr1qn7RLUx0QZ8M0LqxNjt6hEnuZgEuAecOuScwo6/FnLTIKn2yJQ12z78St4zZq65U7z
8dEmRPPFIwq164ztjI0QDHrRogacl1LU5eLMVmAus/iJYpvGnXkjWAuaV9306NEWaxJ/rxoW8lgZ
+9evqR5XszGvgUt0xeqPg45CX7JqUBsoHoADBNKEQnhHfSBKoHJ7OmQ7tF3eH7YcsusFRLB3caPr
2hlxa42PvjqgR+KweS2upctTYqh4AYKTUMnxAO8brS7mfZUWx3bMR9R8GV+OVedQ0Efnl2QXNzJE
UZL5vhqG/A6VeukWKBNaFDnEfkk6RfZMZc/1zi7xW+7fa6c6lDMq6aqSxdgG6pboto4lrYmh97Ku
3ks8smKVbqoFW4iBHDQGtCRmj6PDx3cOFVabgTEVycer7GbLXbMQ3ViRfO3TPaTW4rI0u6XPfBCV
Pxysl1Fi+h/EcNbI72Ye3cVIBYRofAYrrzkYRU+u0LUYKV8PGetFvf0OqrPabFNu4rbyO8ur4QJ9
Op/p6yiPPXwf999OTAqXd1pPqIxbSbkS8vEIiVbyLH74Aay+ybbNQbZO+Bsyx6uU4Rm2w1+oj/VM
URVSXSeWbwlt7zKE0kykzQwXUnoWYgI2kqtb0i26ydI0IeDOpVCJm5ZZ7R0lLkDZX/jQMOa9CFSV
x48b/OdzW6CNJkeR1qI/OGa9DA1uXtZmBz21efDuHX5Vx53xVj7CMUsldSAE3Y7+Sq/NtjQtPg8A
KccSGh90aQSmPBz+xYK1YBuZ0nqrC0Gumkass/TEh8u37wULWCtbivlZhvULLov+03G+AvOfQMwc
mdTymO1YCiecVg7pEGJGL32vNuYF55wYDcy0s2D1YJgSC9AYWnA6QOXEh48vaEEMvokkZ7v8KgqM
AuMb9ewSR6h8QClmqeRuLKRkU5fwFvDN4BjhT7E7H26/hrXLm3h8Zrm/Fkwucgdn/ZqQ0bm35Pvt
YSSPWbET+7Qb7dUdglYqJs+7oME56jemrSsafehKIhYYhoGMGyhROmV4PbGIcWCk37sqPPMZtH1X
5d+vnM4DNSBiBLzesiW70yATKpq0Sh8fJ82toqo0KUUeY71RBLz5Myn9Y6y+zGzQaCWK0SbblvG9
0KmrkWbM9kr1p/KXo8mUBBkqJKHqYPpTi1tf+AMfdW+qL0MpwyXBUuTGDft3lvPJoehesm449xG7
DpIfSi24ZGWRkZK7Rn2dTdGnMZtjBbetGVwR9qj6XYCHgf4GHIR6qdaauSeYecm+HikyOIWe7GRR
cwc0GPSse6wBxyJsU5RMwVHBWdqAbemb8FcWVK7JCUvWS83cPuJ7Wpm2aWdVMPfo3ioU2voPxXFT
P61v7YlQvNNzNo88qUTgj5w0VUMCmmURj+/gAFVOzK5j5FIDrZpteYA+gHH0Ul57ml/3skhI/7Qa
AC8vK9fqpw/ZWMyPpTusMXd44OdmgozrcXbeH2Hz5EabcIz2frxEhCa3kmHMTWFuUo2VDjNxDNPH
8i/kRu6aZzZyEJe1WInvpsK0cQc9RlxZL8ict0aSUTNrOzjPtb9Ddj2W38+MrAJ7yGRbO7nsnFgu
eREy7pBfsyHAGiaHPO3EMLFC0GKjDc4J6d3W1csmJ3lRgeIA6KH4EQvrROonnUZ9+QX5DK2qWXz4
AO99k/VTu45WYnc4SVAOLtEmGSVREi4ev7BalO+Z1XzU383UNn8QeqWTIPnHGFATGnHITSBLEqt3
yWR8LhYzY/FmEc33PcT0QOABkbuo1bnQE0Dw1Kv2REohnbLpWK/yP9RJ9Kq1Uxfne6UkLLKyWfZE
p895Iy0jjAT+gwJ8rqUBg/9aZe/02n2NuBXBvsReyXSP/k+Nd16vy1hi0UiOJ/La+WqeDateUXbl
bk50qfdZO2DK6RzCKYUfaF7IdzV8Y3s95+TSY/WR1b6RKh7w+WCocyAlZiJ9x6aPnytyBlgR1b5M
h1ldpSlRpkk2F2Eizq4J6QHWyAS38Bx8yjCFmsBJyOl+aMYOqQxC0Zb6LMygTMxYzcCO/djDIpt8
mdzCKKYF8Ww7KGeJIAd3mcs6NagVYnKTsmdaHzj9PmPioX5RwMmrrOdKHS9S16dLNqcfO3bIldty
AF3YfXaHvKi1VxrNPApwHbWruqkOLe1RIu4+BkaFF0wTOzmy6VYXmjd3PafQP2LYzj3g24bupoEP
V2jhISItvrNq9zeJdPYA4dBRFNBrPYF47dgcx0KCxQaWDZsujbtjVjmHv5wc3YCXjJnElfrOR0wi
edtFyg9TgDDhOFcQCeiSzAiLH3A3NzfyPeS5Ya3WNP8QcNA3sTDg/Qv1e3uyjX6nyGzNX0pyCr0M
Fmm1z8gtM5nMsa5Y8U3Opu1ku6syplTuspqSGJ7s7QlNAyMnbuW6V7feuJ96O5r2spEjgaimfNUH
E+bhjlFZEI1eeRat9QtjqmNNyl+Mdl/1RPsgr6rdK9OV1cQQMdVXg1n8JpUHMGOsDTLiANHfTYjY
VMl8EFHfEM5NkyR7rhkU/FGKTVO5MqecI7SMTLlybK5ykmzhW80+otSctyQyQCp8MBB8uCSLX3J3
lvKfuMK4wk/N0KyE6a3qemGPCvHjZrJhW2y8biVbw1g6cj4bevpCQK/YYVGRue8n/pAPW3f9UPuA
rJ93SeBrcMfpKpbs3CLuhgwvzKo+0P0g8FMm2CqJVBA8wly1/pkuLCIt014uTBtS1wLUCpmkKV1u
lfZrUCgydhoBm0+dmI+XPONNmIpfCimzM3Ib9x8WUaQ8uAe9K5aTW1lGcnG/wdrtubG7hMNR2y7B
4xSqwT1N5UOaWDZ1GexkujO+jtvAoIGRHD4Pe1cwuLzmxF3sbXknECtgLitrSmcf4qNjq/KibBZd
NKFEcEp77btgoOtpymT2mQu6SXq5Idz12tO/bqlD8OHjRNNTJDRxPB2mMEHwt+2Y27F/XQpMr8JS
BmvdsTuYeYiq+hR+MUKBpCC35ayI3E0zGhkyBMXfQxsENtX+WFpNa31GMkfGX/fdoi1/gE2Et2Z0
KRFbGN1k4/5XYjsa5CuIQaz+DVeWKPGfCY7/9zwrLz5v+R3Q3KGYo5PgaC9uROUqGxF7trvw7n+W
0LyPjOxHASt3Gy56Ul5ZtwMtg7GeAo+54KozAWlYxRPph1J1sP80vEht3ZOgVVPKbnsvoSDJep12
jMEd2+ZmA1Di/X5gJfVEuKMu3F3d81uRRbidjPUGKszjD6USRSLAtT0+ANFukALpUf46tSJ1O5f4
UwpJUq5kkjK1mUWlfCvcAdm0kBFPSacwGGxbHINVguqzJBjogrB+mtsGxSHxHR29iphHWtBGQEv7
CzYx8c80CX0ux1cnq6mQRmeHdQORRZeJm7wl19yfdWQi7bQQveNOL7cjAhCY+nRYIO2QssP9bZO9
d3w2yFuyVTVBwedGAWRwOMDXiasU9trzj9Gwe26t/aV+GSIdskDKSynJJHEnuboM/NsMZZhwrD3T
jIdr8pebByPJuxELj+pjSdHTKSiV6sM0o746d0vF3D/XHp1HmkHNUHYtg35pN7UwuBVOnE3ONN0S
DlfbuxS/mPRvzuz/6XZQ896W4Eo3kPtw5uXXB0WPxWzfw7F5K7q7jXjuHMQxOvYkXae7Ry0Hm1QM
9xzmLYrCOvazFViagKCBhov8glaHlcIwiFK/9/bdnxiIUPyB/8hQALyTV4dJto2a2hoPSQvsYqDd
U/Fh0t9y9kG4E6IaxsPc9eSmdYIEvqYrwK2rOijLuQZ+mkkCkeKhEmuc47WA5V+abpc362oyL6jM
RBpxj/y37VQR3+Ir5fwAqbqxNXibDG2+JidYapXLZRnd7iSswY8ALorUFJj2R3kefRnZgbgfGQ0Z
9lubf0Y4wSNnV1X6YJZOkiWNbdOqFekAZzGj/YfPUMtbHTgK1LNNOqJ1MDF/n3SbCtUTJ27rms4X
mar1djvWcmP6y+SXGe7n0dtwKOQt8Hx2NiUQTrTQnhdvbAC6JfpmvvCrwVJMP9+p8W5GeaJUIrLG
D+9xbXmr/WWgvb9cbbWzp+0wRjB4Mhd/QbG8se1N/CWWr9X1YFka2vXfiABsf2YAH6K9wWikbmLK
pVyJovD1za4X5Mnf8kx+kKm0Y+nQsUso8VjK4CZrTF+MtK8LOiA3yjh2rvMve9Aod2+eAqHhnO3n
kGGpWRiPp4TCr8CrEoFGvZA1dvlFTlTq9CdZPnTlowAw4rSnqa8EZ8yQabCSIGnHMmGHeMHs72ed
PqGdSeVMQYYZdKnBkz6HyURxOEyisJkNzU+sMvQ1AHoy55aTPTnIjeqtTlzpOfwVhhvwx4/P/Fkk
63ITjynm9MhK5Kkwf0chxyvSrG/gnQhVWmcWu8o1yOeiGUFcA/Szzdzu8ZYtG7sgnVXv9XMC+N0r
kBra1/vnj7XwMG4TXi2Tg30Rt7eiJyLzvJCu7Jife+aUIhkyP6rNrmjHOvNxACaQhYMHUteHvURV
nK/jX8b26xZm5wfz3Tctu8OBJ8WnlY/hiMfr8gQGBsfh1vTwJUFCWvq8R28iGn6diSKi54ieo6iH
x0LmrHJ2bJ932kpob5h7sGWpJ1qgNKtlMcLfiZBpg3oRxVb+gHENX6UKyIHQMaobqo3QrS+TlL1a
pod2Vwd2nkggljdD+tanV+eDvMePLmdpfS+z01L3JSAaZ2KwHovOE1nY/Rt0cW++q8YhUPJ+8MgA
3lCRr2oPwNMBZIpHYO1jTBMHu6fy8kdtkz71yE196vd8FBacLuFjcPwJbNWDNznnoYxtT2dVtJhc
T8Htx1pTkg/++G6mjBZYDTQ0xPBsuDEiQ9BjfR1PeV9MYmFtmDYqdRpPD6kJHTB98KUl4tdTfHQB
o0q3ugWYterZRR9jjI5+J/7NkYyZ20C7QkVcaSgMuJ7D1WyG77j2mp8rJbGW/nyoNtNxyOuK5uvz
R17ztLEIt5kv6vJp+B21f2pUaHEHxS3DyaBTLe07z84q/MNpRP4iUyCfA/eeAnfzDF9URR21e0Ut
nn7k+xM1Nv8Mt3MclE0crQ2rCBY+fvat6eZfFV8t6Z69xnQLLFKxxQtZpLlddU85xT5WSrz+qWvy
+4NlrLiz5wlZtHbW3oMpn2MsPYlVz8OYwwO939GhhXV7lSg6W92sS9nFczhVDyD3Zp1dNgYKgLF8
ko56A0uJBpxrRDo1C0DIdwD46twnMGFNVFV7Eu4mbcj3o+yO/zNY2l2Fg9pdtRoXu6Tmv8zMFxYC
kFiqOay0Sel3c0/hl8MVjTVGzXTN2Eidb1Y/G4orer2llvtvBITqhv0WkWdNTeV/SGVVHE1y5Fej
YetVGC5tkWyJI6TJJyJ5i/Naa6lNfx+VXpZM3C6Re4gy/X7tUF9nxj7c4FBZAPibkV1qs4BdOERO
YJEdeF+LZOR6jhW56/u2AR3wkR1KDbYbZcaZpmQUDhtxmt8RcLxEYPfp0ilZsJAL+1PPKLd28+/F
sSpJwUowa9aVTiUZZUgdluSOsWEFHn4bz6xWV3amAXlcAZGhCDWOI7We6ydlFwLcL/1xgtQJ9JsM
raovAU+OAZcPwP6jzgP/y98QRJt4WFT93gkLN7KoCelDMSdtwv2Z5fpW5bIo8A7eZOufmxbSB7R6
ixgUuCPUEquiBGXfzUDFg177NC/bM7y3wipyLDeHWvbQliPg2ejPiemaKtCoJ5cyVrTclS8nujFM
po1Hyem80yMQhxY3sZQyxIt2iBrT9e3kZRy+cVTk8McmxDynztbVoSgQiha3500hCNshcVxII4yn
HvlDoFcR8DsKmreJEKeuxqi56P8Qm8M1V9nqM9cTKPYHKxkNSYYVzOOFs5+RsTjgNOzZ96w47Nno
RiOGAARiP8lMkxbr69vNUfC+ucb8XQyicPH/v3nuHfMJ/Ugi+GQ0xZzEmTuhBKHCPB9D+RvtjXnc
1kA8WmKPwcHW3zhZvnh3RdWVnMgBLoBoM08cJdEmsC/yz7u8a+8s3M+nrI7/CiMjY+oCk2yd9YQy
hDUmk8fmIyDN4WLhMJfRzuFSsnmlV2SukhuRA1zAJF79c0VjBPMJFHzoq50UYqcYoOhfK1btzpso
HKIzbRMhnh90RNu7B3KoGpsZSbouLdNb6EusSQ/2XPNILkyXfQF9mF2PuZqhdgP6ZvYIIjpUjwnU
DyxbbU4+1BciilShjoNDsVcQthVLg0+kGW+3HzXvvY9ZZylOB42t0fz04GHVF7qu/FeMvOiN0P9l
BXcSgPYeKl/LCfHUQObEud57H7J9/ZjlelbzEBkq1Q8QzK0sO4s1o7t6meUHdosZ7NOa79lCuHSd
goy3QNsgXRsBXDz2z8T1pukPR+yjHab+iKtmnwhotW0NfH6UzEjmA/N39DqItonTJloCKVy/Yq8b
ErH1qswRU+OIY6AX3qzExYxsbu92gZqKeqMalaL//xFknDm2YK4FztkWxcHORv1VoVW9mfNXv7B7
8R9IvPgmLXnbc4OEwwPk2KPqL07o2TL8Fuwzknm5EFESa8Qbwwws1ptAZRpt0Y2x8PjjNKelGW47
0YTa9gT0aqu/uASXfROeBbct5KK0hf9WDwr6XbPS6BFB926iRL3e4dSg9L7XmWS2ACi/41UobITD
Ad9k+tpeQxalm+ZNNrVLdPdvZDelI49uE+1lClQPTQCONeRAwvHlY/DBBt6ewChNUezxBnUe8hsH
BNDD65rCyU1YwitY4kerfUULZOCMsYqgyxKGqZECH54dVqQtxzjaLoKIF7vKij1MJy61XPg98Myj
xIjRFZd22ESfj3rym392soeiU1CazmWipb14dnTxSj+zcFtdZ5Mk0bwL5L64dUDNezW65GJ1NVvW
Jook8OTU0RgcmMpFbjkX8vP9u6kB8wqDaQbvD5hXITluRAPjpI3WhTgURhXojPEl/oVPQfZEcRBF
9kfw1UF5nL17UemlD4nLyL1zP6KN6Ad3KSrxr+22tjC9LTD9Vi1krKSoG+REW4x1UqpAZGycLM/j
dOiFeMD8X/l0eb6G9UO5tvAGj10t72Ar+4vOIeHc76gWPANM6XYfGrnZs3B7IV2iQ5Byc07tVMPR
jjcQOJj7qXm2tqwcd94wmEt1CUTeprVGXFxOrjTBcGXa9WHEn8Gx5XP52kHhvNlVHK1p4o4ll0re
/NeO1xkDBReCMGaj2vUtYGeE3fdec9559fMZgn6I2Z9hmPQCqek+172eiQ5j/6BV/B9Ryy08CK/z
mpj6Y28iRy2Mftx/Btj4OMctv+5IaKlU9Rm2E6NdQ2j8NtTKllGrB3io21uwBjUkui5MLFzUBBcq
+WqAHKcjp5Sq7uAu8prNiPqv0U6UBOt19OmjIhfpE5UjSKOu/WuYb31jAHSlGA1k0Vfo9/hFitPV
FVFK2iPi3DjlI5TZDNR8R542Twru/4KS/MJ3sz8EXR5BxOZ2+q5GNVxyMmXYMeFiILEvKaZi9W63
pLw8aZQKpfnaE5fy4ijsEp1HpvGPkdrhoibjaGRE9BFXHMwuE1uzV3gTEoCADd5faNL3tkiB7Gd+
cI1m8uO9AKvb5L2J0ZewxYA44cebbJt3GoGlBit+3mJipJCvdPiaqrK+95/G+Vn3/R+KVUpYFlYn
iGRmlD8Ta3oPbvuPaoAQthzW23ZjYB3WQ1X4JskRfZMOnKxg5xIxGNnTzrwoGudSEqkFA0uQ4bMP
XVcFqZ1KgPyjiw1JQLkQ1L0Ltp56svX+wsAeecjJP2ehEi1TiMaxZuYpbL1PjVCiSR6u5an1V40+
eg3KuqvXzB54V5ISQ89pFF9tQ1qaNSFzYQ2Ls/gJH31oenM+mVq7d5D1U+whxrFErNhKhvtu+ZsO
NqNQ+z1fLFP1fErWLyI0aNCUr+yU0t32SDX270VQkHrUaq3QcTUBssd8d+qZsw0Ok2da8H1czMMa
tKLP7jPED9p15F15IrswvvQyMY5yXO4qP0/wk7U4sSyKkf6sHCyUbPjFLB7SFNif57iaHVdBCwI5
TsPFfCsWDjTSGVZqDtFUY/cL0Rm/WK7GFvPkIlgN0AeRvqPMepMMSY43ZBtnzuiTwaI5KnUWT7nG
AIYRvEgjwi3gpW3v8+535UYsi4ccw9ywLHwe1s+66Hos5nl+FJ6p+d4S0IDYOsIalFQTSXJS7gP+
XBXSFB/zE9rxs4B4nk0NCY0W/Ve6N6ckFIR0mwR6ipTiB98CZvWldP0+u6ACCwNqGpj8OR65wlud
7NVUKUf25H6Pk1r1oL+kcEivkAZX51FbW3m9+h3A6k9VIfjz9v2RO8VOzwIyjkedTgPZLn1Wb9bQ
VxoGoeKckGks5FhBHhW9P53wzmWgZReV3U/aeBKAPktgcYzGVBMgph2H/DzOqZWLqKnUA7onsGdl
kdHlcrVZWFaIqSQ3pFJKSsIt7PorxOq9Sw9KSmH5ST7iriL0nu5y+Ucgro6NZ2yST37FuJUoDHjo
rRtogeiS2WUIFSLg46A/Bd5du0sj19F0wrHDYX2umbqpxmq8KoSL6WwNHbGzTWE8qRCeOBawxVb0
xwRKfnLtQ7uXd2JzulDitGDlukyDp1o0RzZDN0UwjSPn2RfcAXXZQLg6schJfci7MNx35U51TrP5
zENkLdcIK1sdnpltssQp5lsx1BBAnZsO6WNb1/bP+BaYhi8DsI22UF6+/0ABe+wbnV/8k6IDjOEH
FLQXpvH1uw/Iqwxt3gpbRQbz0MyPqllPNjzf9+EIugfbNPfmqamvR0OAKtELg/GSfMCX3HOqzM6F
2dFejYj5aYOvcjncfrOfB7Y9hz0GadUq1ZMAXhozS4Swl7EdKsinahDxgt26LoY9K9HxseCx9lCU
O1jL5bLICMB1fxKJO/YnxM0gfjhVLX2L+V7bmex0Jej7wndxePtt46kclaS9mWP2bIEL9GSIEo3N
KYqF4w7WlH3OOF4l1TwUwb8Os9nYZWHW3G1QFGswBlKGamkIjh4AxrOrxb2ssYqO6x2D1XHkZ2G4
sHPPwEp+k1BbhJDtSImJd85mYJMSz3D6DFT5GIMn7GUDa9Kv9SR8lNJlU8TVNpBD1x9n4JrqkzZx
ulf8vTHeomuzSYu3lpbBesK/bVYZ4NVLSKMShrXPgzU4i8FD/0jydK8zEH+NUdLifCpZdp+6JFQt
thGUQiV4WRRgiMKdZ7j0BODPH2ppIDL98j26Lc3xX22PK86OUvXxSDnFi8yYRVvvxlCkPVaeh/aZ
dWOn53K3WgWl3AKo5eYV7MvhubpynM7BOiIwhs3OruZH2Lcs8BIsN9/fA3rRuuywtbLwPCnbYseW
BlBsWDjFOKqIL7LPayia7JkhynGxMNWFIQPO1eI3FZIQx3w0m2O8JDlnTov5vFm2p/LpV/n7aIek
wmvF0G8GjuWH4/wXHjcSx5V1hfofENu744fWRMf4zUuGSsBt9gla0pbUohWLZUrhShGTvcOiCVhZ
Ym7UGlec8FUP6NKi4owH7BynuoS4gtUUx3UzsAeOst+hG012xcyhDV0GLjz26e8zC8qpv469GeUO
rFM7LmgQZaGIzNsQaaiX718iOL6PnBP2298Ixxkm20+iRtz0GQXmYk5/oNc9fcWP3dCmIdMLVlcU
khuRBye4KsVVV3LtcyTL8iyK2YZUMP6DaW/pu4HwNOqUO76ypAH9yso9bgSRtKD5IPbHBFoGTrqF
/lwZqsid8w+4BqOtt4A6iy7XPPJp537y3W++ZyqN6mCfBjiorKGJpThO0r+OTiXGMezdr4M06T0l
148CZ4o1IdhgVjmZmKg85g0vVHGT7J8kGZQ7NHGctUn6/1b6PoEpQwJfY5PBWOcWV2vn+irXSD0U
4ahNKoLsuQDCbwL2Xx7xFifXXKbZB6eGbOrkFwgnEX+cCzutysWTOwEquThm3pEQDeURZS4SJRCF
fSTJ8J/9R11/FtIaHVQ4P6elkuqyr2AcQJt3kLpF0Q4nWGO+q3cRR5eCm4E4iVZMkQhkPQ/C4fcx
e5eKwZaqrYnZUgRnWa/+uxm8YXWMCTIcQRcZeZ6XXAuZU0Pa0Pvw8kfE/CdT3UFMgBt9aUmYLcDM
6gHXp9po1JEuADyV4Qy4iz9CZDf9TAMXNXRvc8n668UGeDPRvYlHAlaBogLVjCRvhjdRfY6QTfxk
NYlmvTxEpY1K8CN4yaK5lOEQoQUV61ojeOfKQWLp7P4EOuR0UkVw93wRAZBVcAkwwj1aTj2xQAdb
IrUAKCWiRshPNLemNiknB819OF6M6TUTSwX+BWbf9EVHSskNIf6/m9Equst4SHW4lw+4APWGz/yf
nDvyJgd/JzbVNX01WMEC7cekfp0943EIQ4ipzTluqA7teRbBO618R5eXf1Sbp1h3rkCZ0SAvPhSX
SNftwU3x5k51QPgpRaC0niA4H1hba0qy/EHQnduMiJYQCcy24Et13TjBhPYV5i2GgLAAVlnQ0Q87
NTevkPM7BD7O9gGUCUV8Iz8T7XCm2XEnoCvhurmMSjv9vZaUiIyq3zkvSVG5+RGkynNcOI9AloZD
rneKXswYi0b+cHUrXk7oM0BCGOQq2tEFCtQ6JnCDlE7V7cfZDs9uvxsb69zpHYWVdCtNX/Jvmowi
l1XWQyEQR82w5F8CO62UMFUxR7YpKDz17HE8aVM3y5QPowNO76kyvJxJlGy+bd2vBFRH6636UtFJ
QA4wKMvE+aHy4tb74dtHAwga6WlIJuzd37O4x6j3j37Wk4JQ552HQGtP9hZUuLq2CGpMWXAWDQiD
LWGyohN7C/dIUJNGggRe0Q3NzQlG5SEDNmVmAPgBl7c/be03hPinXJuiHWoy13h2q3GkuDswP6k0
rj5v3qAkUfaUnOs8a4sm/7k/B1It1NQtjIwjrBWSjn0XXj7Cw6H521BmJz72YMyEl9j2XTDFArJ6
layys5jQ09Rw9pmvoI6slmmZ9pmcCsPCuIu9V3ixhLADhAzRoIUVLZpmVL4IiXUtmeFmQCnP+Wah
OoEkeeq0mJpSBund3Klr61VY0jEk7Y6UKgj9XvnKnj87PtQrtac/5BHmE78U2qfQIkFYNSkOR1JZ
uxcOyzfacc+LQyfptTqdRYwbuQxmCkZCPEhVn1Nv/24PwQF9ShhkaHMVf3VlNR++UUI0HJWGmuEx
S/lP8td8+IAjWg32HZKqgWtG3oN/xp9oR9IGtWz0GFUQTPFLRKAd7QC2uldYpvmctzoOet8VI0hY
xvt9dCvmTAWIy55Qe3FsWn5iXhWNjclOFL+eAf6H3GjlmFeXbemdwCWNy5DOiQ31YqalNW5IJSZz
shr0tit4wyW3/5RO1s/4ew5/21cSWlEnb402BjcRF3PQJZ4f4NQQrc09Ba1RQnYfNRrKsLLLm+bK
AiwVBtgI4oA3mo0M2WXnTtJGqVlEBnRnvISyhzW0lOXnT8EYvcnV+pT3wIAQH/V0Op/On0cMz2Gb
uduW49JjC9feWyxVSdlOqrm0PR1t/UdIhrOD6G50UI43kklPOaz3Q52Yg5ltLbpOhQNxazeyFV0u
qH5t08UzCckjZIfWPJSYcV6tgTYYvII7cN+ntJD1Y2g09tDpnRbPvX6m7/iBwI9uNHZHDfH5tP/L
y/xI594fOh7VfCq3YzUxd2YZSNYMUes6H3Yq6soyTnZ2H40/B1iwXZ6AmhtUnAjhvtQt1zEh3dLR
5fGD2uqEwMdbGJZxWTHr3GjkAjujbl1XyXpPbRIeRlajPi0rHmH2p3TbxJiJYFmgE77PlljzWY+4
zJoin+CNCKtOIvErC9K4KU9g/ZP5O0XUA41KMeiD+9cSV1RgrMe2ccmbBrGKmCbGlz+znBCEjbaE
81a5FgPWZqK2a2edPE4eB1r7YDAxHDOIl3KTJgj6tb0M20vxbjEVUfNUABzECW6Cbp/ruSnZPjTt
MKCROOBeThYRm4kisnqsNW9crqpZ9BrJgljKfYfAyhlhylWjgaIywPo5Lc3jJf0URL5jzlh3/m7U
Xruj4iSxTdY7muoXJy3IDXvMunHkk9mtuhTOBTeACOlL3EFy9ZfQaplBQfpRTNJ8o+4ewHH7SMdr
AOh9BhGWmWbOtRQCVkIKKk4se+Apu6OT9KZe1K0uY3nYXc3CAhLx5tNK6q9Yk4wcN7+2ka32b+an
OzQSkUwkDG/jb2EmN/EVz2Cca0ozUa48Mhi3pjw3QiO5+Dt7056gZt900RZITBM+83Ui40Hfdqxv
R/eIxP+TZKN21GLWMWLJIDdIgfnNCmyEMvJuvURIS4wpiE//uPjLQy8KB5GiX4wjv2LQXfvZLhiy
qVHOKUb0c2QtaCkasmbRD7GiuRAr9aVn/udw8I0yjNEO5QlotA3Rpkd+Gt91W9jdwCgske0zRgq6
cK5eDydp2Lo7FOtMXB/Grm0nVDiJ5BlLxABb7Bl79PkEJST9B9/juzGHhiIwZziBAunM2yIaz7oR
vms6RyDgqWvwiV52a9gQyoJtLkE1NGAIOHrPyl5yxrFMuJbQGqliEkW9Ctc82U78aMVE23OsoauA
dLuBTioNTGn+M3JGRrt2k/C22xpNN4BHXD/ExFoepqcdhLUJQN5UtcJvw3Sdhijw3YSohireKJj+
C7S7QaJdmwU4MrKd9qIr9G4Lsq8nBNxjOXOfc8NruJMriPWm/dsyC4i3goLPYptOKP0Vo93IWjwJ
4p/At4uJbgF/8L3Uep2JEFa7IW0MQzeTfLtHV9Xq2RnS64lF+hy/Mfzt9fNn36fcqe+PWyS7NkS1
zq2ctOJS1tWNK39coGXVTwHC8LM5s5VM0Fl057JFT9jDnTRYACii4fe6Ek46LbAElr5pecJ7HNqE
bs413kxbBbSzRermPhKKgRZkul5JkMMGCW7IdFPPCqpzJJowK5RhMDaWkZBZKjZFnsx//pxUTwqY
xByqBheuEd4bhaEBKGxzOQvUiy5PlI/SxDAwqA0RBx2dOWWoKN5L8YaSi1sb1FJ0JxWFMysysb/p
2AxLfQ/CVaMI6TppMsjK7X3KM1yj3yGNljhdbm+aYU6vck8O77SXHoDob3GC9hYXsHjyqgwN9+F+
UzaXP0tVBKwLXtqDlfiTif6PeLFX3vMQB42t0xElyraOb2LcsGuFzkB0KA2XK+eN9t4OdGx1UgR0
R+tcyNP3NUrNVe5q1Z8L8gjvW6QNU9xK9IWM+QpCuiOYK7hIR8JS6QMEqrCY0dINl8YEAyuUZbu0
yyP0bjclL/tvKKjh1pjh3hTP9pUKTm/Q5YGewJql3kGePRGv6/MMf5SUE5p8h6robOmB0dMnCbte
v4BEu3yrHhl1nVhQFzG9eyzR/6w3ypdd3oR81ILx35yGz91eqjMmYDh+UuSODm+VLIkS0E974RYJ
hF9n9teQmvwJWq9yOEnFCOirV8QmaobeOANZs3vbcWaKDBJV08LeX6k2dyfkSo9rWTtHtpCg53fZ
B+GimyySbrxvGukTA6UoSjlolBzT8CuOr/KvW0GSaRCQhuK6FXg7FyPttrBmD2x3UHYwzo4eweg2
czAoXUUbKrxn8J/LmdLfWSvX3Fw2MV3n2ITHbqqXCyGodc0oSNjUmlCeFWyLPVZLuymV45jn8eDn
LY18/JXpiPpXqy9r7hywVoknx04gq/DuZLc20vJibzPmoj8e7q5nlsU77fFfQvkZNXoAedSFK1/i
nvan1Gz0QCCXS1c/h0Cdb6BHKf9NfOvUQab3vuJsIgCB6xGHjii6BLRYDfMwQgaw5SSS0kHO8hNs
kI7qEuhnD0Y0gxYz5fddV608dgGpjV5rCFbpIVH7y/bRspzmaHQ10tXOgx/gHTt+/xnk6drHHDc1
jtGf7zCkUx27jzZwnSQsAyEJgoM4FGExoKiWg+tvjNSYXd2xWiEl2dkEV7+oYR/4Zdfvs9SHlReX
DWrViogodmULTtcFpwlrL0jO1eBMpjQwfLFBbtFbEHT4KyTq3tM9/0jE9/8I2GUiJXiZQBXHOOKK
0MIldcIRFnJUGuY/S77XPPrK/Xekeog3325aLLsH/K7G8GqfA8aYnao5WH/wDn7h1D8ZxIaOVy6Y
KvWQw4zcXUvs+R0GnRmpjRznXRDriil7N8IioEBd/aPqMIMpYuuLbUJmSMznKBtFD4sLKpdlwYTn
UN2DGI+fzSc1iMba18ItLzU4O1WEj6zzN01ThbPlWBITUmRhFAcrjHkvGi6bOc8b46Cpu3YO9hgZ
YoK1KGIITAl2TLKLwIYkYmBoTtu+0aaOP80GOnTmd0wEIEz5AKfTsEq0CyyXO3R3Oo5M+3mcvjkY
FINXlHuy4nbnrT8WVDW1foAPLP7B6n9wnKnXfgX0pcn6J5zMUyR1ANQFKARFyOqamNwV216awWTI
pkG2LIGIvQqEsNVOYYugRtykYwZQWvIdYOVCXco4xY/HDzeohVxwfrqltau7dNdaPjgrHtVIRyNh
1MftuQ2mW4C+PKVnW3Hmvem3O8cS0lycyax3TTm89u0P3jKQ4cy1tg6Gu4XytwQy5JrDbgR7MD5h
XSRGxfu0yZr+ysGaQ3GStrqA64Dky+UH3Gjy2KgqL5RgHzDtHBAriel2rw5tSwk+VmacfuNU1xUt
aedD4Z3T+VFjV0SazP/DDOASPc9loEWZYu3a89Fu/3tNkvlqCzITjVYKKlhVvSNP76Ey2X1sc4Rc
SGdnEKKQaq4EwZmIH/mbuEo5zu4CGt1q0mWzs7PIyiAjsjGnWRythaqdTNnmTiRVwhI90xb/Hgyl
/5CeukWpKty5Ez916mCDd7FMTmXMYxRqSGqFEzNmj+Cn777BFThL+YYKxE4TvdV3FqtfV5xY/mNO
Iw22v5ra4P0w8SyYOYopDWszlfFctLyS4MrOWfQ8nNefpWWnn15VrTPl6/7ieJHNSVPmtOfEKk9n
TsWWOBrFYRhM7iLbQNCChOykAYNnagjX2OaV0FWo0w6LSyqtM1ovZgJH6GgclIWxSumT3oLloqLU
XjffxUlUEFGgEz1TU2iE2alR0taDNyezzME9gmH5iiBELkmkpmMq1QicZNlxGt4FxFiJb8fYc0aC
aTFQWIMn7FNDDDiiYU36pRv8ueKH5h5pKSy6ALJBt3pVxCI/rBptXLJcgkvZGspUz7U2PsKDPEPv
/RUG7uEWeGBdD0BqiuCYrSFok6j2F0Zb+5uRkxpuAONp4vl1oLR4oykIJQM/CRFfptYKU0jlqJgA
sxGUnRgrtG7AMEkW20oFxV8cjTL4+nWgGuqlSPoNipWV1Rn+bKMWoRgF6iWipiG5DL538LX8YRwv
nABpPu/+aJqJPWvIQMOqZolf7qf2WglAocj5ab07/qqKCYW5oSZ7T79ibER9aYNJA9wcA189MA+f
dH2GdDDqoHNX4t7kSkbDqHbTk1f+21NbtFzdILjTm4yKEULz+FVTXzAFV3Snjl9hcNfBfti7zB4F
J9Qi0pFqiz6oliF1BMGT0D80DN0WyupvloLgU8LiwoFoG1xDakD6zqaludIVT9EnnAVvndx27KgJ
VE6V2E7CFLxoOLoRcdpSx3vM3ssAslf3qFGLgtLld6uKr0bjr/rTAptTMub6Z/jpYkwVOor1haIc
nk6/5k+UL/OWreUqb63nSQ4lgmkjFn8iOt5KSApiNj0GUG5Up8q5DK/ANOrxvIT5AlEsQRDPMSmZ
YyvNL1Dizd3l9Ztlnm8SMsMDDxEhngH/Krfp4rzRjB7vcF7aESgtjP+8Qj1SJ52AiohnvvxsLNXa
7h2fbF3csVp93UjL5Hszi9VmKxsIvUAMliF6gZTvhrwK9h2hhbuZynEZF2RE23ecrnw/MzEJhw9H
82o205cKHMBYdgET3fNQgJ4cAkKW7lFv+G+ZWXUOfQEG7y9/2i4OXYTEVzQ0dITodduYggWmPDzt
0jR8Hst8/OAc1Z2f9mmQ7K5UxyZ+cm3i+0PsAhX7gy/dMYhANmtmeo+UiVyjSt3FVkRfyZK+3crr
X4GqWvdvr2hyJDCgBiqzhI4wZSvBW+AfLnKRsZ38myma+VfXXPQawaXuiCUtYIPWaBHtfgvCBDFX
DWh8yQRr/BLX2VkfWGEO4xOuUfkdK02ftYOrTiSJ8GxPybuVnPEufIOt7/p1XzIFB+0tE6w9cTjy
3I6cd8/kkCxNJLr1Dk/+YuErVuAAG+sx4B+vgOCgBpKLuFiiVwauficiXOO94dkVcce/VqMT6FjY
BxD2Styn3Q4Y62XAfQ1eJscp0gbsNUzHD2e8ygzXwflDPmwVLK7AWa0zv2YUm5iHRMmzE88XMdEe
8+oGLByN3enmRTit0F+6F9xnz1I99S3ivxmdy2TfpSSNWYK3G7VGFMytVqT6qQ26iAlnJUyx+DO8
uCkXu8vbOcp9gcPbsqdBLfGHK5S7p269FbIOzh59CJXyeja7WCQRHGvy4tdxkr19YyzN3ZdiMs1l
0QFAJLqMkLReb0KqLFA3PyC3S7H7CtCOlq0L3f1oQ+tu3CBQgFXjTVUIZ3redS/Oq90haslmYufr
+r1Ng2UptUd5Z4DdEjYnVgCslvLXC81KcxRwJyWg3knF9OwILAxnL3NEy95EYTyQaipk+ttEmdRa
C92dyPXqT4Q50oxh2/gdxiRllvL/+9wxo9sGiS0ntzX/h+SrteadQuUNdsvXuHqjooPso+SlYzi+
PfoD4CPHaoGdeTRjZRXP8LI451o+qIOnNZgC41ksEFHXOvV/Xeojd32ocF8wTZsBlAXrTqTg6wtP
t9uW9brHtBuUvm+lXK0+8wb6+Y5gOJDG3qd4y2J1Y0no7hZvvQKJopD3AN5DFB8wmCMj8YZbioev
frCoqzY6PCNOwJ6UA5Jf/RlDcM8iQa4mnqCubZ+Qxbd5Z74tr+ig/da5urnRy8K9AQw5bYUNS2/n
iIXOab2Kvck0sGB/TfWdscTFIEMAzSqDp+ZnXDHHrmtwk2YaHvbzyJucZqhfXnt1WYduYzU+/fo9
HUSeTllzNE69WTe6Ae2yVQ9Gd3y/W8VwrNgJbfsJe1pgESo9i7nkNP4z0Iz2EYsJkGlBapmYWLxz
xIFMUQVqmoOXHwuxQiZ0bdL7OZn4//32qUftI5NTnErXixMbdLuJGn7K1U56NDsdkNQithEZDQsd
zVN30J2h/b78xr8P9P4ETWHSvdIlyO1hqBXCS26M8ITiCqO3F4upLiNkfUVDxS6uTJL4X5ZUeX9C
506TYcJXEr6BEzYgg40g6kSLMHK/phUrqVc2gI79Bq79FSBRxxsEpvoisoCZjA/CLmWkXCmvkGtN
ADEFm9y0yDWjY30bwAE5p1eftJQv/v906HvSLvZpML6WxsIAwbwcAjH7c4VQvtNg92TkMK6H874a
vRKgncXjtmvQUkceayMqFj5SUR5beoM4UxRRGPvAKvLqzYGdRwIDJx4a5+aJFNNDfnUtbkii2c/c
pew2kw375paPDCClWIQOvuo4pyzVNbAjYacECkBbeuYUE238m94UMbTWgWyAz6XPiN9klcijrxLc
uwxuyBUJoFG4z0bPgM6rvc4TmUkCrAaXtC8FC9RZD7NhXiuUcHbaKBiiZfGctbx/COmjlIelm7Nt
FZljExo9dp1AB4rRbsO57ygwhfvsRg+GOherrPf4NM8RaDXsTM2Y0YpQnuU+X71C6IAn2K9Hjp3w
0BH22lWqE81Ok+J43Jc3AKiaU2MpGcuu73IXSi1TI59r0CGF+RCv5UylgcoohXzIti7dL8lX06rn
1W/F2lBs0kTluEtxF1SogjhgLP8cB7IpIqvPYSl2oc4QNGSkeUZs9YJqNCOfRLl01CEcAHpuiU8O
XPM4K406TsGG/nkRvQfMa0kg8qm8503BiS0qPV+V+QgeOPtOyvbZz6lL39GuIjnZ8DDiNv2iGkJ5
YSpug2fUjDOFcmubFUmOxBMqtW9obiqtTQxlYsOwkxSArGw1fwQ1DDh/TpLGHC1OByyG/je+qPrk
SRcd4/XFK51DFYEE2F7PArdjhTmLq0XjjYW6KeaE+9Zgl0PSuuv+eAkn4HQYSNeiODIIbfZ8cz6Q
/weg6kUCnmp2MKQhESkzR5/6Eqz6qekOSDRHWq79QwhZU2TdEVSS33CzkYXvdmoUea0JBnZ5h//B
tICqF5ALictidF7MtoMKrNEFd+2y2ONWqAlL7iw626fPMCJEOOKvgXzVoJlflXX+Iv7a4wGPhIfS
uS9YhoqWpEUUPVovOAsoBhTxUUPJ2FSn83aJs/rldu6qmAXaHa1BAuGdLZt5xIGSQjm7HVyqhSVb
/gMVLzqGgsn6Afc0qNILeqxiE+Ahpzv2c9Q0z3lG+vQnB/KTZOBLXve+Y/HEOADCnGUqdf2XtFG+
NbmiccOgfzH+7ABaxpGscrsqNJf6FHWu/yAS9dhZkUMXOxoB0HgNnoRZlSnOTPmqiztaUZymtzbc
sFH0qBLgdwok+2rBRPn5DR9PvRItcTXWaHhBvgF6UAxUbRG9pigU8GnJFrzZGpI5Ktif03+wg/+y
K6Rn1A71qDWSE50U2A4aAO63xnPnCuBsrTYZic2NziAAbeuh8sUW2PbAyFuJ8n/ABQCSLPglMa3a
XQyjVqZeDYlBELjN5zNdXTDxxFfZ0sAtt8DUfTn9qZEyOLykcf0iQAAe8xJYCIQoSs4s3yglD7Xk
u3gaqnJ077mTGXLd9tix2Q01Snnb3Cll6imFwmnD6T11ET+MyEBw9MzggjidivjiwIZJ6LJAGjVI
nqGPSW/ChkiAnKxEFsXlEfzKgyAKWhrTY6OmsKLj5GWneRblc7tDnxh0tzZ0s9JQsdjnVkAUa2XX
xFmNe69ngrNTVrXsxqI0bXhE/9efLXmiFpWWizZnURwkNXP/E04ZlYLDrL56Il98tdY7W1/ZxyuI
KCMCTHjr0YLMkDS+NAfFfq2rEg+ikhbMQyzrGi0ThmuctuyGmAZngPdcvS704PPesaVnMIW+JFv3
oUOHdz/FRgtAepIQW4WvMAiBsfm1nmmD7yeykQHWgF9JX1GcmeXFWTdOtYed8ljThhdGWOUWMbTb
CwR+WGMr+StS3Mx/VK9dnqrSMf4akTYneM5Yw8af7/dLHwAZOxXq6oL2jZtKUskayaH0hB1o1BWQ
T3ZmdH/0ABlGz2dMTxhJZBpxpQ+pZhcu7eCZaGupEWf0zkCFnfDpvyHEHkpt0KRJjQqrcLY1Z05p
9HkOezSRd7N+kse31SGPZLxAEHxgXDs7qMxlAoH1+QR7kQf6R6N3MwO6roZuvdc6but1VJQ9oiGJ
DGT18IgpSdcykmpqN6qzCmjFRa7HoNICD/D/wdoqo+5ODy4EJmcfQ+GAw7VLLdjhMLWlH1GVUc4S
G+TWzcSncig+1Yo2BTa5pI1scKbhcKjv3D4OtqsXeWYNHKenGEgawP/Y2oNmAW9fvwPXrxC/g5uy
Ks8E5onWUrvSmnfX40Q0hEA4rM0mHLW2MaasId4NtsD1cmL8d4Xsp8tupwZcuS5Kciun9ZnK2Nek
i/wXoJrbxlHsJF30Y7M0Lnik4QplrVE0qkfJxzaKqfQV8HpNA3CLERoTPuPqO6nBu5la9dTapIpU
32Wgta+uwP8U/+RqRMJE3DpUMVIwunvyvqAc6yMhpplPBXu3M4cpC0tEYL4s7i4BSSzdsH6gXsce
NILUset4IpUfBZ8YwLqNjD335ZUIn/75Z2JvoG7AHrYc4v0psKtSsWBvo74Zi2Ma3t4qHlbsheNg
vD2wAT6A1/DAQUi8hU/En8Cgo8Svzsly9OZ9mdEpb/mX8RgeSt/q28U6eKriUGk5vlv72y7X72Ue
WmI21nWz8QRx8XLxCUBBz6QiJex4ZsnyPyH90Lh2LDjB6NN40+Mcejy03QE+ALlF1l6KKzmFSz3a
WoXlvHsbKprScJCvMaGT09TR5A/gc7ojFC7N2/OUuczRvKU32jVCYUPre+o7MfsF3A7XJ5R0ovaO
vhqxkD9FEtWyuBMdeJ9qF1SMJBsSzXwLm3sIGKsy6YzlC0NKUvQZWQDtN9uLHaApq97bzX7eGk7X
WO4OvxsJTV+pCpK4htptDXYSl6byS7OlhCB4zjzYC/iJlb2mWk6SczoYF/9OGmPJAwA6eV15meka
Y/eUUV7YA7lGaCFJ+1iPmD8V1c5Xp0Ldu0vgDdieV1vTLOyu6INXOxuJAoZ7R45kEoSRt7gR/Y5r
mT/BY7hYaA5t5HjqsHO4QX82ZI3CS91gr2/qk/YQQxhSAOQOTKHl2xBLKvL9z2SYvUxf099MCCPc
KwLPC3ASLw2c0ceR8HuE64FFVyRHpAWVgeDy3dRlfGP8gJr4vAaaB0y7mgekKz6I9LkFEUmwyUBw
bmG+chX4wiyBKPL9jK4/GtWFLL+/BBeYAc5wW4IMn/AcLCjKn+UP1MesbRQBUzeodLruVKXZSFZb
DyaMk12ZNePgcL/DWfcdyctF/amDdE+9w6xdhY9qWOwwW/YN8OULVWcQaNX/ES1Dk7d9UUWU1Dbs
vN1Ov7WapkBwiYv+TWsHTRPEmmuuylrJ+09rBDXtn63kIK5Hv3OXC+3MYa5rkUe4BlkXLXTxD7cw
ghHrQ1YTHI/HMo6yMoNKumI93l3kGYi5ehEnDOZ4PkKbRMfZx0CG6nU8zdW/FM1KqpDxnH0aBCFC
Zu1+X+HZm1qgg1arg70CQFlb6bDRF9e/Hlm+C2BEU134fwm3zZLQLzQxR4Yjo1VX9IX0GiLwdNys
nQxpVJccZADlKU1hI7tklYhWSGHzjsSP3WqPCvSqkQQJ6Ks0jTWrwC1qcvbfer/rAR7bSZ1IB0nJ
VpVABvda6H+dC3Y80Q8hsRDmEHT8yB5cSNiJVn/X6ure17RINsPfmrw4FmmIpMO0FxHUZfG9IpLt
dPU3SDJm/7ws/7H9R6fyEuibZ44M3RgGVTvMh0RgabNTMfNTXt+ADOpqLqrAXH8Y/R6qEtkKk3o7
YaraiHEJLxQ2ndY4v/dstJFpsWkDErzFh0gF3Orw2pwhOirBmEnk35SRxKPYXjIz/pCE2bUhe1vp
uV7lyoXJA7KcOiGfaC4uleJhFgL5UkeeN6vpiN34jE8LGIMWuMFU0KXBWhtzGLtYYBDg4agr+4Wa
U6Rdq2vamPb06cox+HWCET7DTGzyXYhV99NJtM3kb1Kug/3nrpdETZ6Y+bRvq4ynEotA5tmSmZCM
ON19jWpsQZs45mHmv9vuTeAF6dR7rP3JQcgQROa5O0bw2iK28pzQdJC8NzoUV7uLdgq+xnYIt9oI
NMcgiGo9ZgjkBzmE0EhpuebZ3RLgbdkYcFjksvgiDCEfOJUk7Uho86F8iHLZu6W7RKhKhlJRwWLj
a3AqcyuDt+IF2pKu9BfF/Z6Ny1t+2RqWC0iiOQhlK61lBXTVXPTt3fR6yCTr1N9IOSd8QyHc3TM/
kRAEoBJiBWXfVztpZNljgpBxRjBHsRIurkwsbpVXOP/bZ+/91mT6tpCEP1AeZlBbqHIZ1lFbvWQJ
BfJ4Sq2RbcpCkUu8VlNNUxnRiejohL7ZG85lELkc0dTu7NX4+lE4mY83RAKO93ILFYLpSFKA8EZG
YAPX72Rvbo8/EZM8tdY4r5OJc7Qx82SW2uZJgAHzSE9XKeiq98937gtwIDUAnF5qXvu03YyIbjew
CxkMg+KMqyfesQk4axRKrhDGbP9KYTVAu4Va1NZNgSSlddEBNukx8+/6PXhIMrj0tbKadbcntrpl
+vRx0NgDSJclzX4YjWC7CEJiCImOgK7mCR+3L2a7eZlIUhefNC/ULisrri8vARgnkqU6lKrASJAV
Owckl3K5ygabaNHtTXA2l2mpR21S8yt5wxtZfNesMIxHfJAk1XBKGi6OaDVAYfLfymnKjsQsqupb
XSpRlOhhOgk0fFoBA0bx5nTCElKbb+QWdRkGcEUUz949tYWHpeNNay11EQJiupXtSqJvDC4Xr0kB
Scw6/eYq4yDUWup9faN/KmMrcAmP/hUfXRZvBKj5rNzrAurMCtJ62RxXZn7lvKeXU3QcqjI+obYS
IGDp4qI3ZTIyOAkspn/B/4qJGDAHoFo5hBK/4nNKsF+jV1EFFtec3wcPn+86ZQOLefpP/CKnsXb/
PmS03PzwXf5VhdqzLJEokcw2pzk37t9oQo0iMKv9ITqC7j12HOV5dixLBK0IKlhJ2taxOU6nDSgb
b1uQRFimuWCKi3BbGLy/+q3bYe3UBbfKUNwJE8Nifcvrra0+3o4bpDFOsy3uJgWn251UMQOpPFRY
177h3JNiWzvxSdaO52/PxqTCPz5zFhNuxneMe7snw9x7p+9xK8ooA1Q5c0alVA1MZBOYOrIw+eik
2OKGFsbaq2M7hZ654ShdFOlwk72+eSNqrjJx/lx83jhUXYpRcNILTXDNcCHwt/s/yTl5bxM59rSA
cLdEcB6dmYlB+TZ4cSyztdTM9GV0M+BYv+p0OABy+v8uYxl/88KW8hsGDRHVV88+LeApo8d1ZJCc
oL1NjwD6ph8ehP6YhmJwef26EHcmJ2GfZxX6rBfeakfKWLwQ6TzezfJFvt6T/9w0ojVKQZIc8+4D
DsncP4Qzbuynb9jg9i5r7zkoSpChuCl3HvRVklc87c65a0Y0zJ30+dSMs5QCd1y9rIAhq856hswZ
zcXbFrXP7I3hgFAtCisq1AQ2eFgqj4bE6qxANvy70U87GlJQCE1H4BytPCHeNdVJltn3ozXfxbNw
5Dwj3mqWov/PEaAhnZEq6zfqNTW8FvWAeggyIED1cKye0YU/S3Q3HAdmKHZJOKuAXaJh4Bajdx6F
Jum5TRD4y04D3khJdjQf3NjFDcupj+Fzek+6ZLuAodFW1sRdf6bC0S+78tdnG6KZbr9AVhfNgRn3
wwqENZAZ6zT8z2Rv/E2aV++1NtOhFp6/umUhk8TX5noOH2zP9mdd2hU3kVRBx+CrVZAxYh5HjXeC
8WQcBl20sFhOf2L28yaQcmEEoF1EXNyc8vNDpPCNVbQPXxvETxx5YAch+9QD2XaM4yX1vCfQYCFX
cFnRHiNS4Gj/YJGnHBTpUjBfKfLTsC83jOszn7Hti87iU3835Qfp6uyQH+KqWyYzJjF0xZIK9YFL
s+V/aDXq8Nv/F8MDWRcqN4T8BSQ8cNajM6WeXif889wa8FQum3yCYLRhi7eLO0urDm3G/ud53YPw
rIkI0wmZf96HTzc+ORoCBl7Ms/xZlu2pvxi6wKndA8h+Dxjua9uVQlHvzdFm8nLTsCcKdYrB9L5Z
qw9wDrQzflJTkdaVtSu+PC9sEqa5K2uGg04xD1IlSoMj6VoC3Cs+SSH7c7ZQYOyjERbrfLKQchjJ
OQxkFlyp05TTDicGjwTwsofhYPODDfy8yI+vgUug2tdahUsXRZ7eXa638IUgFOVzDvwwMyGciXJm
oH/s4vyHhBTr2gxKCArUL8CnVDYtSQQrm7IXoOiuX12OkX4lcYCnYPuYU+bmXlCT+zhDsztzEPUH
SKbV0PWWmfMv8vwY+23WLEn52GdPUcfBGc2baBdZkRIrH+ri4cG3kuex1gFcXGZGgLzzaBhRLywF
boWmTAkH8rooB2jNNPYYj1GVeiZEyJcZwsBGGpBTP0nOlkB57KU26SWNwD7RkkfbqxvODoir4qCE
j9Ulxsqd9nP/0E9odxS1w2XMSZCmISpspycFCG0wSgfsmxkL2i189MvUzNKWjCV5gIYJHjF33Qw0
H9tE6ur/Pz7G2m+VN/koQOs00B+Co47pYwbeU7VdhKUBpZWvDoh0o4H4i4nTvvlSljeuhPp6jf8o
rNXLbDRH8a01cZSeph+PQJVbD34oZGj8/fxWtz7KggXfUmmsGG86ufsUwyHLefA366/3JCkAKdsa
d5jTTHCHS+1k9f9EGBcOF+iUiIxSXXl4tvru9AAejUBHkt5Uamdl2ZE7Km6P+AyjFerKrmgmRbWD
S3nxQ/g5yxmml8HLkZrhV9ppxyb6SHbO0Ho8GoNDBWyNGnV5B8xmm2gmS1uyxOgEs+IpPYc6EdZ7
wGFa/608c91XcP/aSvy+qQd7exVSc490FqEuOjdfyXwk7Q6iEGAksxPypOgIe2W91anrqO9q7CPe
5pWz7jStK/UbLwj1JuNi+JVDQYxc4VWJRS5SVqeLmVgQ/U0euOjKThIBtH12rjirjMB9pkPo/x1j
lfUyA7UzTpGAovQzQ0HR5/R7GlveSEubLyHHf142ADde2HM2B6RCqyPUW2YsBCtVJnE0vuAa9vpq
/qbd0vw1tnL1bm3szxB26VWU8S23+J2Mr2CO1z6aQogmsMpMC4QL+QNEFroNNDc4+pzZ+TBVpod7
rr45FuDZbY/R41EhCr+C/z3FByyNWtXFB5ncE0bDDBMrujfLkBwi1/yjvgFZJYQJlSytY83gdBng
Kx0VxidkA3FUlLxKBtpatvoyAisEgaP4/NKw1XandPQZmGMx6/jHriP6r6DLhsaCaI5OeA/CZT6z
L/CKKfW6XSJ3jYSbLk7Z1+UMRMlgXgUCN6hywKDF3SKR5NJbll71dc8a+kSV11A6Oai0C2b9qyVj
QuJzI9SlTRP7rbCQo1Q3QrwLdIOWS+PyDZQDw76gDs5J9D4qAw1UGhc7s6Tk8M+9IZ6pHGE3K9ND
8JFvB2lEKwCz7dPboUfv+ZWRQcbytiEuEsYV63YhUv1VgySgqfx+vMxxL3HwXa/ExjXy7Vb8MhqA
QS0fSfnId8UwfJiaZ4NcAtnbFpr73MalFmsPc2Dix34enyuB+j97lKHoNXCThd0/m/+GPm4hisZC
d2nJ4RNBosgNcC2t24PT62AcwHVDCR7jocYXlZTloM+G2iB7Squ3RvvG5emfSO5vQQ38LmZe4RT/
9n9zzURO2Fslo2ZPM6ks8tIPyd4g/Ipo/jfGMSgdeqULF56o+GgtnPctPTODyjuIaAGGsfDqZlGi
pvRUmwD8fiiSrRGomhyS6vjrMuO6+GU5bl/d7YqKospSWVSs5EXW1Mg34er36+/8SamhrnRSZv9W
HrasIO51tz42zImRJlUjaVV8PADfeXWpchC9TT84THDmd63xhQcH2ekMkm/ffuWQmlFlnx6w30wn
wRGfyTT7iIPQTw5tXDaGd08v0FbgPhCjyapYHqRiorf5apQmdb+7djaRWyu3vv0gOP2/62lz3ChS
twjES/iy3qATYwQ/6TLTN2KhdUKYRI0vJfNfPpAze/pYW9B1sLKan9IGOLPddIJ8gy7fbdcnAFAc
ARNLCGGZAQq+QN3Xpi/uFqafAn10foRO1Ag+7Z8Z2AMqCyeFfgkELYXVzlQW4Cbq38ubULMw6xYy
JF/fwlXO6nLsi5l7YUxfOGZJLcM0TUYqtTSUfO6REnwn965wtGd6loBY2h0ecX/lZ3e4qa7MrWPh
iTf7aG75EQVZ+cCMYo2RufTIcGVBN9rW8A5LRgE4SV/O7Kr7nUuA9hGjvdWoPxD7LKl5+1zsuuzy
LuARWQexqbbDxnWIVZs0LyVaDzyvvMa7bXQOZDs28zap8f5U+K7tp9R9IN2GTHinyV/+egXGpZVL
67sTAvMdITevUheoF9WivpwGOa7vAkVM1XKz6Y/WIHggTxX7fd0AscxukXI3aTJtrEEfNHvqhpch
uh9DnFRAYiSsxxU8qobSMg6s279/nJqBhN8Odn7DT1neiZqG9JB3FAubaueXmshz3uKPGYozXri5
opb9PIVkC+CFStXsMpRhVqUKYX1ggo2hR+DFVSQ0KqBCc0+ycweu91nNq5VJ/mzp63VmXJ8X1S4P
9RN8XI8zZkWdEUluhXo5A1ZpCnsEyiki51dC1uT9KRORuGfNhTpj7UJQrJa43N3gmVr61Fyv4crK
PVeAVOxFwl9H+YS3+rKs7hqbputvyCOwL9/mW3Ika6dcLkKRAviGfVSFd4ih6o8Xpu17KsAVpwDi
2PTtY5xnsmkQdhraj+JXtZUz/xP+hkcxM+UWeonjLPk5PUrWqd70W8zbdLvumblW5vfJjoJFKK8E
OS7tKhEbpgs7C5nHDYdKL4Ql8vGPoN92P5JI8i0Oow9n3DgNY3SBkmJpbWOE/j/x4ZQCZLZsDLia
7Pt/wmo/k1NKDqcBRUahhtkqO6r87c+hvEVWIcKsikEdddYlDrweJs5p6Cp0i+vw9wZlMuMS8JrJ
RyrPIbW9TIpmaaIgm6avz7dCIPwzdpHNUiTMhoObpiRduH148yAGPlcf5vnT8wR1O3aBxz/pLdsu
E1DW+4c+mCuHZAzld513ythufqg7KP2qoel4EcrxvfQYtc8lr0McbqRbcPgZsZWj2nahpM6bVDpu
x1k72V4Z7iNBbRLCUfNqd+5q2x6T+L72fmF/eMUG6Vdj0C5ASGk9FIo7K35t4EYLEXzUZtjx51Gw
VnZd795yMN0vSfQKu3c+h2Am7nvpyrXxhDQEeFHxux2m9qHIeukkaOnIwBM6JqAs+0bG1SxEaQXg
2/K7SuJxSa0jgHMh4gvesGmRCFCKfQDE8FeuxXrmW3TIRa5zcPbYtwc2JWMdNsWhn4LqIhJPFRAz
4cyDaBwgcIbmhzLW9dS64yroiXyww+EN/XW3AV3G3Isn0naxcrEYyWwl+VCo0/Mi8z3N2+4q8vfm
kHM3FbQ2BGOg9YOVowrx/KKWoFWEyQ1Tir1DKBgzwupg1uv2scqyJt+at6j+kndtUNbIBfkaeKvZ
3KyEI8mvF4M4WL77KFQitVzD9Frau6trI7lp2LKE5N2oQt7L2fNwDaN8wuHjgDNC+fBY9E2FbF8H
bzY89dB8tbs93kVWvmDhAthHXvnDA8c5/B0vDa2aF6E5EknTCbV6CyYDtVV+K+hhcamqTsqb8pb7
EOVFbJLhfVpFRG05BU04wR4zL2YLF4KZQ61ruZ7D5OLyCI+klR1dSyCjXqGxWduXdvdKcFTcHNer
eufkJ2LuO3eRrmrFV0jhQcvXxJlTOYZPiSzLYOWYIfglNLuog640tcMF+wUyn1sopdLJ9vKEKTWB
0toUBQcJ1+7KxQgIM9ImRdbGQPXRO9xriHQj+kcFZC1dEBpYxMG+BBiReq9gc0XotiI0ULenepkk
7G1kcHY/94xbpbP3C3DUAe9kz/uT+KG6tixcglU4kBaTSQ4nDyf/e289cV5T7Rl82NaRe6PYeh9a
pVnt8ZmTqi5hoRqDp/nETtheI2F/CXsRw1kEdQgwAD/pfHk8Oz3/7eLKlQJY3LKr5eOhyKZqbWdS
kHGm5zwM8uZL/AOD8Y790TYpXELRDXlA+ssqa/xO2d72+U5AyWgr/fgRH7sirfyu6kjIuoEwKdH9
YnIyUNWIm4msG793TfWoSziQTsIXy/lMffY5OwKdTdYRJJk5xjS476I0J3m5Y0GXyTBJJVjnNdVQ
hiyQNNfD8wu+/5XYG8X2k9Hlk8h+UaMiT8UuQ9DIPq2Zw2+vPntP3b1ajqh8a2ls4Ms41DaX+8tD
Iq5CwPi+hFlYxjEQYpTc/HzTwzZJM1NVafHv3FkSlmAuevP7N1wU56jMYOS5GbGv9bEbLNgNU/lR
baoToC1dgf36E2gXx0vYC+8OPx7sd7l9aUwS06L8ZfoODCfumXYGdWjADP5RxzX2kMjb9c1BxTyE
gh+HKkShmlwLYExbTCIXxoO1ID4iuTSXOb/f71kgKB50S2qFqjk3DwlK9XHnNavDG+P/NNfu5ztP
s5ZBodlVUpZ4EjiSUXrIuO9ikt+IIvIkqp+1Z/LrWz2N5orWW+tNABHNvg87ozbOcn+Zzxojv4tg
tdP1bfzWvg+jeC+pO1tVJfU4vzS1rkSo27tJBr9QnTVOp8g1I5nZ+/wDwfaHeGE+81w5QjeO4hgg
51ZemawxD9sOtHBfrjL2pWyBLq7ChesK3mt0BscYvrGq+om5xxgl2NsWI5d7u/5vrF6Ai4BRVMb1
zdEobxPkOYQ/IlGY+7r4ZTApgjpy1ZZSLHdttTAqcU1Y0ZqL5X9SOkQiZkGCrqeuSOJIQUn0SD/9
syo+rSBV72jYQKo1o/bdtr8W0S1R5baQDi8QePs5oBs5NQAWqYRtOWvmnEr5NeAQ1eYuJ9xR7etr
xb14JeWnicxw6XlkIf3o2tbABGxuXDQPlb4HVKKVXylJ9UgkvmkPSkpGvAjFojKEdZDmq9vuAJdW
0UW968AdmvhB5mtz4nH4pT32if/65EjY0FrADoWdLqDFCzJWcWl+KD+B/QDM+/5XK7IMVGrbiLU6
c1Qbn/4IGm5ICufzS3zUnqXUWkTeHq+rpJlWMmMKSoEL3LQQr/ppA7rtnm9fBMIBVxD0nv2uC22B
fVDACw/n+GPCNxMnAlIoZvmy14bV2o1fJEAi8F4qLLY7K2R3p5fCWQXUkoN9F8RScY1oOnl29u4j
+JPLM8aa9uf/nFtVFNI1TIkTDDwE2OLZ2kkqtVS103vTdeqEZjvhJ8SSJjkG7ctLWkFixQ1D7mMA
b13sWIgCMWpFzNQkQw/1N6EtLOxoA0pd8ra8uco8wuAhdFK8diE8m88PbDq6c/T01515uzTW8v/d
jTApR42+8u9II94dThcpjbsGAWO/9nAgDZ/2e8DGNqqgMMYGYdSOaoDGwZIuLipVg8DUj/LyLB8q
tGEb5c2ijB7rC9aSCayU0dLNB4113kTxfl0Pnq9sleoYN9fVyKfyEA3t2+1gEeFu668Dwe/lvwpM
Q+1eBLsIOg0JtqHG0EJbqW5R6WLFwj7f3qv3NJ0FQVSXkXpm/Otsc3xKuYwf9gzO0gIIe7Cv87xr
xw355IBZmD08UbXAmnbZ7B4PGgY83b8JY2M2qdJV7XNLZq8ecx0TPAbwOPub2RVgq4F2r1RSyOXk
g/f5irrVARRjtqbslyTlXrEM2+wmJDa1DAwyjUXVaIuDkB+Jkco/MPZnI6U6npODu6bK9b6bkoyZ
BUZGMg7s9S6ckiDgwVkdBazXWCx4fcGnN/zMXavKe0FWFHwUa42uGr7C5BdlROpaNC81kuW/i2JJ
w4vSxXlUUy54Oo43KEAo3RDLE3rnP1jEc8RdzUbrnUtFtWusoa91q/Y3o9qyn429fne9VIQxuPcM
8cLmyJtD8epI6wUD7XwbPCvqFCoyf4uuiPtJ2UAt8jA2h73wnQ3DuwZSGhBDyc9LJjNAAVbs0eHo
jXR13kTyK+Gl1FNsgMJZ5EohwbMBJCDS+V615fThMeNZQjmUZ79YPygpGJe5DHUgxYsJdInHkMFX
VnSmTqVoLAhLtlUdwDFgp6z0DzDAAs0UvUqfVDTaXhIwf/6f13FsBEJCuaTE7cbuse8wz0BPxQQS
C2rb/APZL1Hum+Znkw+G3dgWcM4TonvpWeEOqy0DwR5gxF2/Jz+w3PgyPsV7+/Cdhj6mbJCPp+Bm
P+SR5qOWIjJvxga6+kpQroWkyvudWXjoW3ByVTAvyL89d6u5zLBAVEFvdmUfgU6XpKrI8Xe3nTXT
s7SfQxYRetlOOWKBcyDiBIDZaJsS7nxcsLAr7hbXjd4aU22scoJx8MGF6ZibxThSPnzoxR3HD6U9
qTazrV62Q99gR2igpRAaTOJ1VmoJ0y8bhe7Czmo1n5ZcTMllI9RjVAzGsX5KEK4xFlElyv8Nq/Rv
ra1Byqx9mAxopmr+SLfvWgQzaVncA/+L2gH9JId2UVh70Hh1F6jjsK/6Nm1cYNfPAOhn4CD21hx9
3nGZHk09iWaiSIS6L3aCzrBq9X16n1f22gS0KmK2W8H8bd7OS6enkC3jAZ4Gbo10ftqogDG7K/so
/wuHi8d+lsts0FllLS6yY1jI2Y2mHg8rfX8ZxLyyPUi5IjDJGizruZFpcOpeVFHoA6ne0zPNePsW
9j4d1bUVj7hFQmcQju6N4EVcky24MR7D4du9a37HUk4JlFjXGhFV0U4FC258M5aPsHUX81Mh89DZ
eHteocGuyBdLuWcQ7+QJa9nmZfBThhFJlO8Ucq1MawTesjZYc/9Q2uAQExCKgIc09X0o/XY7A8Rn
94mKe8r6KEIt6vg2BL+5q6IiEQx7ZTzte7MMFTCY4WKD8armgq7ic031uDUOhIRzGHwlFuD1w6HU
jRJ3NrB/bwyOlXNFZwLRcdAuWf1kua7wpC6rQcabNrJ/h7QX+dbqwL2qXlQHzUtI1qZ3uQzpy013
ZZla+CL54KpQfyzsYJxXPWX5LZGtOAsj7OyEZUlC5YiVACU2TiGkTBxrfvJQahU7LIPMmzQn/WUv
ELg9HB/rYmadtgmqv86S+DGcirm+GVzzzjsdrXyqw7+UybAdVxSe6i0aESVpl9OBluL2Sw1dBZlT
6nzfBbbJXQ82WBcgFFxWsdAuJbQpG5LyfPKcz84keS2FGNpErYdDmh8AQ/XMJECt3wAVcLNbHHgM
fse0/6EDbBuU0SxH0l4e2fHfgFANcE8wLdeWVmb6PU6csW4fee/i3TMD890Oic78rOqqUpKbJXaW
NFNW6WICFQzslPErv098at5G/7Bgn8Qe0CnBLx3g3egLfpwt5w2M1ESqd/aoA1swezq+Y2Q7py+a
pspVglkXfKVJInrB7QKXBZyhnRchQlUI6CpGiqayNiyKP6wGreyvEcTNh2BeTdFXNpzSZjJ5Asld
sN1pW1gfipAJ4zntxgH/6Y7SyzKd9GyTHe4239m+KcQXnXpuSgPhWKcBKMyVfRUBCjfwu3qIHco/
gB4bd20wk8K1sN84GNhq1/2PL2xx07hgm2ENMLMjxUA8TuEG4UXzcnHzvfS6w5ID/0JKX/DLSphL
k+erUtNwVJQfrfh1rVrWLfuXnwMEbBAf5DQPJc9hdXWT1A707MNeaxMqodd+TthJQPfqJh38Nmku
PoEkNKs7FKaxRrxDVtbwddYcBtz3lt0FqQBsqx2KpwsHfIgt3DavGOHJhtnI/AKJifWELU1glsoP
SpIjKEl+ZzlQSZhPuPpXtagGtKVZXYxMchEe5bnYh7b5gVNNKq502z6yTzw3oC3jm3Fr/0Hve4Qr
qpPNIaPxJM2NSdk4w7JERSxQfXT5j4giAbvMfKq5GMYUdycOHAOWO77bPj/ApVsRZFQ9LLoAo7pG
IDe+otD9jo89pkItWKhrj3PW6dQUiqj5Byrp5tmrtdfDq11nI10YpVzdrHqBYT1SYyXrX8W9iFiT
ONtEXZp4LmWL/WMZkkVDqOvdZKbtu7DaTpKVaiPtCzEpU4+wm+1yIUAZPPwLpWMPLbt5jVnN9OUi
RyGFO7JYPfy9h/x/emB7OpmTQtVP7QnwUP4opULqEIVfT3CI4ngFOWAPRgM3HYK4KFR8Y68vK1V3
IH4NesYlu3c/FCZ2QeifZ5LZVHgNYzzz+LTIiNqJsfaQexnZEcLnYCPin1toiQczE6PjJ0BHKLlU
u20kWQD9irHttMIRzSfyIoXoTpC5H9+XDLpdNZk/PkfzNZTXmZbiqegIvKj1WMuo51cxNlORhbX+
zCBXG+vf4LdAuUN0+Lgg/NyG57Dd6wzuln83t/csw/frPpf8Jcr+G/P1LchsLa5sGWCOa3NBuVyp
xfdf+hTAOiV6KSjqWLqYLEb3rocMgrdZ4mPni6GExbbseOGY+t9lONQJ46ISKVPJGnIukkH+47UB
UC5kc+XrFDEORBjtFOLFeU73lzMSMOwHtMnT+TmyCtp8FouK13XMKKgGPDdlPzQzXksu2D0G1wIK
N6rxqSMuTEqfsxdicvCTDpeq5zu5klftA+WSxYuUcj0g8H0HcqGrSwpllnOUN/ACQ0rQODAWKk0m
JFCXnE+pBts1FDUij58oDAcbMbp+c/mBsIkgLhZFLayFsHX+17OKTy7tkDotNbBsgL7fw5uUBcg5
HFM2N35rU+wpD1BEfnf8KbC+mc2MqPaCF66D+m1c8QMO95qBUlN5k65GFYXrq8wj8Iq5hCgpVvZT
Sf8rDm5iiLGDxYdkrbWHtOUHAeE8pWzlY9O+8hymo6gydmQ14rYISZeCtIns0sp5eYN9iIICTnTW
yArkwPeigv31EgbylJeq9Yv5PBAAidsaC8WBG2pwyy2RBdmsxmUZLMZU94yHm50YSKIPRzPdIjYh
F4cW0HNSVUs8esQfyk4B8Wa9OmupMKMlxbj+fMSFomR3Xy7W8orQQmu5c0EawHQ9PuRst70Y9jiy
wElBrv00Bqsnvgm+k0k8fYoZ1oDLHD0j2xhvG1uVijIXp8Nt12roo2doLFXVNPOTROYp3qJub4uu
8ww8DxysuSb74z1rOmPrecdeIQicyYpVOK75OgqhIWRPJoo+NVSRiYUfFpoFEB/17obXzW94sh7m
/gCzPjILLw1Y2rNQMo4eNoWpRgYF/pN/r07IC11NRJQJeiS6bXYrMM4FYMFuIMq39dv1FNMS+zvh
eQuvDoDL9fmVtgE8BbW/80qoCvMekf6oKP7FGdW4drcFk0Sn8s2m9P5p0czrBgiJx5GHETD6yvy/
Mk4bhDFour5nBsMreeTR/CzGdswPF1RrEfjPR6o+2cqfhXOTqgzm/SVI+UmUmBh0IppIL4WUyi1/
QaipN3TpgWc2kAP7DTPX0SLcfPMvziS/BdltzzXP5nFdLiQegWipIwWswywfhvUo1MF6PFj7BqaF
2+hBdGszIFZvAmF5nrIA6WiaXthbUU1clgUJ7Xf0IYWlffkrxlTRlG9kF0GEOQOlcQD92QHPQCFu
eKTs8NzDrIf/WBx4k88UQQmCyFutVS+a+WjWw6ue1RcyW8V31PW/saMpsKAQrCOaJOhXjYFgkE+O
81S+AVKakW8eOfMAU3PlDc6xgkyGz0mE8izAVzK7MHOfdcjNTIMh7uTN/4QeJimtHvJmztJ0gJWQ
aLtA9Ca3SlbLZQDgz3WuAwpyIvx9VWDnx5UMf7/42cDU/m20xpzvw2/lF6ejiNZ4CzAyrfUz7RQ8
VHdd14J4K72+PsuOBdxSLSYsjWAZfqtryuh4CuJJ24GCeIy0buMVGvPCIKFtpVwrJzw4Ak8jrOKv
cICEouzU7B7zYVM0r5tL+tPUztUxYhlbv8umA/z3AFndoS6GKJ4VT6i8zF0s0fxrORGCxCdJJwWA
EgqV496c5cDwVcyVoUEbuvB92hBoWAyAkP41jQjp64cmfMpBFvh3nbhW63fTbmm54yoyqz+iGvAS
xMoKepSEMbkTyFXOo9mPctQtnOp3OyGV+t0Lsd09FxhYUC84DWRnZkA9SyPi9x+X66/7vrbZpaZh
Hsjqr60gOlN+c7O4ZFEh8HAUqOsCauEpsF4AeizZ8rDSqcrGKv7wsVAsUGHhnBet+LvEa8kBnqxs
aUL7ojbdDpcDP4tHSm+GELDiO2Uio+53Z+2Tdc05yLGOVVtks7R6gCBFTyPm9qzk43Rj53VYnMQk
Dn053Ey8JUikPOXISKN8NEy2YUeL3Er+9gDEtkQo5sJDhP/k6byEmL6vy1NGYeMPEvZ55uwSIiHl
wl5ygwOy7QUp7LVZJrx9WCtxotCNqNdrBwfnup+lkz4PGG5WU1/5QefhEOdCyGsqH0vdQfgbgeS1
5mjU7Ypv311HnNXyjtpUltWMqsJ151TC/W6IQP69qITQgfjKahPaa15UNlY1FfJIF+nC0JKqPz0z
5XcLVXOh4c/+yPqu1sm52xNOzrXnFgEdFdDQlLn5fCMaTmDUuASg/qfSi8oi21FXykceciP7OMVG
NQpSTCO4dK0Qg+g4Y4mZ4r81vlW1QmHGI1SEx3w8+08Apu2bT9O213BMHzDS/GdwRqvgViXRlWmV
PLzd/rWoj/1+UkHF8w7TpUnqpolskORHdZ09PJARdiTIdTAMG4Edwws1B82z/9oWhzy5z9CIO5Ec
h7+ibd85ykynt49tZ8sVZBcnNTPtUPNgNhXG69NEqJBZ0X6ys8tNLAh5McqjJkC2KIIoVCbcCyP+
nGuY+VqYvATuEiM0De7K8AbM274vXIuyj7bt3dmGx/sfud/FBhnY8EEHJmdFdQ+jj+YgkxQQTzl5
Fr8QaZifdzwiTLnd/QoWeS7MsA/W/hbPYcJRGbLMQVH67EARiuidIVLiI4rHDG/ERRLVgThjyDPp
BakLgeBseTxAAbSEHQZqU+HZ0okzhI6Qb0kGUsDOzKs4ZSHTWANG536LF1F5qvooyCuWY5uBUz+I
DfTTh0srr9ww/gd8Q/0mKNGj5hnbe3PelxAkB+GbxMgPr+J/RUWpPCYr26FZuKQI0WaPexCTl0zf
UfzGajEiycNokxHNVP/wynAhPueF3LLX29r8WbIJyvK8B9KUZzwy8zb79RwhrfungCZex6SiYlyU
gGroQfMSiO8AHY1UBHfbNumaiu/15o9sK4CqDLLPTCGzO9J2WfEgCdcLZr4XbNqvkLzusqEnh2G4
KJREk+izM0uYqDMfYlazqvxBZ8SMa93gGUaHkr8IYQ7MyRLwQ7KODiX5reN5l9808MJY3eduLc55
mFDRGGdfLTd//Xd2YE1IbtXzA6ywF+XXAgk0e5cp83Rk8xE4mcA1DcYEFqdIXyB55GHMV7vE6quO
AVAIeNTueWEtc67trHTCuhrg1lEvMTip0aHr1clKekRlwqeT6p3OW8+4SEpG0b9jyBjSL3pmmeQv
ok1txSl0+547vk6+ohQvppfkqJSffliQ4QBr+N3FO+RtI18xH4H+MF8og+JmB0y5gNtugZNyLYWP
y8s2hqlLiC6HFzIGN+jShEkqsGlNPcAnc0w6imqnFKnad94Q/wYRqtfPvXSpepUaU7lUHD46ZNJf
I201wjcIPXVGlnCUnlSFO6z9b4NYcyJy5rPcn3rGRJYQzo6beGzZY8K/8m8+Wq/yWIo0DDGdCXyY
XQzjhk2EF7MeWScpR8Fiu15zqNjx7tqhwPZMj39QBKKQ2Q5KN3KEwESrePHdl5pqwXoJphJ5J7GD
w8CEmxYtxLaSxTyCqdDs8PecdJNDTCRi4Ypzx/iUjZl4/PfVoZRl41cWglvdTgs47gp2MY6aiieN
BI3A4qE2Q0QUOkSNdJgDnXRnSSfhM1/tOk0UqJJU4vADyG0qcS9qGyCtblGEtqFCZp9wiQIyXDGu
SRP+sBqd8Hieh4Hul9UB2+jdj1iihapf7dkUReXo+JhgiLyZeR595AULidAxoOtziOCAVmmcv8no
TuhmArDWTfavDTZPMLsSd/k9nmB+h+O5ppJ2pBTnm1mY0u0gOgFPWdWc51j7olMyMEq5dhW+Yvyj
388JWaEZZ6vb0a97Ep3Nu2J4yOKsEtiGET7Wijv3KJlhwsDWfKPhGs7SIxvJv8uyMS1B+IK4fnCO
a6G1b+K7PjvS5fh6Gz4uBCsZ7A8Djpovoi9hrk1EGoENIqApGcptSkhzLPjuyNfhfWRzuIQEtbzf
CeOczkoRpJVBjB9oKzp9fV3iv4KxE8GRGne41QWNLpyjnxijNqromzxar5jjZ5WU6idLmznHrQWJ
QrPNGJRbpCglhbgux60+oN8zsEc4Ju9M5rCbUVkUlegvG0IFddmK2SVoOaz1AqGnq7HPwDY7FjNQ
ZvuKxdBOIlxzK4XE83soWUX/Xcl7k7GhjAAr4JijQBM3qJ3v74MrXAQMZxxwiDQT3xzNSBQ7jhnP
16kjoeKo1FSkxAQEaTSI05QyrkJgQJ9RGU4KR5MCe4CfKETf0HpjYYNWzeaMrDmqs12p+QYIVE6y
a9yLmW3l+w76T5LPfFyMBvdb9FZf5xrn64jWmdME5MPk0gpqR28QrtVm2lfE6duMe757bh5Rdvrj
ThIjTQl+CymFUf0jwk9gaLBkyP16MAcOzzKeOQUTLbu4R8TGd2pO8xx4y3es73aH/yJEV4GkQ7CT
GqC/P4gTwBcKYzob/Lodd0aMAV1KEuTEIvdSDDHcCmXao7pD+pJJUL03d2qtoTEHX58VeIF27Jli
kn9A9hCACRJ8O1idPaSvYP4PhQG1dD+1byNCYe9ywommFPUD3RIkWde2+95ylmY+UAXgCPD4ysJq
XNBc0GHppxg51o4NxbRZTqfkMDvdijrDN0BBhVQoWFTa8N7Kuq/Jw48lNitKK1sP6M9iehknS2HX
2haMuuTRO5Pj90tCyAplfngSiXbwJRjI4eeej6W8bl7LUvUIzZMUZJEHbM/yL0533RjbNbmSrFiV
s/FEjYEfFVoRAP9LaD2g0nPqdShVYoTBeQWhm8ydQsED4cx4mxaLMstMOQsK1wvPpDbH3bDssNXR
OGVCn4/PvLHrxi7ZksMqpKRJscQZ/OLet+B+A9CKAX76CJfNiPcU01OjqI1jIqPyLIXpt9iaHl6Y
4YIyJYTkHbIXLRopUojrlCToDW8mhf/c9YRYXqB/q3lA1emgPIIYR7+PmatfxTiJs46K3ZKVD6hO
DR9RbLqi2KefbsrtHe5vg1RxgE9UTvilH6Rr7d7Qo+4wI3IhFmjq/ZMIv1nuuR3BEzd0pbL5SNKb
Kqj/PX24eQwiL2YKjSnsRci2yCOcjIkHgnIOCfAPWJod4E+qUsuYJK0ny/VuYA6Aipm03bQAezAZ
8VHrJaDnru1M+Qr/7S67tAcOYt9NJmAVN9I6yLfowSD0qu2djPKD9FPJigWOJQg2TaPZATZkm2HG
nBSl5IoNFDO4D4j7bOAH22lBd7dxNQf2bOCZDKAIuOiYURr4Y97FuO2soNtRudEk6rWfztL9VkZ7
fTJjRQZZ2bJaa4W8MyeYEMg8m8Ci7AbPxXFatl3mGyQuoRVZRGkja2SEWWC1ew8sx0uPBCeUjeHi
wDRpqyMm4faKYi26l6HT2h/76svzV4+JZ06nQmSsNELZCWAjV1ZamrAeteLfZ7WVB8mOIxgFX67u
77YuTg2UsGnhDrvXj9anwM3iU4hTDYipwFJAzXLsmdi1WtDmoD3TgwZE+b0DySFFxRzem+EyYn5A
65oqIsV6SX4mz6jrkL79GFE8HOO3fvM7slv/AmLVNEzGcBvMWY3bgLzWh8qCiCsnDE4/3RR5syEs
ca68DUpdCeqMzz6A3Y0glJRZ+dzJ9gm32VXYpOaVaX5IOIm+KqjzYKjxOxAJskcgQjbYCc1uFrQi
bcl3AvmpM5m0dyvaboQneQj3ZzdAO0zCar1zyWta6yAvYC74dfo458X8m0BHjal8khOgkrE0Qwze
Dm89eE+4wIwJPhbm3WzzkYzEsO59AaZzuzB1RJUCtMYPp4bDzK1C9dNOv41o8d4XXcEAqZLVVQhR
uRY9Thy91BpJ/enLSNkeenTl4/icKUbhToSqIA9dvDIErnJqpmzvs0kkyk2PSf11rVhnhypIFA1U
6096jlNbAh0+vUd/qEU8IOuuIskAPtHC75en+9NqhTYnF1wHBjYjaDar5fAq3pbhaD3jfh0KRQ55
tS07Rj5nq7OEeJQzq4QNF6facv739ZEu9H5TpAPdqsGHMyF4jO5+MJtMI2R4Q7mp5WqJuIySU+MU
IsYLRcfmF2L/Gwp2W7WJ9NrzH+GzQhkscH+lxnPpOv8nhyEF5XQJ7Y7B+2ickVEWDzAwHg9O3XQX
S7Wxur7Vqr+qhKfBwahQMR3kZQLzU8E+aGaMRftSpuHwpzcgaK5a2E5uVm7w1KDgIbYXqAbXamYh
PVwJEcbD4sSBHMAy2hBTo43zehg+VKWz6TWtmcUtNYq7dK9BCtAdrnV7SkVJr2J/YioJoEltcP0H
FGUzhawa5IjAGKEkjYHkM6m7WBzmJDj/qKiYF8AH6NzCcGBm5V8zK7Eb9XhIPGY92h2QbjuVcfdV
QtfkVOxpEkozgnDMPpgHWlbX3hOh6xdQAtlyztZg2sjAU7dUQauCR8ebIymreOnKruZBxDHY4IMc
Vc6P3XnDX09hSO4L/6yMY1P8e/aRbBqu8Ca3xyWSDesJNBZKEXN7vR1egwgHgAolEH5++CEuQ5Kd
9vVglggRFusoJI58zTtUtzTsBA7Dpw8/zAbTccRXFsYmt9ksytes2KdXatkGvzSrh00cXVW4noh3
3S3UU7PDvIslU2xRSIDMUR+tqUjgn/mP2oWI2qColu7zYoE0IaHHacJ1TBLakK41cbv/7ds2Qs2m
+PlMIlgx6hbR7qe+8u4VRryU3JaM6Qt1EKohqysil8axmbqA/yr2wVJ+SRbbz3cco9lWNIshmTIM
edhb9S+B6q7w6fpQJvy9576e8td3ixdKgk+vnoSNsMOQp9gXZc4czRXT8keeZkoudI2L3r425Y+3
C7UwOxkrU0aWTPr191HzxgLNTwkffOG09/Wwhxb2Co0bCmJ/Sxa2aoSKXr13C83hNb7s5NnDlM4o
bhcao8hXZikIr88LtPVi5h3eFSD15SrQjJSGxEt7M31mVQA4JJZbORGEcLTO2WAPWJrq3Hulce6W
N8aDlh/ArorI4KcXllN8Vep/uIFeuLTmN4oNnjgJh4fpK4Mcs4Ui8EVehS50oiwC/MFNvX7U76Bj
oTg1SF0uz6npWvkF45dJ9vuem1BSpZYHmACZca7UWZ6d7L3Rd9HGh8BDyzLgjQjwZhdTfBGOgiOP
ZTw1IdqMmlnzLekAYDu2yv2+OZ6BVPu1AitGLXqJ17YfzTKiw0XnZfGlRhLQl5nZw8RHto2s0833
2v4uykFNDm/D9eFddwiYeDPjnvfpMFIdvVZjpCA1raSBqN3qtyClwxq2JXrN0u4LW+PbFIAAk6hk
cJrX5dFNJP1rStijeV5pTh8dkEEi8s7eHHYSUUEgPny8Ivwl4G9xFGiji5j/sZcKmQyoJKp2LENa
t21fIfClF96PREc+GtTQFHtfjc20I4R8CDXUT8eVDUrKfEAL5cIntycXHQ176NoUi45x797mXKNH
H9JBAC5ktwqtRRNaaqRR/nGXeopI1G9RWBX07XbMUsdIEJMtcK42VboeFcKXJ3lBxrUCUtYuz4Sv
HBk10VvCxVx/XZJxvBBV1vhp8Aia8gXG4tUnnQSk8SK2e/vToRyG7JPx8s6GEe4S7sfMw5j/iMBe
bT75Mw0hgmgzibqGElvliSUtZxshM5bwuM9FyAHUiU2dZaaFcOzNGij+73vQ0YYXabg52HWNK0co
CNoxWTmsOMQTzMo+HRi81R5//+WNu/71+njJ2PLmSApAmPlkU/gC41N58YMcEUrTxHEgLLJRxza/
2dqWej/jI05sifJ5aQh0QWBszzFIVsE1XU2boC/yyqdCLcLeUYLcLLzR1kttaB0r4kKCEesr2Q0u
a7pciVdGTDdsKC9O0KsTItBKZ+BPxeOrtuCdXfhedHEVQAfrGk/UzxtvGYfa4kXEFWsOqPYhXOjL
UMBAdq16a4STDLlGP/R0BbSGnHM/EYB3YDqw0jIJ8Ss5hZqYXUxDTXwSfVf/qRtvwtsjHIGLQHvR
4GAnCFTk5cBTtfliebDh8vlMMmf8WES/btdhrY676fLNuGT1v7x7p+AkI2P85AbwPVlcfDilTsIC
L2zwzaKRE54E74PHVyQmj0tCcOxCGCAarLTBF1qCGegKMA0sDtjGXmLnwohIaCHoakuanXrN6MH4
Q7qXDbqye4wgSCp0OZolckZc0DOPpQHYKUEoyr2PYMrk5CkANA+pN0w5SnNWLXOvwGLlU/qG4wg0
M4aJ8b5hyvJ1EMll3T7HG/RX7W9fbUuxjug70DZ01U4d4LqFa/vVozFytVMRQ2mYnvsjRxdPPbV1
zDptx4gVLSpQayd0gbtq45S+fk5JS6K45oZxNXMZ2KaU0xGUvCtFl3oKyolDaPHUUutX5Y3L6oXB
WwIKTbTuN3ezkvUKiN77y24+71swLVesN7Zz6QcbOWtUCBMv9oCuZBZvsBUvy8cnBYOvg+fGDCI0
Je/hqnZ1p3N404TWl3TjJRt69BStwOL93AolpF45/1Q5nv5lEhocxHy//KlFZ9eFBZUjzW5KacSL
fW9LKAZAhDAtz2NxuHHUYZpJDpdsrOF7+3+5bAT8LUcGiADt2esLXOGtunf/8r/eHU5YKt42fvSE
VnxEDK9iYMTwhdrWfgGnaWPu5dItghnuZQbuqCVAgYkJPy7Zek6x/+UUQSRE4MiVVw+ymzNkndXx
ydAIo1/Gb7NoT/5bAPt3CMDMzoyuXMKRAYF+X/wbQXHg+XuAOHKTU/y+FgKjeqsp9bFp+NfVfs5o
cFga0TBjsy/Q8N3ygkxoeY3YfokZIpM5Y/wgdSHhqO5Ta0Ed6cP6QDFtw0PMsfcBdsUd0xbdMbsz
zmzQvFlbf1M4x4XKTDl0pWlaJ1cfT/aj0UQ76bNnSKn0+od8iU6cmYWuDYsI7ko7OciUzqvdGjOk
uCQWakjehaPRgTeotyvhND4vDnR3J1dDUPkIPO/tJI0SNF6B3xKMrJwh1WRBomGp+YkKvnYSmMkP
qZWEHt1sHuFbfaq2/xvvq7kTr9yB7WYmnR6FQb5vw8Pz3JfgMCGx/D9M/04oimIXND5fbz6UFfDn
SD5gj+AeDzjgMeQV/coPTfMFPO/9lpbikJmYKsPras3h535aStXQ1wcIxhA0RxbsxID8nlVbkphk
IkigKV/5wXzVOWqPjVx15rC3StrWJ6LrcqmpcohLhYLPyyyup0BfOfcg2PfxUMBCcC1SmmCF962N
v2R+vIpIEMXgcMLsP5N48IJ264UBDq8A6bOPfan3RfZxSBjL44GSjM0uIWITO/GfsrfqA5Kg+1/m
iNkjf2rIGVs1Ly6M1tjy1JXhylgXkkJkS+eRsz4uy2M2BJ29EtFzyp1o3OGBrypH7kl6TtzabuUK
dQ6vsCgYNiwnAStWQvcst8GnGTTRAtOEPJ46DaZb2v2nMqb/zea8hH7zESD7hcC2I4m6cVyjhIua
Q3+vktrDpdJyFFpemTezIYuU+1t0wWZ9VNVEV+NtUSA1uR1oyJTVJt/wyoAuTABvj57YL37bZ4RA
tFc3M5XczkTEprLskGa+gQC+FxpCohnCzgKk3SvQ8OukKX3AK7t8kFc5KdqZXo7vpPpE0n0sqeGw
bM6f1XBvb5m0Zmjxmg2drFurNacc1IpBsV5+Tab/Ky9rI6rwNkfhWZgZ3vkRDGoUz9OeLt+xmP9v
ukqLeaEwjWJJp4JlMuEDelnV6TeSgLumbpfuJCKDHjZAWs4pIYPcQvHjTiBgDyK4II2L+GV0TOGK
4dO7SCp7bOWt6NK1GE0F7juI6U7IclXwfhAuNZm8uSNrj4+yJ+nkWlqvuFPXVC/y/ksHRf7cSfNU
u7XJavyv6DpLNOpz/LYqpxl9sPAqYk/q6q4NDxPzvdO/vAEGKVIolKk6UukihSxLypTVYkAY8a0v
r+KQixZJRjwo8Oo7j+rQvN2z5ztrCn4R2uJybFiHpAND7o2Q2BtOLzE+cPn5RmLsVl/9/jBr0PUI
kSCm1mr32i38lamo6BqVQrH3Z40ZLuQnJl/luU+PacOhtoFg7Sk6wx0KSsGOYXAfyMJxcqSVO7gv
dLntQa3kzLSAOhM7T55uu8BA2UpZyggBVt54+RpaASR3T45D9Tptl1zhYsd9TNCnYvOx1QYMQ2rL
CNPVjTfiMEATnGkjcAKwOddAiu3nY81WWh2uGyANGn7Wjn6rfbrFZmIY1Xf1zVvYT43QaktlxuDr
+ft8X6F8HmmP0Tja/fmezyERAEoaxmcTMYld3tYWsAUKX8M/x0SBjZDJdIsjzmZIjD33zblJoYdy
qcliTxSLaV35P8eavRWMFyYZFK+W9DQuV0ATYmh49hnGTW8tN6llTgGd7w+nYEFO2qXspQ2Ux14L
+lkPZ0+Is0F28PtQMLE/FHubsCSXAZRLOeG5LD02ghs7XruMXVhjR+gxdywgg+j5mKgdx0If9BuX
ucpXBdW8HM/CgyMTrt0breytE6j9GE6pt3NH64+eI8Mka8+7+TfGK0syRw02Y1qVJeCbsbXQbd0V
V+0iotbICcMolSy6BoPsq+Oe2c0xNLr69z3rTgcri8UFu+FxWfQ3DppL3gutZ/1NE3WDvZ7Uc0MW
Pu3Si5ixr2wqV+m4EmmNcf+mXQA6gc197ifH9YCH/pmgkFZU1UveMLuhC+oFE206neGIqtimx0+i
9s9ROm/1VajGeHbbeWZyfkRU0KN8M4OTW8qVXJhoI78nXk/3d+d0DvkdKPzNo2IgTT/XqOBXOP2E
1k58L3jbc/K1hbLkzwjvRHrCvjfQYFuKUelUMCVZljW57fJvUXq2MhqPmz+M0OcqLNzk3q+6E8Ar
vMQNs7r4h6eg/D51Xp9b6klqQXvZ3nsPxSXajqfVJQl/wf6OKpgU+oe8ANwDLrT/qVsleCwDI2gI
IPJv/ykjb0/JPIcIYBeVzfdFXg3nbLvmDWttLbpZFxY4X3Y8netUOD8fVN5YfCWqiC5y02jet0EJ
YGdTBF/4iqtzlDuZJhwI87NhjT4SaOXQZ+0cosFAV3HJZycjosknwLa9A/A8oznrmiamx/IrLzia
rqlAG8N5haISydWLvkzqKHgXQ1sOJCR6Cxon1bZ55a9/mIl4ORQ3dIce2N0AM0cnKVIzdPQHdBKd
TFMjpe34MW8r6VfPwAGY0WFfwFO11FoqZds1sfwE3Tk+eRqivOnvdcg3TfypmtXH9n02Pn/aJegV
l7n6k1hfBTNWdIsock+IccjSlaafXMUAAGmPub4D5h3pyiNpqkX/eHZV1PG16Zjlc9Om5mEwjwA/
IW4oTaOQcEXMEUsU99SSSrvW2vTkFuFWSJGGSyEKbs4ze8mmOqtE1C0nag9UbOCbIPC0y630vNls
/xQ7nHJoZ9lTBnr5szvcFOLaVlU947FfoTojXv8AOHc19xmTV6T8HIJYyXMIKecykU/vCAJ7KWxu
MQQeif5vllV+Lq2IlF/MS5+SThVXRtXw1FaoP3KlPAjwvRemqtKDnYQDwPj2+9NCymyqpkd146wu
sx6KIPAD4R5Ffin/VNYTydwxEjzpB0tGfiknC1DLekd2WCG3jMQHdZ/S8hJax0ApzoGaJ0Dj+Hqe
jph8d+SbteTOTt5GB2iyFqsN7NSyFHgUu63tjqEcEy2znMVGlabZ4ULEFOKL97Rkwgs6lafuzkx9
DG1BrjsHSgQ7I/lDYwsHxdpZ0MwK0s0EWKr+sxLpo3cmWtcQvIZRh/m1JKfnfWS5O37dHbsRGd2d
4svQaVlftdHzD5tADLc2qNf7lvDPtibfyRa00bRcuw0/LTXrDM1ge7fYljUuQaqxv+qWuIr7Uy7D
EqMzFs+fjpcr2rPS2h2M3xCdYEzo3Gk20tkIwx5K1Lr0VFsSLm2LJu9SruV7wRyLBPthRNmt5vsB
hC+VyvHxQt4ojZ1KDcSQE7EIzXfB5TD4m8y9vrJHF0HWuZ5eHunhe9j3ZdXdMstNMtCC7WvkFq7h
nyTzR2mggzd4ogVlrNuawoz6TcfTl+ppbbkoQA/FResu5+8NHMfytr9BEZCGFEH1pySkj1MSGlOP
mT06C6swqSYyc4aMgDQQySa4PGXJFxrrimsNHdOb3kxXaWmEyT6YYIUTju2k/sSLquP9pZXRCfbd
CZFxM9pzHBY8LIQhb2/cJTXNu358pL2aGxuwd9m2RPjVOU5pK2hh0bjkw58af8PZAVSOgsBOKOAH
4tUfVneRCrnlRiOby5wD4k3u2sho+GfrRjKXiGs7W7pYw4sdW9UHUpJlpYuymvbMFJETKodNzjxv
RmzErIckZCN+jPMQk5Yj63OVTrQHm8tJXIjdZYdpxuP0rB8IJocXrYbuOmFCM2zNx6EcxXFfhsL+
kZI06k8MHek21rnkfQpYgfRI4knaBc3x6+B4jI2TUpOOw0Lk8zzMn3yM4XfmOt9htltaCqeGO/1S
An4dAkjm9usoYTgwDyDD7oxgZ8D6S3tqLdYlILN1GbbJD1kYXomhvw4goSMd+TkXzu1lVy592Zu7
slmPiU7lHNZDbvqfWWNtP6LUa9gKs2rG0KLfVJj+soz2SxhD64PDEC6xbcSmEhRvUu+faFibIcSu
75bQRoP31c7suc0y9vWFhG8R/0bDSL7jh238cO59CFmmgFnsmT0zqPIc8ItRjoKrXUiZEDDRDI2J
jaaIaoqR2He2GCC8bOEoQmHjQLgUnNPIJe4RHKrHfRjkxB6Ki9wD3XhDZ9lUfs/EGMhZpVCastTg
zTRAp5Kh/f+8xeuWJHKouRzeTc7IZtyxUIOIh3UmqjtlmRMyIS92nAo1tFoQGJPT4wGBXTQ17p3j
GIHzrgBH3KWBkf20iycHK+d3TrWjBahq/2H8FdqbBreN7htGAsNcD6ncVjtbT5W47wjXi1Rsow+W
Qm4c8YnavRA1fzYhL1MAeRisxaq/Zpm5eTuXdWN6eyTFESOd4x1UHF3md5V1cD93Qv5vlWR1Vg09
KcLh8i1xu9xqi1MAfHMayvvb6s/WrMe00tvpAe7g2Kmx8Hs/wmKS3JCouFkQmbDiW0CvJOMS/v7e
hTE4unCqkukAFfc8VLjA3ZraFKTxvjMSQiunE7MocfFbOE+UMjvsDeqnFS+znd8FAvNayosN1wdT
i37DWreemYNclZiqNcGJvS63Ivl4Ofvi1icmQpDGbYnxvkhf5yxCAQRioMc6p7Hjl+7dcURyZV/e
Xr18aF1dRqjErW85ORzUqRiP6MdwBvKiWNihAwUmLl53wsAmF9hwqG8cIm66dO35dh9OEqfkbfFW
PxQTJtHk/4TCvisBt38SUxKmTNisdYPsXbK3ygNd60OflskFzzMKKpQrdIJjFvaLUXSTj4nAo8ai
JevHGMuBcUx683qjr+8E0K1Ko/1PSYoJIhHkY26Wn4QmQInCgBHMZBpflBjeROh+B5E1KFabFwPE
95JT4KlSDhgV50IcWdLPwwlfwhvwFIOvQC4lNPhLvDxWm4zA3+D1NGee34IyfGdKkDvZtDXiRW9t
X7/lYkCYELSN59lDu+lxgWF/VrNB69yls4VwxAH7eHlDEPe73OcIrUJ8yemlFLprrrmGEvokjHZW
bfHuYcvjojea29L0cT1QejPLQOS9BP7kww0/pe9plJglI6EcE0VK+rx+80vGGPMh0+Z4zJzpEgs7
Xdg5op6JqMd0drpucGtSvNTA63X5OBmu6ic6jGssx33WGIkN+Zsso4JponxujgtPnY+1vYITB3bE
Ts58oGK71DMptoPYz7QNQom/DN3Fxy07oD2cdJt6fKaAoFtOZ6J9uiu2i9U2hRpHBPRNKrsb40tM
zBzShzpJf8vwjI91BX2R1r+TmdFIqwSxmqr3nhsvrgRpUYOOJM2B5Wk6vumNLkgSkgMxL4bi5yj5
Wfxc46bRs5XlOqaU1NyDFG4fMUwXa9OgkkU2668LhzUp43ubmScoZJ/mGH9fCs24bUZ9Wbk4XQN/
HEVK/Xbu6qsD9CSXNH/fMGzr3Hulx6h1GkZc/GRGq9EJeZrzQKDXyhQwdGcd79qWZaIGaJzYMfOE
KF2rf8lnzp9OIpMtTTiXb/IFodOkBH/dDN34uj4MkpJijTSN/GRZM0YmEw+qTvRMJJ03qWxPElwB
9Bw2mMiW30Pg6mRXk1GwIVcUFoFQRjwuzsD7V32miN9XQTdoac/0I0j2MFuqZ9+VCDx29euCDw32
2fW/z5pJbivLGLFJ9Se6KGA6ZMc0tc8/TDgHLGPVKzurn4ODtc7JO5DyiQ6cH4+F4k4SIzY1qAz7
DgXOapWXN2QEXDjelI8VCTH723y82daL0qk5QP7R6X8bykONn9H6uSgYC3Z2wXH1Oej+7h6FNMAJ
uUDGxvlPJbnIc5jMRVfdPyL8GPmYGHDIjk+9wpNsOQRvv/6grrPtsqxfmOohB2EXOkaAi1gkDJMU
r/O8KhYMxOZu4SmW5XBon0hF746kRkzy2oLjM+FOee3OM+VimAVZKdBmX+UDyKsP7UMSrKPMAfF0
UtM/XAyDwKUUpwoWWeV6AfxfJHJEGySvkxFHhzwj6qJvk21JrXEEBVJlj8Gbm7YMAEJf9ZjaS1k0
bS1qssjZ6kPLmo5YKq8TmonDNjB4s+4fadea5BWl9P4l4FuapnppxTmC04hye2jWpIkolZySeSu1
HM3N1l7z7dvtOt8jJfBY7tokNi0mjLBE83tNwaTwKlMfwbkg2fA0zcUgWZo33b0ye2gBSiGPycNJ
kIP/M8ClMlVEET6pM789Y2ZouQfX3bbatphzIXv0zfwXHBbwKbnwYq2Y7EkbkhedxZTwC9N0M/Hu
pS+LcGZnANr5hAb5Oa1qImYdT2suhpWNiWVE0BnOMIlPB6Nvdeq1VsXPgxduxlibDU4WUbb979e7
Csk5lVC5dRMdbtR4h8PulANqNi4xxMaJXfFf4bc5J7u9PCH7YxGCe6/OKaCuVA7oxWwtoOhOsrZ8
KY4XicaU06WIWmAPWYX9JZmdrghfpZgFlSs3gl1VgNnhHxDgTZOoMfcmY93d861r9kZDskdsF3GR
QsQqRn2gag1HSKsUJEuqUsC7KNQOrEQMpNzafuIXJbRRAB/N5UfJqhL1ftYxiHRTZ+6fZo8PCaoh
7agfjdyEq3h2HHOLJs0/DeT046xmuypVqg6XorYrDcL/bRYZ5e15jREiI6+0ty/9Lw+bDeDvJo8u
ikYMV8kzm10fCPLjDpv5LhLeky2tQ1lLfOTlcPyd1HQEYxSpPjXBjMaHsT8PtoWr54LVZNfkTt/d
AXDNQ337+iynbPzumIM8yXhrH1RLaBFpwj8xyfvpFGoCGxp/54CpdUaqC8NsOJI1pOuhF/8LDgUZ
7q8FU75ZpHK/0wQJqC5P4EsLRVlkvca41HbRuX3kDw6gafCZ59v4N1Md/HIkDtd8SeyoV+y3Qb4k
uicGCtswG7wm54YNTkvDDPw5rVqw5XOcoiElfZ56NP/UpUcNjzoWCz+pMksihMdr3h1afLRyHtPC
0UB7k+4JB1gZeR1Pebc/xuO+jaHRFRnUBgMkwuuk89ulBSK+/ixuHqVYTLjyadhJIXSGbhpkxEQa
/FrQfyyKCATpn4RSJRJeUf8QrQszUVzXoSrwnQpjGCJDA4HxaNKNPkLASn/v1qiV3HD+hAwEvCxd
GmigMLKsoDPBottM4v2OYNQ6pD27F8F43thntO4pQHkAaW5B95jZLq6zrj9Tc8KguXipRnMjIpPu
nhepimCKhQ1cbQvygSwDjT7mi76suPE0MEJWLb6S5fSj7Y5ypaPr2JTzWXmpmCbBQ2ung62+BmAB
BzSIMSBISKXuxDA9bXDnty28dnrEPg7nAKLhk+CQeZEKogNSLN3xSPxmNrHpVjgt8OBl6Fl8ZmFi
NwWd2xZk392aIH8XCSRPbAl5r2Lpc7SuB+eDz7ieTNQTLlim+j2LhGQ/e0LpNaSwg/z8fgvKSchw
R7bl6sflH8in5UMkRWm7QPw6A8ju+SxN60y+feULGIonI+HXj1nKAMjVua07o41h2WXCaux/jvO1
oEO3+xmYZ3/CfSBl3lEpBGyjSFdAY6B26DPX1NTUOEpNFk8DG8XPX9WGQ7tlk/rmRdAQSugBWRVp
gB5/XqZ7avzh7D376vEzdCU4IpafFR9MK/Ij0JPxc6LM0VIDt5/AOG7XnmHHrE/e/GDePANpHXKf
Me9567o6+iBrvwqiuDCUkkhntAlu+sK3rgIFh+0SbmDQ3DevsWzYA3HlLfQbF8PuMfA18Mlw1JVh
KZmVFKQLdJBL1zREnq4l03mcBDebVIuJjXFyZf2zq9j9kQCKCH+aVEbCOO+kEm8I0GGbZYFwf2nx
IES+n6rqpv36TAi+thIz8PCI9fojuGAGK2mNi1pU0PYn6qtu1mzx2iR0XdD6ujwGne253YKMi+5Y
PRUfQMs0AdDflhJorywUy0icA3eVZII9i6gIuBy11pc7KscP51LcStb7OzELTtTEw0rOUPq44H6+
Q7KklFj3qOBQIa8J0KtKcUJUVN/ZSx3TTtLSLUAvyFnX9N1FSPGeEewCDWzQDNAzuKypAi4OA8zp
8K+5R1dnS2smxaVqqFXzH0n6q/oJDiau8wm2TaPkQOUowxVlLXcyIbk7BmVF/FpPW2cGL1+gVoxF
zUXtLtfj1zP/fmYSGW2CG+OEDlw3F7jBlIhcKgEx/mnO3M3UvmY5tAXpLq0VAWzVZL4GvYpsWBAz
Pyov7PCUTBACbYsKn2gFJkP0FvpSO5noahOUm7hOgywb6Slf5TXh9hjgjjtFj98fPqtEZ6H7F8zh
mDZXgHwaIPL/GcssGjuOwKCkK8g7axsw+4IwrTCteYAruR5pNI3qNheq0kM3F44FtS2W5e8ZRDYb
8ZYv0p0Z3U1/I0qnMU+UNlEETbB8ZmT2Z8qhLLwOUgrq/RYAL9PMIYd7paUS4+ZMtoIadUn8AlZe
dNR6Kn0AdT3UJg41wZixairfLXd/0Qc3Yg/N1TVbI61ZsivrFJOtx4NzXqOoaaGGtTmCW032cy41
nIkRPTc4qvfBb4d0uTbRSxPdvQV4aDPD2MMQJu8AW7YBDKW4pzNbnESHZb/s+K7BZ4KQ5+CC7OLT
nJw9H2HedueLBXFFICXkS6g9CQPOQmFeuOJACPQYSPGVwbarf6IYYT06TJLEFWl5RjR1icISYeGw
0+kQDP0M68ORH/V2Qw44eJORS0GPysZSk7nCjSkBhQJPRhQZW3cptxy1zcPWhSTvwendAYQPS9/N
8LIdcWxd0pTxYo3+a3UeD/BUdysB55cDqPnNmGiLAIIt5RFKaD9nS2ii9J6q83x+qgTYgFTBzF4v
d9JTSLbbMVFwp4JywqqmGrjGLNZI2MP/IAPQP1jgDFiQyqmXR3clDNf0a3nKsCBPWa8GUT7WM1Yo
e/43cN8bm10xlQPtbX3w4fDnlOAUUefjMofnLySFez+sC/Ho8+oK0TW1HdoGd+EIv1XmFIQG04Eq
V2wT3+3Bam8h7kawvRUopeXGYNAm2q4q8+ljGic1TDVoE89bEneXISaRuEvucsw/OKN90PhTaXZr
XBVCQ4r+BX0zLzhXiwTnHy58SEieCDr3Q5RMhyp6CfL8QPwGb0zlO2bI7CTFN0l9BoChUlNFQMfV
nyzGy9CxH4m8uOUMOpvzacIcu01FMhkuuk8oXmNbAxknvEYmhyFl+RFsQ7++WyrXBlyezaG8V3tE
V8wu3OpWb1JMyb7j5fN4brA6zqx/I3EiVd58Ox9zH84NCl7zAMDHz953z9QkX6hYwCgQ3B4VdHcl
9VNWVC0plXII+3+UN9ZhueT8puaKbYHRxQzW1XMm3zV9DVnIu2iv4deMJVy3A7eROsT1i4qj8EGn
GdBgNimhuoLrDfhjqXxQgGvQn5VMEBQeni5dr5rM4WcHRbYuOndTy3YnZXSQj24My8N2Y/oXy3oH
tExd7+wQWoq0RLDgy7Z/CHqe+SGCu+FVEVq1BXVzANgnsgdqrt4VY/H1F+du6kO7q2hEyDQtvqRH
QQwWIZeLYLYw6mh4WWl6eA+V1FQlhiV8QoxXa8u5eNO68D2JHtMqRduJe0UQVWVfb7FiOJDBFw+A
JnN5fKtnJl1axgYNmGup0jQ7MPrqVOZH/UdeMMt0E4CbnirqNdWNYPlcO3792drJLZsKIqXt5xBQ
afAmO7P7FH3Qa7CCqxxn1egnNeNaFVU8kisS/6iC2liER/iI76NKg/rJOIEJowXInh/3yM4ENxPV
ucLQEgdECMiHxI1gZXFhS7MYv4sTEbdjMAnuwtgsnINDpRzVa/8V+EJEQ248k2wbGbZ7jYXHLexQ
ZKYTITf8vS+DvkXFOCo9E3WJfs/oWVdkilm4GsZ1bi9DFDlEvZ2zPQKn0wsY8Eqm3MzNyRI8mdMV
Tj9doHIDcPpvW+wam6VA2NtHzoOgZ3m8UXPkpeNr7Ig3e+PBNODqxsrosVmVbzC0BmSuv/Bf42AW
bNPhsVCaAOWZ62e7NVc8Rqf0YTT3rReCp/R3DXoUtGw8e8O7EyekxNiAwGsmoZ7bnAhJDf31dIK0
z9smGy8i0f7ygfa3TSvxb64y4WkeaMW/tIdCTseN4sV8Z3mwSnXyESg42awD8SVJ/1UvqxWaW8SZ
emrMjDKJo8kSGJ61MdvBs1M6d0l2DOEOfbjagy27CJLj97paepwd6bxvHcUDSeFg/YAgqR5Hndti
EXF4N3O9mE10Lb0pxIvzontRN+RLzTh1CrbaOmltT1vpzznIspy9eQv/hcKhe3IFWbQ1bAlorxgp
XmYjLQKhTpA+PFU5HuG9spV4s3/uW3SQAjnAwE7+s2MCt4+/5aAucVfSHD1gpLNXLq3r3X1g2Ir4
lKRhBn3HeRcaEd8eYDCx/CviuIV5VMU9uYQQ0wgR9JnkJ1FVXdERt3V5FOqZxFJ/9VtPXHGzmLhI
NZDD4lwLFemOF05cCip9FpF8E7QQhF5WRI0NNThCpL7Ux301O9PjMslFEOBZaDdRW98HALAIGvId
UkUdJ1nMCwvKaG/wv4ToL4MZ1biqQ/xdQLnPbM4p8FGlDBoGuOF9nhfDfh4xwY7uJHA5m7te0I+F
UeLdJVKVjkHOw+xdxVh0TSU0TDHX4p2767bS/0Ww8h/5NEtyWkXN62E5MOQ1cMDwCyHWMNdwsuET
ElL219zWUiiYPBEI/i6z7TGIPUurs4jEp8dBPnVxuyByF7F6gtkfyoxEK1gt9W0XhrXSYyYuQu2F
3Bpv8giXgAaqZCvYyQqiU4K9syFswv+36jSc64uj48r25ft5dqLFPsXvibXdoKdILYjh6U9WeOXt
b/3iuQZNQkXHoruj34hZO7mXLV5Zpp8m6d0ehd7g8z94Zfy7vb4Ozw2QhUOevjyHFs/xDqK/wC1f
pG0p04e1fl1D7d78e2x7fyO5V0rBlE5DpWxVt6/lJFk4btJ4QMlznLb2fIwCkof7KsOPqYqIo/Ly
Nargq1vyI4b5Dv/m1b1po/Q+Qh6/90L8rVvx4nMGGn8klnIEoxQW36UGD98AidyR/OeQb4A2TVh8
dx871fRtbxqflXsD9aHXOIqVbmyw/TeVI0SbebjFPNfh6bx4oM476gFSysqKlp7SKpjVlQpGDfwX
+Ydui/nUkDrAhHiXp+AhVI+/C4sXImeyEEl3v9jjBvHHC63b4NtZSQ4y+ZUaCVo2vkx+2oYjtThC
1B/OfCp6iJy0xbsrMYEFLBygavcK/2/3bczMfa9yEddjNfapSYdXsaEZN9ZG3QylEt9EXaUOuuef
rPuBNhB625iYly5lilRKxlfBtxoCFyQp+byJDK9QasoAoxiluB+KbuwgWqOFeImoAQVcediFM8FF
6ablbT+DEQ+bJyDewmmx1Jp7cNKnm2/hJi+Z1ETjgRBlmg6mPfz8gV9UOW73sjPrg+NDAgqqrglj
+y+iuljG/jREqsrkqdB7ykoiflSf3AlCwTAqwuNx4LiAAB5/fU5YS6hmAD3JOr6FLRmQu6ha3w7P
ZOoSr6SvucRLGGy8JG0GcsE6c2qNZt0zz+qxH86U5/t+l9I0eTFR+bayu7RhpntfMT4UyWX9eE6o
GEqauwzaFIcnetpkAzRsHHxsO2hgLuyYDJRh6pMRCSZvQyUT+eHg3yCRiVHK9MzoNf2va3sW4dAd
3XO+wFEdGTW9cv9bZjwOmsKz9PAH2uTG6ITMkPn6nTtH3Qq01Wka6hD3QgmuUdQWFUYid/6qF7mW
9tJ0o++zGXg7xDu02gtCxq6aHGO4NJs8lt+rMNXhMAzwox/5MQu2cljObC1ZYRtV5j2eEfQwTrHC
0CAG4G6oijAkNu8MXeAvdV1HxdNy6z7nv+VYmX1RuoApX4m7PCIkx0ZHLnJ8GVnJz6MBDQSCIX6A
WbgHabRf8zJQauRc2mgXH+GpaOYdqo82lbTPkfFwNVAYNUNpewdiZ1MSZ1XEAavinqvCgz/kK20y
Bo/vVYJ9t87QXjk8eYZEv+pVgd1Dfsdt7xiu1Ci7w1I5kLExjq4t9AbDUPjkC4sk9r6crdQ2i/5b
a7Wo+RPWs6LwH99Kbut+H6ZLHLawm2fmFivJRUNd9JtuovHzECd5vklCm3E7HRWnhfaFtj7AewN+
D+jzH2GEFWInN1+aIgKTcoFjdpzbLdbtEYUxLLn3l01HZZ0xqe9RuLaJFq0akfYJa1oOKYnB43Io
JHBzJRKS567FH5gxQlJ0THy3HOhh5jenKOB4QlGaSb6HhEa60Uz6ANSvqiUXTYOsgyMEuoMncCJk
yn4DLJlMO3aYwvttJpxowyqewXKNzB5+TrRhivhCRXe//CSkHmzzeXZxstFxpW9r/MEZqZy9nMn5
X4yr6refTNxGuZINcBhx/JngHVaOSNEcXH5AE9UDkiaIeXVhTzNLfoagL1zgfGoWOWC/BUArAQDn
vrhDPTv7/z4X6J1EzvwEeLgvnTEf/ZVN2KZfqPb2G7JsPDPaP4+Pt1Yfim1hHG9FAIuF5AAaQH9Y
rPOgjT+o0cZB9FzCJCmGrPoMuSaGG/kELEXCAvgfOQP8dRnY3Y/rGwvl8h5zJkwNkAV/f5fGNpzQ
kq25zoU8tYLKXZPUnplS5mu4xtOWYcHF8VTmon5xSE1IShpZB51K2Z49B22kL0ZlCgnnNY+TtMOP
BbtdPVEjHUarF5571gySSiqlI1xp8uEFc6kg/+oiHQbAT0Dp574Pbo6y7zDu/Tl+9t4EOH5V3jRv
Zt2gpYK+Cg6uQzCA0sA4EDE1pYJ9PqFNKN1hz45YsL7s8tw9wMcf+GZf+R/niuGGoFfI33KD5G+L
wWM5FmEx3J9HXDODxowy1ijnICzkBrSUO3DXSPA4/Owu4d4kiI4uc1ZOmmZJO737TXEyPr/Wd7gO
mLqj1QwY/HNPEq9GxvWle023fEE9fgKxn8hWpIa/gLQ5vqNr1DoixwK7hXT1bO2Bdu6RlQgipAZG
eBmzapHU5ExWCRWeq3CrJZuaWvsH1t673DSj8LYS6ymL7nMmQxlWQEDqYpyuRxDfRnmwY1wPwFcn
D2nvP9oV66a6YmXlLmrD/+gCJdpYDJuvIK4Nh1oo+SpvN79hkE6T3/439heRmJGFGzYTdQv7GN/W
MfZs8CPyTAdjY8EoqbGrL0WaHRjomuh06+69bB9cqhQxEGlhff3GBy2lpJZkRJcOFR8Uu9Kmv54H
syYhAxHm6GC2lWlRgagzHEXKUsUmfnHF4j1fP+3fDjt9eo3ARqNgT0iLUgMwKxnJoJKOKGs19uOb
sQ6SAxJzame97GSUAYEfwr/0Dj67HaQwjxydTVc86ziiMvB4ZccR2y1YTSq2caSB/yzwBICxSGI2
LyTg3JEpRZEIf7+Gfc5BNCG6a3jATjlgNl1jDWrynegTSGHZ219gBqYBsEDOcXOPPJT4deBpBcDS
oAfzJ49bn+cgRXlj5EqDTX35irz4tBAgUMJbZPoaTy+ct9mXR9hw+9c365H4ZmC0KGpFb3QyFzOO
pDZQ7biIGc3jsQdCYLuzX30pmbVgavYlLLAsAhSdnJW97m4SeUZUV7MD7Cnmr+EqLVyu7jg1NiPG
RrJAvve3UvgpeThbUY6HrdfF4HI/PHhhVsaXPYoSLXSYonI0uAu4JBFNsKqK8QyagEOawF2SE618
x+GXpPU5v5XD0n3Q2HmHSBoDeB0ietG1BG8iDyLYeK8m1porw66xgqIia5PpgXL+CsusYiEekGQH
s3nLUjlf/sfAF2yEvwk+/3ITLElTMbxBVdG7uOQRTaE7zy9vkxgLWVE6Qac/HKkw3utLd2V3H7Ei
AC7wWhsqLAiF4tYY4kNjCYKmhCdh2dmjvTI9gjBgh4eQ2RWwjvOkjr3Owij+fyr5dh2at/oOzADL
Rv5Vg5SqfZORaC4ud5pVpkyY6/RaLu+0QjkZsDcyF98tZ2FqBS5UW9zQt3/7s9OROv9TnR0dr1yq
snAkRTmpfxz/IyVnYmbM9DnEAu3Yqz4xyMe7DMm8c2X9DmS7g2mF8Krn4BOgALJQs9KDPwxFBjuB
he/hkG1lWJUnnYXIlMWCxM+QaXk/UFhCMbtef8D36fO6xWcWwrn/pQzCd6a3eeembVWrrk34zq+E
1uiboER6CQuMDDvQrNvJGjkVOmVedkdpgwBRY6iBjj2JVWRv+agELvuLx2geOTphOGE3WizuyUJc
iB9BzbFiXgL2+0wBWD8qKd7EAY61gfvDBz3uVuvczJyNsA5pB6fWjTV2oaO5deMJf92Qy4rnqchs
OzQ7XJZJ3bovKgVPfDvrHL+gnXFwGYq8v3X4h8ecPIxM0BKAZOUyyld/SJfZm+y8SbswlFjRyq7V
ZoTxqAVKnt7p+E+0H1+ILLwL2pSKnwcRdfGZVScDsEB4s/FI4avU9jEqyKOCqN93jEPAZSN0LzTk
fC242IEUCIqmKiW/Pj9Eks5b3ySBNSYsYMcFh8kYEJblx9/uSA8W8pqmC6GiMqyUeY0zeRjc+sgq
7SdDU0S7HG/cfmhHQXE5NevaZ9zB34q/o5u86n2uCfRqJ5JikwJsVTNBnfh+KzOQgbo6bZDBQBFm
PYu43tg3NN0LuCgA1ZDwmKtE+a98bv34xG0wWZz9HzcNP5v/gFVq3ssaYaiqpSQFwhoOPH2MS1qY
mrRPzKcoDYeIZkgTJS65o3ny+QoDdwgUEJGV8lqpFgZj+3zC27iRKXZ91O3R83dcHBZM+EuRdufE
xIa/YS9LoGEoeImjpfmTp0WWpy0qmB4ElVxItPJWv59mokFPo51qlVw2L3ATUACY3MGk80GETgWI
KJWT0hnzHDi2oQdw53xjJgBRgriTRldBauBJyDotk91YacIJCihkV85JmbYdq6N6Jm5sSEw4n7li
rQXX0lzDX3n8oaU8ieVEJAq+G9frJxL6MqBKK5Aye/7lxOsyunRHE8J0N/+vxuJTZP6g+rxJ9U0u
PJKJ6M054ruWc6VU/Ei1den131R8WuoMEEpQ9a69k1C+cTbaA3aWcuNemLWYVvdlgroiHBlOFlzt
ipwMdf+U21c1YIIb0uMjFN9xgXHcImw0u7FAPh31KrTVFwBCcpN5hnte9XK0lLTJZDz6ihXYQsSE
Blqk8KaOA56Yh7Oe2g/Qd1T5D0wh7lMeKPF8bt2fx2xcxRHtbypKxZY25gd2uoPtB0yiOTJylPWv
we12u0SAKEnhlMCfdtl7k0YAJi2RZRz5bocBH+MrW9R2wxVUL/qTUCgCSA1Kzo3S5yJ+Q6WjypNL
Xe6JRK4IXmJtmUWqH/jkiiVdrff1j+KSvibiBbiygfo250muu7sXmNdvWP9lINRV3/NYf99bysuP
3fPkGYXQuHzPyQz1mYqu54V62Q/+M/0n5BQWSBY3VyTjoW7YrzCX09DOlKc4mOD0ZKq96+IjLHo9
OKo83mVrOnyPiHun2kTMB5G+O7qAeLm4ZaLV6uUgtE4q8LKfQKxcJIhgs1B8lMhj7THPPJ6n1EYf
c2+mN1lS4RxRRLhfX5EF1rbKVKID0q4ezKbBCTVWlzMbgkGkxiPtSLKS/sxqS555anhd4qQ1vRLZ
sqc4jUE7dUmt0aHMszN4rUOZsBJJnhMXc5HCISmPrxrvu7HjGqNnke8EG4JonIFbVzQ/iT/GRQ3d
yi1wzxfkPlwrz3sww7+l1b3J4Arob1Oym8hWA7bGVN2pD7wBtJVBC/q05iJ2Y98FZKGIXz6YhlFl
c5o5DXdWL63y7E3dhUrVrud7+MZcoiWJJthzmuVwjyY+euCIgv4itpC7WbrJFNWEZNBqXIc1Dx4K
TWwbCsJFQ5KSzux4p/TMTUQCTzic0046N2cjWTtS3oTE8UiNC6FtqQuy0BXuafwUusQ3CuspkcSA
mviVdV9BJfWyuxidz9hg+qCPrKLGNmBau02J9yvtiD0EK3m7e/GPwXTgrBRqPkDtHhpV/+vu0g5N
1Ye0RjBUx7AKQKNGqTgEAik1fpOSXRjzTqcma53uBrmgui1m1CzpkzZBB3SMMO8M7lilNc360QY9
ufcqDhBDwK0YdL93RhIbGlnIsvUDMcf1S5IDlbLC332PiyEFWQ2aKIOKUH0K9tRg8/GdDSrvmKHq
F3xEhm4yY7iHLBlEaZN1PmkFIKRQUk51jLI9kdJNsuoeWgvliIL0242AcPSLI6nJfhODbzkqWwrB
kEk6+ZNxVc9UYJGW67ukcPqrpHQJwfoci82fxkNFHsK0SxXe+Zm024QcnagXJMcYFJPvJzWVfLCR
18KXhKrRaB1ZsjtfKdopaI5lY+K0rpIpQBcWAsbVCQGyb2dennU/jtxKX0KlDkf3d80S9HSz0kUY
D+caZAoJg4bhiUQwcaoMxHez+GPPTd12rpyBo6twRtOvweRJ+/m0i0Wk5114lM+p8vcf9yRDJKpb
cAzHGlHnQf6PNrMpHB4NBOSAwhKlmq58dE5obQG9teiRQw/spbJfTM4oSl7DdB51My+AEprpjOqg
Ld7DuCwmkLZXU9zwzGp05RU3WMU2FpoFxbiBicujlqXb2o70dy5tznkmWdt25szToSSYIFxRBBsI
NDAm6/n9d+3rJS3duCSapOczHhp2iYTRxD4z+dwNpjDV0Flbs1ocORWcYXxiwQbhMvfdnoXqGmQl
0pXN5vIsIsh3QYpQxi7aY0GYPnzboecdgtC8kWsHEPAZZRQ0bTlm8hq1FoQ8nN/PmHAySaDFPqXl
kpcR8t0VJUSh8ghKqV/0FK1LQu6I4dYRrB6wjdjcHNPC/mcNJXsmBT0ms5FhXVmGibsLU1ZgfSyq
Wa7FYacAjuGlmIyanRfYEOPFpu88lNR3BSXmeqLYaL1JwAqLwRLZECtaeJD2S3QlnyvzlVXD6XS6
7q3C3YB9f/ylM3tbkOQyrVsRJKnJp+3CHO2Iq2liVJSiQCuSS1ginBQOPx9rRlSriTfveyrJ0kfc
CyMZGEPuD3yn0D+27DfZycX5nmf70/stMPsxiek3aZPco7GemDW4H4/7ZOlLVo//qyqQ5zsQ20S7
NxvZulnSWYwskYy2kn0uS9C42sPg2AXHbNcBCgpoMSRkw8e66o0CHFok0wRRQYMy02FvN0/QyybS
HMrT2znKHln7Svoc3VJwvl0il0hRbVoaONcME/bTAcgN+LcvIboWnWha36x5igvYuD60WJJdP6pL
h/se8q0wnJeA7iAX49p1hBFKvlmJqUTzLBWn0RS9nJTIfvByta8Ajzjtk/q6Ly39EEcjzOmoz5cz
hmCUO4NzCB+QAqz3XbWCdtcBiFPsE9kELScnDaagsfLegIAL+iRdNCOqw3p/XoNf3f9suVpGdECp
MxjhWowvk+waffbag9LcD6Ok2oWxnTQkkqQ5+FfPIaVshswa1pU6QdQlDSP3XXNGGRTqUmoO/JBM
s3GEcsDUppjmt6OzN2gmmKriWDy9MNaLDp7FKGGFi/WPdUfd2sr6l+saYue31LEfr7x+g1Muwi73
UnEm3IxGb7YUdEfim04Vcg6N3WIq7evCgYwWJM3mnkX2WHi45/FZSVuEzkkEEOafTI09wHt3S1RV
awICXcWR397Zwo8Qi6Rw8EVxeDhJ29MWme5wTazoDvFZQDO2NJm+ovOCS/qSeO29NGStZa3VwnIE
lYPaNcKnYi1cwmXtv1VJ/kbdzkA7lThzhE/2PMplGVPtYZkZG72+XKfFazseoz7vGGrjIyKtBBMq
APM4vLflkWNFW/otMLFXnNrNbjAGO37wQhdfbSVN4nZa8jGs6MWN9eabDzT44LKdwsKShyVo3T2E
8CyUm2LmTxURvVm83SwVQZkerEmt7yZLJMjkJ+HkHB2Bf9w+VtaFPnidZfYsJXiQWys7XoVP9Agu
DoJbHNduUU8LsUde6ck51dlrIwXUb/Aa1XTHNAGXkJFftBZvc2R/Oz481civzAePeWV1LmcNQp+B
oV1NnWtyf3h/NjdTmiAe7GwaX9NOo7G293JUNyfFTxb7CBrJhYRCgVoQWAmmvgBrOdlnmkUqOgnT
yKPG9/XNYho2pK8TgPfSm736v+0goLF7pw3Ukm11TzVPW08IOLSrrX4CLSV6a8PJ2Et1NogBAaav
JcuWRAKG/iMOcrVmu5WeKDNSnc2C/vMVOUhKJtJXV4ig6fIR74qlogjsV0qge4gwEcD9CkI9h+Cy
MTajRee2lsJkRWGt+00PHyJmanaMn1RX1i6axnBwYiYMUqYaSbVq7MGbZeFnXujgiZawPTRt1rCq
UYTepaFJGXGLX+SOqaUJ2SMOsKRxwu3vSiGTTXPz5UqsL+ltvXZOHbsZrscy/r0OZ3IMYqBoRJ0L
zMj7kuhzrQxVkzhM9uDAtzPN7gU5Fxp2cQCPUE1v/DnemuvP3R37kgS0lRRNCGAzg6DO3/kELq/w
D3vYILJCoBIK3UZg8CatZdOQCEp6mDVjZPuELVyfit1AGanIRTNcTNf1h6ontmbIqrMt6ZosFbnN
i2ZBqD26VvfKO0IXYDV2fTl0F1Y0NAtnmKPqCBZjA3zPg4n4LQpPO5SekVrVae/Pk/RhXL1XTXeL
mUitG/PNj86d2lyU/gjdF4KIjxtP9zlGH9ICR2fvhwHtBu/XFNeYkKUHV/hXzARiUtXGpa0dbTuC
pNT/aAw2Fa4BELB7RTQjeXO7KwXI9sE60BUgqXUEaP2Qaxe3H271kj7a7lNo9nRvTBm3qBK68hfF
C/mfWv+I4j3rrVC821OU5KodjHd+m+vCkmFCaj+TZk/Ua/Pr3uRXK5JEbAeuTvf8o+F1aDwTeTKc
qeI11ujEOGd9P4DUkLbhHMcQrWraoBm37TmnmT8rqIUl00GIysCWTHZO/38g5HfbuGD7J3Mb+CZU
aCYGE/8lApiIBVXzf+8Q37f5I1iARHOjVI1NhXvGP6JcKqDd/5zX6gFdKNHpQW3t2xkHlK8e822X
2jEZwUW7LYOMjwL/eqZvkc1+Q9He6pZNva4fnQBXYhxNm6zDkAEw6bru0p3+O6iANBAx9U4HdOJE
4BqftIjDOycbwaJp2ie1q+90jz96D5ioudiLQWfdrzOyeBLSmtfVcXfW7VT7PDBv5nV0HP2k1pD6
GGK24H/j6PNxWQfKG2XjD3eKLIiofvMVOfqZ/gs+qby9VcS4cI+faKj36s4DLZogGApfv+dACUzf
qQu6PpfzgKZSDwMFzDv3OyBPBPHETLm2kj7cQB5kmBzV0+0+9SLkWSErITmaCZE9H9Ca+eWdGSGq
pZ1jel275t//Gul9YdiGtFDBnozgRDUMDMLWTl7GAe9bWGWqK2dTJFCYeAtKM+qVqhOkDZDLHw4g
4FrsLLCwcKOoYhbb6in6okYFwgJuMDJVW+crjSfSoEiHvPreEvTeFeWsEaAxZZcBzsP8ov84PqwF
jh6CoVT0xfHJgqtnNcM7pxCD+XJx3Vpqk6gj8WwVsj/4MjXNdasLOgGJ+jjzVNhseAx19iK+W+Ds
HzknNJ+upeW7D6+YBcy+8+Jowml34QibOC0surjMrUPdLq6ZOq7ne8I4sg2E/ST/1L5/wQlBj0eR
bxMs3Hm7PMou7qqTFlqCPkRZFmLt0vpZAtH24kbbPQ9HTl5kHZvdLXf+hpCnnUYrkOHoYMAdM+Xt
wyZb48idPl0MTwGvRIvLXLu4AJuswZgSAo6je2/RujwtM+upmAzsZ7Ymp6T7LbA3jaSCCYsnpOx1
ZV1dlOfyHE8nXVEhebxIT7xBhfM6O30tg9SOgZ68eT7ULknbkQN732ObxiuYqOR1JkBdS+zA0zqR
4qFi9HILHkTj7Vw47jsjH+syDX3jxkFO/HAjEKDhi2ePuaDQIdTmHj0aHVtHlXxhC+NiSx+E1ssi
tvil1OWq5fHNpX6pEVqYj2wvu/4V7K5OwakQ2kLkIDEC7qNDG2hq/7Oqbc0JZnXJQ3D5YEstBbwU
uerczTLp2OWzpmeqRBgXoxUEltlyGq7meHrusD0jc8xAGk3WgwrXHO1CPiom8ZCufX+Gen7cpSqI
Fw4YJQPx8uShxTffNqo6n1RoEHp1/u2FP20tJ/rt4YibfrBU+tmzFvCtKExyiZIIJhkyl4Fb6Nsp
Aa/vMAkOYw7eszTBjmdTVbfR1sjYeyP6o9mQb55+RH4pf3PjC6CnmKqaLrIDHdOl7PJ84qsWzkVp
7wBTnk/0mJvPgw5rdMKaQpUgx5dARilK+nR/B8OFJu7C1V94ePuEqVW6iKwS0Et7LPENeqLYdC9l
m77zpgWUA9K2Kum4AhvK7vcBvmfOxh5hMB/EFZyl2oGxdc3pPGmDA6tC0z/umvUOGabyGdXqtqEP
EMF9LzempQzQdxflVSJgb5VbOpJ1Df8BfKtaog0qPrI5+KQq05mX0bQE9EFuX2g32456n+WmfhhJ
1QVTnxquT7n7pxrdifXv7jt8axwLhrVJtfu1WQNMKQ4fgwSYvVP6tYkIKoo9RG3dgTgZYgKSKMtX
AMiRmjoE9L2xCmtdULq2zURQeSAFPOO/DbodfwUcEkfafzRYzU2+hE86emvcMfSqBM1Xd+0P85RX
MngZ4UbntiIG1RcETFQrsD/jPu9cE1CoqDMXL9XY8tFqGP8W4lV9hhMREcgrwryq0vPR06iK0/zR
+qkNRPEuH9rmzhAOR2NPNrca+Xx68cZPI2qbo5zuAG5Tm55AX/NHUCzT+E6NdC0TbWeL3KJ3PvP4
o2COuVT4wfldr4wWQkLso4y3FrVcyqTNuNFtTgtdvpU/0RY/LKroYwbRFx9G7mjduypZVuixLnkh
psHloQVtJ1PSvEEjQAvAmZ0acaFPsdV5nYmsphXXWQrxbJK++/VSlMELd0I/yjDm8getd4p9jM2T
MmbrBzFaxOr8qqBs6X0NYg7hnThtLfwHF7mjTPldKRkCqCCZXv04wrUX+WxiL9DsGwnPnyAdRjrI
+AN/QLhoVHZeB/0ZXvQeBs4A/bE4uU9Mm/yDaDVTlZvnjyPGVjGUSi/zYdRRtFA2asMuUC1v5N+Y
mMEU55idzuRhbTmrkKo5S5GtDpzcGgOvcsQ8hhyx2bZoUqlxI9a0+6+85Tg5bwO4FStg7zftlOH3
2Fi1vH3M4nEbSyMCqw2ykbforpIwxEyaW4XZhSYUNZu+Xq4S3yJ63CCLPsTr3aO/TnsPmsdnOgBA
liI3wP6LmkzHOWhTYTisBs6WQpV0pu0gs3XuJi22m3F/87VJu1YIetGccMQdOsyTV6HFO7A29ksE
dR2kF7S6SsQh4sBhgNdpq3cWmJOKenH2bUK1q29mMlXkwr8iA2CBK/I3bJbjgemdgDZiNT8jedM+
tR41UFzi99nBWRQRXy1Ud9584bQJYkbKHJrRzCYwoKDhVBM5smDwBHQzUZb19GA2crf/DAP3NGWr
tHL3P22f/yt/wKlf2/PWW8BdvnCSf1aHvBDDhhJVceL3QNz/i3PfyI4WcXmQWqcsd7KcxO2Z/Fdm
IKTvbdFsg11nRbLrJRh9qQ98It/fpeiaP8b2OFVe9A3uJns8EjtItYf4hdIi5i3jOjIxzpNUnZ1r
fH4cL5HoIDSV4mEZnG/L0sXfVuHZ1ssxJD7pE2pvTtIw2rz9sXuXWwaqWHnYchVFi1FjcMWppvTx
SyFnZmEV8l38kaTLRJyBGweAKZTdGRc1u+sfVRh/5XpWb2g9lFyYLaGC+7w4cnE1+8kNeKi5LCDk
5xK8AGUF4yWcSA1Q7z9ZyYTDNy4oii6EnMTMv32v8WmOD9zUur5OegjOLIPOYvEX9ZawnaburiZs
YVE2J8+Z+ZHyHGkJcHl5gBB6CM69rrOPlV3zL8oQVZKxtFhudMd9/uMu304bG0mxpGAySZ5dyPqB
bW2XeAjvGhiEGFmRZAotP8Wk/AVEMlWc6BJt83eP3UmVsMUvDjMtts7TYHtGM4VyBqwngSvXNB3X
bDCcGG7hmGq5a3EGUDEWfDbpBUzv+OOZX2YChyp4zEF18CirEbwJrOGPHTuDcTJWUbKOvC6FOecQ
Y58Ecfq6ew+VpEf4JLL3eWCbV5tY5spMyl04zawUSd5PEC4/VBCeV01NcCKIOzB7/jB+L59aTmxd
O/3RkD4UkuXdn4ZJ9w7HDA3Z5po9aDWsQAVfbhelNMh5aW3p7onvxF8ULyCsbTxBkPWtyRHUza9b
lOaYWPWhO8XeOwmEL3mqKllyAZIM7uS+KA6fL06bvQfDK3nWdz82uK5Uc2s4rOqTSLTosAQyXyvt
EoQfqnjSEbf/NtXUI3LODH5sKLfr0iEq5qnGx8CQ65kdxkDNhez7hNq+C5qb59TS51KaoKBKAPGQ
JjyYodnA2k33dC1yz5pEjugKW7iXSnnWC7GcqjbA9QOv4ndi8s7erhbLdDY+mchRNs+H9XVwiQ05
lqdcXZF01YtkIqsXoAAozYA3Wf9OhPvLAn6w7hDkpnJdluzjgWu1hmwXCunSIFaYO5ylwxssl2c2
yTPfawMJ8kXwZ52cQA9EzJMzAzdjXspRv5Cxai5z8XoBd602IGL5pERLgwEPWSapD6cp9oZwRnar
UpmuNzPVN65wNsXRzIOdmKMmXFdpZpMLP5U0iDkslOqhDFAFJ5Zjl5MMyOsLNjMMz7K0hZrJJaEb
BzDycbqYGF7Mxq1xDYhzwiSdSMR1xDCv6CRMu1GB5tbTee5Ew0zJmQW9OBbkT6UhZ4CSMaJ8KhWT
uMC1DXs1oW1yisB+PD9642/nNj4LBEig4Agwo1oPSNr/eFJ/QMSB6C6SJO74PnZVyYxfL7aXCkRa
LhSa031iKWJu6B5eALnX166g+QM2SNUd+WG3F90eroQqLClW7ikgdJZJxvaeJ7h4ar9zHMRMc1q5
Ms0yicdkjwGTAMUC8kGCO81M7/Ru88dQWrZA29AXRE6JeuK2T8GlBVlom0eTPkJOLg/5Yx8sZjof
bJQCzReN8wKeN0TZbnGyk9p0bjaAcaCWk1LJ6QT2qdhocI7DQFaAXHfKFT2r30tvrXQjhwyt+Ox7
Yd7tC6xZNTPKRzShw/vYz1AdqpEtq7Iae1X8YqquozOqcm2peT1/MnQtxlaAFAmLnc8xSLCwLu3T
R3UhBy4a3HAetrIB0IvaGxV31lE4zXRY2nfJUSnyr9VlJa9sTkahjLb04xS+yAWnukpd8NrJea9s
/QycO1lOxKk/4zMwyYczkBZMkdzvscjKt1hkKmSHFmYb/H6VoxNVEr+ZtObedzVuDXWr21TMMrDF
M5zdHwKlgp9R0lV6FTyZIOfR8X5nDAn8wNMtFypoIfRVsyNPP1PYq8Ce+Z4cxFS6b1d5+oVtSZ3z
3oQ7MfF73DHgiWfthctBt/GXY5PQ7isQauL4fogC9KeWgMC87C6TBnnGI46RCif7C4Tj45HpleVz
2a0MJV8zPfOEmKeBg7X0uy5p83CBbJuXA2EyCHiifnR7kRa7BvF1gRnE95MBnmtwEQG3vDkDx3Av
99qIFLvl5RYrD/kxlO6PZkDJJgPSi9py+hTEwZP8zykko9t0r/iksJljOC5k3NM2olKQzUsZfqWM
4jC9ylLcyMBUPP40OntOZV2pZ3M7H26QsCF7kjJD/qlRP9q4mT3xgBejBrJ60ibRlAbAIl60WkXf
H5lrmpejnTc4j96S7XkqN0Jk3Y9dvXMmF1wlQwKTAmJgffsq7cQ6ihYENHPdy7JFiAZqhhDgbWY+
Ae4wblIoYtSMMqn1TdxUJr/5bwY3sSHu8tUjR+nL4lQGx/F0R9giOwNA8MubqA8ihNMhXXRWrB1c
Xnx+1qkBtJOp/PbShA4Zh4YoSBVYh0hCVM4jD4YAyQCLyu6pDT+bBluJQEYsGTXN/F09x9Yy0/7q
d2za60A4JzCa/q/uzIrcwHKrNdna4Y1b1ZCNVMEsgJRgljSX6e+YuWn28RUQTPJIUUHWneusLgbr
9zDAO6rsg12nh8Ak/b/buP18eIsQYfTGTp9LNFfgA309AMzG5EcFe7Frz1O0EcPyJDPeWU6polea
mLotsyUiF7ahIrIc4pxgiPb8BnqVn1uOFgvcryOMj47dzK6Ghnv+0TKNZ0QnsYYKqGpgTDANkrMu
9LE5Uw3cMfDr4uiqfhGOIqaKcwkNE5iQ19mWfScyZCesIwXIzRRluwiDXhK98eLTRZ862rgzvWAT
ozn6Tv/9gTfCNBsACqr/mxdY6ymPaPr5jOZmNetFbdEzhHX1dM4eJmA6CCUFd4FunO9XGe8qsFMz
/l60XGHYdBM/jkRwwyo1gGbyc3iE4xTILgYb9/9Fey5YAVVATkhmTK93CUdHLmkTaaDmausBEKPM
C2YO81CyVWyr319TaHx1rMbAVBw9Kd3ZbIYiNpdGQSOAUgJZD+xH6nv/wdH2EJnX6QtywaKQOJrX
GG8MEcYvnk3RYPGlM4EKl06NAkzU7lGtBIISEKXKCFiL27cdPFkqFWQQ1EkwvTLAQVRpiVDY8qvj
nSRME0zIiVtOOUgtNebpCsIV+PnqgmcB+bjilSoSsCdTCaONO0NoRBzcVTYUWZCceomr13jdwfgc
psUfPegxjxt+RaY2Mq8SiDXx7XbHJfbzIO07xi4ijaG3p0LpVUF30cmo5KLNhmbnMtnzKQBBptU9
YmvDxMhdIIch1E4bjSh2F6VKL/i9mC6xiuyNlvBqMT3YeGpwJDiaiuS3WW3WoU2HCEJQzzhsX4Es
luiRnh4fCLT5qrcDbTn6ZfutYH3AGcvnxXhKhkoBiIC49FUn/00c5TiZiYf3ee6boOOvVTvB4cvb
1DbNuKCkxTvcZokuzbALmohx4bChHRH27PvfQS1wunjXRMXVWl70QrsU5KSL9j2f/RxAXFwwEvCD
QEJ55OYn1rQbFm3FutNbCtRpyuDMMWQX6XRTxAuP6qL3iQMZseRfAN/+wy0KZjsYTdrt7aeKDgew
be+GzTYt+rocjO0ZpCwLYj8okTOMuw+FLHqhYPtCautOXtW9rRiBPNSjfq+6TWOnSuGpSaapnS2b
6XR8HRPsREJEZnW58/Zrj7qJ6PaTyB7eR0Zt9OrbMYDjsSEoQ+8NebnpE6q0snEoKU1JK3pqncak
8zLLk/IYG6iFkhOibKQlgzDPbTIhSP2agzDCTuhVN35b5tcp9BBDsur9J4QNL6z8hirxd7teZ1/j
F/t/dfEq/uMsTD4v8XOp20REq107j5oNvFS+ENYcpo1J6IhCrhsFzFKRK1HLbkn2d+akO9tkZ6Tu
3Z6UzPXQph10pPRMWMt/hKz6XNu2emYdkUR0UQnW88FGyDxanMYPgUYz8cbpLwEDfgvF89US7rv5
ljLvJtw1rPXOo6Wquw1PN2ibiJwKTqRCdZbbjqTTg9LdJ8uUSsY61GvGPNKqj7gq9KZYXJj9XcFp
BFYQ+nKml7I7rjZexRKegWar/zd5IX0oAWo07/TdBwgX4DhT1oISDs1YFGfDmgbXuPgrZFc1QUC7
DlEQ72yOhS6E5K7FOeaSaDhXNbzJVrbkz/vAszKeDsXd4pSp9/jCyiwZrGrtkDKhdaod7y4wJB5Y
pqTYYt02BKuIPBqqrmKuS22wMzNVw75g1bcnqd8of2N5RvmoyZRBTfPc2y+QmjeVThmN87LVY1ju
0P3a4ltxAga/c34iU3usoeleJOEEhcz7ZK8d1242F8jLSejk5r5q2XxOfuGwBGS/IWkzsEaWafDf
K/utTGcZCqr4AKYar953g6ejHvLb4kiHabgTP1alfHsFJHHVI0RRCB59/vtm3+WKNenLiW8IxGZK
JLKwRxX1mgUW8usialOXHFPfEiYBDhReAuK+njZSzetaLj+Qm1wzixjpQY7lCjC7v21pqstkA/lo
jkyRDBvvm5iVxhzO/CubC0Tf+EpMRaBXx33bN2ledP2QNGVX8BuY6n/YPQAujVernfRgS/zWOg56
/73NV5B+5CJVk6P+D81kYUCUsZKrRfImY1g0b7bq05m86RR6hHTuGD6VO4fuLcrETBPccF+w4ME1
VL5UNNXXPVhqURvn55GFtwS/dix+Bp9dMInBK+ZDUiFy2VUzmJiM1oICTw/E7v3V5m6ieKB6Jj8h
skF2S4SGF06nsPakyO7S+9mkmYXlBUfZh5Kz/rxL4H1mBX8pZcU8MVSgI1DYIyU8/ksDWUBnMTnk
cNpApYES2W9uP7Lleo9werYXB3RFihZXBDlP8swdS8/qLCsemhYeid46gOlYXubywNRKM+TLhcgW
axsv28aV++wggb8R5FU1jX5NjrszauFmaOPhA2JzMXn7WcuJHxinnl1bdePnYur3789sBbaImYih
5DdfPenaFKaK3SgJCvd+h/uKzMhfa1ZF6+0Lg3siXYr2OYK4FNCCc0g9TSZWjUAAYh99T5SPVxBm
J9LrPeRldYyKPY9yzxOpEkXx1d4jJtXtLeomyjLM/IQdXZ2aDGRxfOX2Kh5XBJ3uo40MZUIK/21O
s/ho71u+Uzyb+OXsRfQPH2Kmnnd79qoMNNPdo/G3UWRdMp0lNGgejnCCt4WOjHpoZxQXqHvhgKp+
TKcrcg4tzHIr5jbv9iBbvDgw3At79Waczr1Xz5m1k7PZ0GEGDRv901ujP95o4Lq4P62q8V6jf/AM
aKuTSWjVXpFm+bJJs1Mu0224uNyWc+ls50d77feW45AjdEj+RQ7jtciqzl+ULc/BIeo6asql6Jng
908Vd5uNOozarlduXpKVqGzEzxMvskas5dVjAVFrPgQjuUusO6YxcJCHYDqyI7qRXJWf7i8Br08T
xtpzcLi/dtbWZMjITum0x/cM6zNCzvhGgLvdxM/fKhHFEu69RY/PRQT4A6nksjrPytxD3Jm4DJH0
oamn30Bij7hKedOiQcu3Ws5SLDqFgZTnsV/7W8hIwQqqOputpdUngI91b/JX2VN5f8BmVx7nTmEM
9yekicAoypxtYGHOGE/kRt8MtxMIm97bQBD/ehBd3SVapDR2iHR0ANABcoP/jCNRcW2T15jvopP2
JipASe5GKeIbSviA7gKW7W2lTta49yX3qniMZUpOwaWFL83d3n0w6ozoGWCXmgviN1dTi0CO2+XK
h3UWrUDr/Dn0rt1e+OYMWmUF4WBXFY7/hGALNvKLCNp226WJZA9SRJgKyVSwlPXEFoGsRLFVfBQg
G7L3QcU7ZaEs8txQpaYskxPhVdwVLbfqiRZtX7DWNHQjz21CRCkgk1WCf0jwlm1WRZQpZl0xI1As
GZCfST3Zf7vTC41HRmrgNYViKroSLCXHxCOvGJG7cA8pzgt2pYn4B/Z5TE8DnBZcFJpCKRj+9ehx
6OB78xxuKf7WDbuOr1d8V9aYyvu0p2h0goqTBVmOSa/fwltsmAfz6Gb6kwS0LAdNSLbF32DqX6At
TpRQO+ZWhPupLCIf1IFpIlqzIPVili7q+jQ+3BGwvyaW/vtK85c6c8u+C29q8AxlDt45jaFI20aB
x0V4gLh3cv4c8kyy6SIexsS0o48W6KYrqE/rIdkiNj67lQAElIWv6LRNGmRWFNDYXdypg9b6gZFx
Wp/RTVYquQb+K27CcrXn2CmjP5+9a2Xm3aijCYTrcHFyX33EqbNrc5tFRn5eXAi0BhC3b7xAYRZq
fFTQyglwSnDDmir6ozYGzgqQET7tiuHvJDr+Q1ywozJM5o4hc02d+I7n/OvS9ZZ9P/qoszu/V1xB
cqYE1SbHU1xU2ertmoE6WSJ/h9HONoIR5me+AEs/UNdACSWE/RfWNxvNS5BqZaMk5EuHSqxEWTjA
axaOHFs/UfR/5NfGez5TfDoMSun0vW78tPDsnNhboIKgijeu80fBSzoAqBkF0qfymHdI0wtPaIW+
VPHHb2nd3uNyiJxhR8+wvgIyLb8pV/mhHooKJDvgrgm+JeFjvo0FtAWwtr+19rzGJ/gw7fFgyF3b
CmQ08Hnf+juHsZ3wvvr9nsD74WgdAkW/BPMJf1wYrk8VjXAk8PUu9EccRn+YfXINCA6ROVib4rRm
TeGGBEHLv6jPJAlF+XiQhElmquwU0T89xFdjCD+bjenTxdNJhd6JWtiK24PVVioZOxm/bQYOeejR
1gUvjzLPxD9P+6yeIymwoJmEW0eyRU2FKeRKh0kM9kGy5mf5caKtEVUan86YxTer06kl8cWZYQ5u
kvgm763adzTSh6pgooSIS4EedZARpS3qMZO9xCwc/MAE7cA482JexAR1dq0uIbb5HilaTeITCyU0
+lBqpoVMyKrsmuKFtnQIzJrs1hi6yYQ0AFdFBI9KnF8l7FNpqhJi2TUyGeKI8RyWLcTp8C+NwUVu
GLA/79T42y0PG+9BCUsIsnwP6nMejwWxTlpDf+Rr55R0FI/+uYjtPmAE3wmOt/8Cw+YtY3FKAkjI
DINCOsDfwTgwrTC7Elv/7ytssS+MV+HzcrvSBXg50YHS20qAnDXMFbMPTI1DokxUH74CZXiWv0cP
O/7HZJn43E8B8ddvvA24vXQERM6RRPezYZsoiYDxVO/63CKH3SkF+BRrEwfrhGQUgANFYzqZqS1H
MHysTPZn1OY854UquoPN8DvDgFx49PW5ZR3PGnLer2kupk3iX81tupYwXCmbYWcZ9HBfKBLK+zMh
VESb9Bp+dp3/Pb+dglBu3yZQIbdBVRSFnzYZt7A0nfO67qF/IiIfUBO0HtiOTZDEc1+Tg/6Vkvka
m2k+yxOy/VONTpn+GtJaNzpfZQGX8k/Fxt3VW7hN9C+iCLfbBfGW2HFPxiBgDW1LQ5bADfDuH+P7
FzYM9FTFvtrT1SKh0bj2bKlEZchhVr1eFdNlTRq/cTSnK6F7My5KM2i7S77fbrDoa3csFQmctXmp
MSy2n7HJXZXgkMpQGlikOxwDMoJ+WG4LXrmBytXD5sa7dzLMawRRi0Wpof4BtDZLWEYeNsOaa5T1
SCb31SB9u7mKjo0JPAvJN4g6OIBxdRfhGO/ChjJLd0aQfHLexhoNzvPAF9SE1I9CnWUo53wHJevU
XC8VrCA+lbAcIyIcn7/x/tYzIKuuf796OhGWWzF++SyupsBQ1k8bPrz2hFNAbdjdbklR+UHueZiN
VMYU+6yWlokdb8AQZSQRGSXlfPpSCZDtaN01UgRnpMuyHGKZH+3wci5VlgKpRSMXSVe27V+V/+64
mupuAmTMMIaEzAeglLIPrx4kw5BxeRrFF4+iGvO8y47WywdPLeBmlyHJ30WUALjwBDJ15kLrzkrf
HvMLxwibeVF1V3rd6MMqSao5hVJ/8IWxr61Z6X2Zlksn+v63eLyoZBvK7qkSfx3UeiNie8fYzrPe
nSB4u4mwwsZjkKYFENV4UQyAXaptf+efLIyHNYxdO6AmKWoRpUgNyfhVrV3z4M9v7eZClqHVbp1m
OSHJpbyJS259bhj6D9RXNI0WPL8TLqfGzhY1w+oflWYYvMgciz/WRnzNkk40/8u1MU74vQYsH5wc
0nW+XLo6GtdYzJ+SGiw9Dz7yPUlu3tCJAwPIjTMOFj6t/BysFLmXV2eWwIHXx+2jY9y8HsvfFi6a
91yD7Ig9LSg6DnrrKOMTrWKbX2zVymv7nUtqc0OCDpUIKX2r93k9Dno87kcMcFj4N8d7zlDXN4lV
pupuKgs60bLj6WgxOL517cq/jddRE7C3vi4BjhKm6N5kgOIOq5S9VK5IFxV8dIoQ5SObxxjGPS4x
8UeZbHtA4LpVqDLVrchOKmW1OQmegL0PELFKKDwH6+fBNt8h0bSCBMRoKcp647eVJu3rfZDSo9xr
xe9FdfwqyPFMiV4HDXomRbvJGv6QrZRqr5pUDQ0CHuSCo7B+v9zaTnxPP5GCVzI//cPgfrd7Ejis
QbJ6gh7Davv4qsDvHehaQlu3Xd2LCJ7kPBNSTAGB8swBjyZbhJpUKqzn5bdq8sWRww+ThVM5UCc4
2CzhGCFtUF2lzFlTTIRXbMxzAI9IRFpmueuIniQUoIw4NlJuDk94JoHGy0t/FW1S0rGkNlJOqwTk
t7NGsskSc5Em+tpINcMt3nGqXvriCq3vR+6utLn1zkYBPye3VYYKkUOryWusUnBBxZ/kYej4LiHE
B4yhAnKQytVvLZ112OoTYZ3tLbTJbW9/V/OWlw4f/yBAevr0293gteVPeg1LGRMEuIGJIWkFoYqA
n9HzNEK15/xPk7oGozHylUvpBMe7Q3z6X4X/jJrcevCLkjr6+5IL4dWzwZgEZ8xpBbvfJza2N2Gh
BU3+0l//XtZvpG0UgUrGd2ZHSi1tTJXppbbeQZIznMEvlt7Up7pnkVBgltd2zIqDAO46gV7QSEao
AQWSuWAW72tnTLUp7YxcWb7vDhebHzYcrmQjEd9XTVBwUo5SvpY9DD8Z6FPA8mCvLxhgOl2/GSLc
8gj32UWRbCEZSEGRY1k2eUEX56NAQIPT2xwm2OOG0Nc1M1burnJe+W0YThTBdZooa6Vdtt/1+Czw
kCYf/HNxfmONa5Y1Sh0QEklrq6ai/wDH3v0XenfPWF0rT8KNFxC05DelMpolmLSzQ0NqwfOvaYaf
ThmfDlbXxzZPQTt13YDpa1wblWfJad7SWVRxQDB/n4ciRQ91tsEXNNqDp/P6wt8qolEAhutg/cBR
c5mURjcam0YE/gxkMo35OzEdADsXVXxKz8HRG6HkG7tWxfY2B13a5mlCN7rkKfEmu7X2WgPVS5qA
I5XEFBlYajPFBPvW7eoTHx7u1MY7hV92C3K7e0jq/6FSvrVCfvHME+GGcYWrw0SBSr/n8THFrqFj
EexAQ7CmtL+JKEdSXOmO9vewWgDRchCgWYD84Kf48DMiYWOS2A5pfRmeY+gMB4KxMGqRNVOWq8Fm
/6LLKvpbjQcE+q8tlk/OtroaP5K2i/FG9Yywtcb3ZLQjXy+PJtiCWXsimhWio80DuBlMI5ORa2bk
/s9Y8zEAgI1PAzSShmb5JQleaT0ZRaN3B/QgEI1DU0OFZlhLx6Du00dGELJDUoK8sJg99dNMp6ut
zYNlSnN0GXh7B62Gf81ftsIL3gIZF3qRhdpWLNOkPvxNqRwGhf+BtDz8yR6iea4OK4It7McNyX7n
aVJZ1MT/0aE2/8DcsSWE3wID/O1BEXk8lkUcykk6t4LLx729OIwvAR/75XunT0vlhkFuKcAKVdo/
rooDpNb/XtxMAeUY9T5Vb6JDLJC0QqMSq0Asz7M0G7CeBrzCWP4ezql6/URzPiHVOtiHPMAn+jP9
B4o3SA2mthU2gYvDan8UcpuVxRNVTY4cfrpEtM9VJj0ODaO0HqCI4VG1LHibJongF00/cgdl/jOk
a6cb71cUyQoQFcaZc1wOJANcZhJ02ORi+ITUMtmNAl5BB4+vf+OGHcfCCRYRvx3ZIsRLTkRsYWR/
vZ9g0/Wy22vMDoSLR2vtpHAO4hYt8DLy5TIiJ9TKnOrfILD+e2OsNyAuxUIb860g+ZhjZURBpYc6
6y6vZ6CQiKMZO++RllTDDb+0/lH8Cp8XhQBruMmbFMGztp7j3jRnx/t8ah/JPvnhwH5OTOjOgU7l
0ZT+PjuXhhsqaUO0/nLQ2M0xdxsEROfUU7WMNqT2kMrFPKIgirLwLVvdfWvi44zhdoIA4l4Amgco
bQtFdvJMLrQqUTIqyPUSskSNH//v6aWi6Z5pNb0qbHEVjCi5d2jAXxzkMHZVwqRZGdcIMmpYQTp6
SY0wdkYbOABc7ItNDsNPxMn4vIaVqgZ6njNUqPBLeyeIbVW8b0XcwFUkAr8GPg1gmBdA+2jf3w6P
z6VMcJnyJSC0+2PKvaAj4UDVZB85TTK01Q7ibeO6hlA9fZeHiEMBU/Gze0nRd11F310IasdyI5zC
u3lbHQSyVyzpTKsQlL7gcsNK2RPXgfgxzJzs2ncMRprpUuF+Qk5hui1DEx6UjhgsScVg4O2riBPW
zPDZHaqpT6VTUQPWX7mTQjtf9NTFQL+P1ZYVnYX4ZuASNPBUvtVzL2BHfzQmbE+UXv+YN7cO9q/1
x2lu6YKiNav5g/8Ebwwm9nehhx/jg4wXB6QyEha5oB2yZC2Z5GEE0581k9TAM7m6zK2YtfhZo+5L
kAlFInXkK4Jj2A9Gk8JwLJsUoP6U9RbVnTsIho1AMjqrkZU1gueeZOF+3fL3v2oq9wSKa9GCORza
gmXfSqujSsFME49EA2zmPYNQ+SdXbkSef7VXOckN0uSdM6mZvEL8qvtrVe9kwqgKGw59lg23eMUZ
mcgAJErCyviX3/CNQUfWDUWpWcSkbT8P+zc2lnmSCvf6Wo/cvoXQ+aBe7Zvz9526ovy/7gzPL2yS
dnwxfs2EBm75TfVHuHkTmih+klqWSWFrjuYarlOalkEN4BNsZRU0Kd7w3sZ7W0VI7PB3tV72KbvP
aWWfHWbb1HhhbpqRU5UiApPzHPbhLBcL8ZUP0QpHEvC1ljYNLYvt0NpTL8M8J9f1UrbMquqEocVc
IamwaSRhGlPf7JzC+vOm+YpebICQ0gDzjhuP4b+FJSBExxw2O0JhF4Ohq6F4bhkz/jGWIc8XdKzI
l0HE1Vrywhr5YvbUo+RCmPChEctWWFDDO1yKXRm2iMLaBiOF9a1iFavVInZEap/jqpIIP3QOTu4V
12qUGzOp92ieOypmSYPLic9Pr8LijN2qC3bv0lklhFJ825YLv3I+cqfNTXd3XsYlmW3KM8McRKbo
0odTRZqm5Lncefmm+C/yImiW2mKaXOpQY48kHuWfOipa9op7aNsBt4xkjcbPECQRgPY/ShB0C+1v
z6gjGY+HSudfM8Q9l1KIoHJkTzGGp11vyxxwNnEPkCbbokCdbRUICxWrHv/52Qj17kXzYRcu9ONt
LI9UsBG7hnazhRtc+29khYFtkJMObW2bMwLEesCty2WZaqOfWEIz5Yq1z9ho6AYJz4xfVXPBtlSS
4dePwy/P9bIXse6c/nMfSdxLlTioLNEcYEztAEwkW2ZYcHzpd5tzbCdGGzUC4jcLlRSldT9agaaj
/TnROHG87IirzSmAr3vuXeF4C/y5Kf8nGdvTQ+tsmvMmLmZRA2m4uviRYA6br5EizV4gQA7gpdVi
qzgdHTf8lCwrV4lQf9fpDIyhHeJqZiiJWuWYVeOXvhz0f3p8A2AXaV7c9HBqBoQ5OGz07V29VMXc
6fZKPLjh6PZsDXC2UXYIcmGiTgHOQNTmHRfMdBBlA2b+ZBdb/H/xHSamuxAUgkqA4vd2YmxTEp2O
+vgozMhA0wBmCycD/rH9nilxVuxnBc39Opm5lRB5NF2rl05XhyXj/pFAygsnk28gq5MpZchfMWR3
V0uLquF2OvW7OyXzqYQMS6LpVj09TMkJk2n07lhKPpxnwaTEQdh+Q1Q7+Kj1cG+RC2+pXXd1F2gZ
BirqlTBg1bjgo9nXQwm4lskRcXuwPnGBy4UqzdyNhvUSwRh8m3R710nboYa/eZX2MI6YtEPmKYrq
TCoVKYyQQehalYwqptK/quF+Dd+wW1EcKHVUfcrIKphAtzzXMX6VqnySgb3YeuBIVZfyT7POTYkT
NkT4Q4Gyb5YQe8zrc+GQwso++NSCcQrqwrKIH/oJ/GaIHMJoWI5z7fyuXxqdpiknnSKCCKikVwQK
4LAxM8EqsXsi+07m0gE1sVz1qoJ+5X+RMQe4E0drPkQYtohLNcJ/cDeFigzMfFbWJ9OJHM7tokCu
mGSgEcC7uDtp1HC3VS+39WH1qucfdpXUlbn5Q3at5/cQ4hLYvKZVCE1VQxrUkGpF6h8Off1rT0pd
eFioKJ2BE8WpoWuFXtFZT7fT5H/2H1Y+99yqKSpqLQ3S33N0aoey8z/Lpd7PwZFiEuYhNE5ngUGt
RyXNSWeWCs/ikdJO5/GGJBKLkY2IQi01kxcI7+Z5m4TnMNaVnFLQMCP2QkdXAe7MBPH+BTan2hl5
eTigKFUX5p0Fe/SGfuEShcxKQU8nJZBj3p92fe9FNJH1WP36Rg51ZlFK8x5EnwsPyueaoePW1Okl
LSJgPxejQq0nkzOOaYcIJoyaGOtNsuvyPTr985I4L2HuNogQ4fm+YNfSVKvtGouAYJplBBsnYm4l
8MD5VE+jAzS9rlzSLQNwRqo2wWS15J28DzzJ1QAaMl3bZvmtam6XXDM6KkBs3iPZklbsKJDfh+lE
qcZh4MBnmDMDKVfAWX9G5mvakENNmqQjQOwd6SBrpNKTlHSqUg0PSiqL78MpSTnHjGTSk4iJMNf9
i+VFDs2fiLrNvVsxgcwmHy0PXWZh0HCjboj5Gsaz1/FTWiqLYXSkAxQDHCI3E2v4G+/XUFynZwyE
iWoyNFDgtlQHX13FZLIpc5zZXBhN+Nylw+o9cALjDcbpDeT56in3SEtVKRL6GG5rQnzrC7LTtyCF
e3e7Ze/QHcllj1ljD3tDegru1ZQkWI4l8I4rhyc3CRRO2yW/uN1xkwl8IJPV0BA6D8fecQc2o8LR
JFwrdrzN4b/Y8vkFkRSz9JJcxsBbz4YlpH0MVh6+yCO83yO5+5Soy0v/AopSasfWvLmbI4IH6jAi
r/nyKi4xVUBRJcOaTBiYo8/Izv4EmxVtbqyLYeIJ1KIs0n0jfmu0rJvly4dRD6kh5nKqCXNaQ+GR
/87Gpi2Pg08Tqvocm+AQWz+SD4rGOM0fv4inHsBa/fdGmTQATMlUNBE84PvJzFY9k72B8ztiENQB
MdCgmbvVDUWELPjbAS/Bs8J02pm6Gd9u1NZES8zhgiCG9jPZcpyZ2uj9WCGD5fPAWUr7TakQ667I
jlBxMKBiZDC/fR2K+y1ox3mKixeEI0fS7EWSzPLdF0PJHEWG6FPOy4tathjm2XH5Y/ZCLXXK4U4Q
Ehr0v82dx4f+XHceMIANtjjHy8HcOYX5S3vQq1cOtCkV+1zyMopzx8Ply8ouOO26NS+JmtOEpozI
I2Vwoun3Njul+Ls69bdm+9iMVRYgealZIkTpOtdf/Y1G53gcrp35nNIeMkNQfWsQmxaxkR8Ah17L
wC/qkTGc/kiPFY5b9XIYrYzI8OMMe69xZrCrRH0NZ0Vj3C9p0Y1WcOCLQTn4V92m2mrneMh/oLAU
fi3Mhzab1WKOnKFaRp7zu/dp/fajmMXxZgGYYk3xhkMvdPNHvQyf3jXwzbUX89LSivRu3fkW5BRY
GCqVfWdkXSruPRdFHRpvomZZN2FlOgx/6551faBZ0NIvsAWDMnc0iABHo+AbPBC4FT/+vMK9so3G
GSf0Fth0EbbpqF7CQFveqjQ9Xv0bSuzVhEjf3cVlx0cYuxlPiy7biVK9kJnbs7GtWd6ncigbxXYH
OxO9nhTumIgtH0XXMxpWU24xVnb4qpVOuBuUmDs3fHofY0vYuYtrmgfK2lwWSmVQEDxjrkyJxgAb
PaeRl5GJJ+zvLWqMC4nV0aK/73cNKB0VGd1wVTxvskEKefVL+WhPvTRKz+CdWzdq7XGWdZlFPji/
tuL2ZEcSa+S0tR6j/uinmoltfcKwE5kq/nw0DwBXJxL3m4xahL6Z2QONoZ8prqYfxky3spLJpGe1
DhaLQxSh0fkfZaDPrN4cpzzyEhfG8xzmwebprr0FjFRFiQqcLGqxel0dk3uV18aY//XrBl8Q3tju
cX05/Qupz0MMU3O9w3QeR/KBrhno6exyCT0LC2zeNKWTQRjrinO7ps6hHucTT3fiI08X/lR1lhMU
1q5yOtuKYjo7YtBW5o3Xv0ifSH1k+NSrozRykriVKttK23x0IOHQMlEfH/u4PAlsFw/1dLJ0UhNr
B9l2nFCzyHGhn5DdQ0pDVgfQffeSB03HrJJCehdSWZC5Pl1jBWMyiUfJhcl7fdmfen79P532mJ2d
ARSr0YttnS+1ctu/nhE5b2yJIujyd6LmI+qJX5tmJrJq91HvuOOntNLG6bbUGSusuUR0JcsW88sY
XesugCkNstR1TFI8+fLNqYmOf+lIpXaND6I0k+WlGTKF1PSaJad4hEFhVLqf0OwU/S9jWo9Ojf9K
Tl1IuyJ/fB7aQBJbOU+TG6FiF8jywwomc0VHqHIz0jXtT++exDVv6Ftx7AK5EGGnFYKGGRlMM/cH
KstsTb3k13oSAAhVdYYfz5fIuRQeTS4cLFNTy5FIGc7Heg+Hb+6CIqemuCU9vnJxJZjFjAn/G4IM
roSOGASecI0zV5rrQxMKY4o57CEV3nDxTCP+18a4oaApNfiznXAwMsLz5TJ4SrFtOMPX9p9PFHgr
pbrXRCDCSnJgd/0MPQ9T5M8/1Bst+jqUu+aY7zX/dmACP33cycDMlN6DQReI5kJkNAucHSAraPcU
/DO8vK+Gw4cyjCm8WLUn99xpzDzLkq6ILgcE7gRT3yQUf49KQk3Ev3BP23dz5HWCHBHFvoAtuQt2
iIVSVcVQtLbUhqnmuWkzMDKlU86GejGtMMBnAGUqjzPN1WXPkrVdqUUzJ6RfiHLP33o1mg48KFkU
Zs3b8FZudy/+LUu7CvMn+RmlWz62+0BQxhomtlf0z6+WRZlfHwFoL2T5ltBmrYo/At/xxTk0cEOg
1zhP98r7Vwo7fKPxebvuqo/H3x4D8bu0KZk97IdQB/Vlr+S6xRM/gDrsh8L7IaYW0Fnr/BR8Z/71
kEMwdhHZwPzFqbK8x8utkgxra8fTQgzgpmied6eLjGDIcjphsje/BLMrwSXDhTqIYhkJ0barZRRg
a11vbNweHl58rdOAMNC7SDRj3tJZ1NGEVYk7Gmxrgxo73MtT//S+cUXVu2cTCwdPnflUfHj92qb5
DTReNcccCRNBJHd1VPVNFosdZJsegLD2CzCI3ihJ36HusRTnQxmtzA5uPnWofIftwDLa/0L0seTA
iIA7BTkWPLt6ntJER5aTFmM/E0FUkdzNOq7umG3Zewhq3chQIQjEK/HKGFLSIfduBGRRo98T94MW
sJlZGFnMUt69FoIR2cv8NJtT38WnMaW4CROFUzM3qSCYSIOi+7NF+0WV92BxB62Nh+7T7n9n/bbK
w+Gah/O0/4DXWViYRuTwHTd4owFV4DfaMScZoE4BtxFHRFRQpDYyDrLS5PEwqOCpVtvxPWg4SlJ1
bx8+bVBojEJQWGDWaK+aQ0Tw3mJCNLn7blHEqb7xoeAx33spD1cec7NnUpWf/uScE5J3MmgfF1ls
qzbiXDLsPJKwQrUmCEgPCht+XqvCT+oAXY8MvGDGAmwu6qovOgQJ5etBe7O/dqreCcPt7sR7V41Y
od91+7MRXyQAlezRwxPnpoPTcPszqht0byvLlZDqUtJX5Ceq5U7qZYYcSih45+vA5Hr1c5azafOR
Df0aHGBojeQI8HlAn0NsbhlHGhd1yLVphFp6BWkSsFMZvF+wFeIcUzBgYjtPA89tVkzSDrcJEfdh
gixeQkZ4iE6I8PO85CWcNdxsiqqrn0zkglFHInRcMUXOtrq4vPidrTB0+yN1M4Q9MrRonbIwxmGw
CjcRhpPLynO21kx7XuBG+/j0/hLHL+Iyn3TQbbYear0vkvrrMifvEL459kmc2ilMMprju02Ve7QP
G2Buq3L77JLgYX/CDX4Un4vY/+i+YteJ49ZiM93xsruLt2ddlqRayU9Lgel6argI450g3A6Lm7vS
yfacFEmqBZKwpVDqIc4FQKE7VC8L7valfaq44AOFttQsg9F3QFYzvMq1S4gh8qimHPG1TWa6ktYc
cTOuTiMabdmpD2wLueM3JuOvLeKQ/zyE7XoaT5855qx8VQMYmNS5Qv+EquPUil8njw7Ik5OtKLOC
qiSEh+epamWjwz++NJFVTe02AyDD6n70F47HS47Ru8kN8CpXUeixPUbfgiPXXqtL4BkJuLMJrp6k
FN2RkDvtGPM+rIWmYqLooRP/m+pD4F2r2b38TSmhxZ+nBzWDqj6z76MfP4CJrQxzxEVVApb3jqwL
ajJa0RTzWCJ6pEsQe1g/+gBVQTr5FIkMLRENAVJZ3N4CH9J0lgi5f+aYtQAFR7GiapSKBaXb7Ui/
tEhZuj9NdLQ5YK/VItoLPcJ7d/LcJbBTyjaLUxO12KdccBTdiGBBpeZ+PAdJR0zkZBNgq9V7E+t/
h8Eax/2rXho4mUFcSrOLrnjUAchxlZzrKiOJz3qBn+KW+JU3piWvLagmIpjPtmy6tzYilzlkLd0F
kr0bLkO3VCXzGf46TNEzsSScPNOuePtmGqg4m0pY9AF3S5PKiWTOTkjgYHJYOkKSsRnNCGudcjFd
7j4djxijGVFvYdsrULNyNjXquVMOv7MeAx9W9SFUO5oTHQmK5BmSfwTDrWF3CopIYuo7Fnq71Kba
M49l2nvuD1gg4/QBN4YVw8iHsn5dAzzbozudjPO8gV3smkD/Wcvlc/WAJCY7sAFc51mkvloYiBt4
4aMYs/4jbUfH/A6Us5W7lXPRynUsulxWyGp9sGZEGdwixyy7LZAmNpdEXi2rcOtf0CG5dJIX/kgY
ttW+K/AD1v+0c/jaWudkU8D193+YHLlZd5CUri0g/BjBedRpmjSWOM0rC2MIxx2DwuhGLz6dQ6hn
ugJcn6ZSlK5FgKUCUXPdi5ypH7izpD6aizcBExMT67u1tSP3LtnJLMRpumBM2sQ7ivqr7zeIVED1
Y5F78qmeqNG0jHA8FGyMFOYUv+tWy66fNbPK8LIgMSTzzDzaBFok5bVHVh7mTLzdbu/J1RtA+xhq
sLTtGKIf68B7HJNBpB8EBohgf9kqF+MWBr8eXlCp1pgQcp/8PjKpGGbpRwYtwPGDJUIL3LkFUzAk
6QR4JkGieQhx2ZtuSei35f5lFp5Zc2g/IDFG46kA9FuXy6u0M94IWuGZCsyXnFbYDEHKFVbYTn8Q
A56jYaQXELL+jMWK3NQsOq5B5RLer72ogq6f3y0fgNYkdWzF8cIh5/rdmflYzgZEPYfgmMqo7bn3
KfKKdXiOfnAkfuInhAO8TDOzjlfIhgvNz4zM61qdgPc8ipEKbBriKBxRgle+BAVQgoLM6WPaKiLA
TKmXMoJO0gLUCvzdMPJPwRjDxN+DS0o7fT6zwGrxYXmYBWf5FiFzTGHFG3suRg5jIcxUmiAQiEdK
1AcIRnCGLtxuhyUQG0HNkjrAZRj/xEspcv/5eGO6yu1xSM+taoHvQjHJZC+5CCVJ9ofIqT1dmOob
C9JeXvj3tYwI+AHdxSvsikTqhOC30eqkd8nyv5lvaRuxER8udwduFteqbv6Nz33o7bsfwRRTmtbX
FTauGIl+375jYEbzdATYnszpZyppUMfJLzmqZXd7QPS0dVAiK1I/etkmkPCSLbXuk8A06Ih44teA
ivS4cGsz6zLMsBgvVPBnOWi6oor+yYjylU3y/5MN69T3Bdu3PktWvPTbozkhaIcMCRESRBBO8c6A
qqnLC2F9VJAb7SXoZ5Lczx84NfYugMSt/5j3kJXVdvipSKFS0a+/gqtMJvewNtHHKkYhjMkKvnKp
5HUYiOl3Pp1ledwYFoK5I5g5VxalIOXWRFHm3G9nPyUIBGJeFZ9bePH6D1qjf3BkMzu6klNxuToK
SFYCP2DKgI21AvrX94FOKxb/iNB3iDI2DL/CUTteaj+wynCPSz33B8ZlAGruV76nk5NltSQ5icX7
TmQ/mLkF/pv/iPq4zWSDQBF2GvicUi8riymiM6ZQYiPQVodrZxH6tloiw9NMq13wMo3CZwRRXhpc
nomsXV96FQ0kGeNGPavQfuZJ1rKRVAClffWBWtysY573PcRs7kB4DDnObOTYnlkLLsKspB8/qtNr
15d+y/vxUED37nHh6pdTMBd4T2XUIG1RCf0G7t7gGvlVuGp0vh3dpX2fP6/F3tqGMpmIMQVi04ki
dObhEQVZQTnaQN4/aXMb+y+Wou79jZXdv/B7CECl3kaCYvOzbVU3vUEYktpIa0a0JTBWr4IdBzEx
YJvtgs9zypNJOCzq8mPZuWWGjuCKWKRUEwTny0y6MB9LedhFAWAd/p/l1cM7zJVQhk9gJU8i4qH4
Em3mAV/31KwlVm/wPfenbw5uEAl0kneR0AxNQy2vvarbAWhXp39mmXO/vcpP1baYh8Md1ISqOpJz
mIp6YW8InKE8I6NWlzX1ZzT9T+n/AkhPZDFa/6a/NqqwYm0gn1h49DAloUE9hhwqxGLjmwDTWcTi
+w+TbPIPY7n5s14RfPUf3Qp4t2Lo0hFB7Q75W4AzJzzqDJR0ao+BAa1RcNSiyBncuJdvk7K+x7Ct
/mWY7OY8iOk2cnH5Zq+4DHVac202P2cXrDlNMC2WnxPu+epK3HRfgGfAs6ZD6ApzX6ktdpDnOp3A
A/wX8DJrxr4K/rLrZKE7vtHrAS8cdbK7l+FBKvbPQwUYB/YHPPls56ttrv9UvEHBFcIXl75TTP4y
iuaxiEAfScBicZV72Pqa/ektsldBTXG7OS/VBftX0lIO6LthqnRqm07HcBGBo/C5PP8YO3Fuh9DA
I1FyUHpyperdbE0PFmXmdzpUe0RZ7V7C7YOOcGrmOSL9q+QUiLxvnl0/qc892JNj9NXiBucjXh3S
KzMT+YmwCvl8bir+upwS2qXu9YHeyFyNZZgHtxQerg1/edWqGVLPyZY3PSgtlv17F6C/82OvqIWP
W8NVFbn2CGzY6QL18AlZ2KToPv2Xx6echP6efFQWsSLgnhu0j+lHuTWzRlLxwOwGcvGKe/WfAP7T
5BVnpi4QfVF+Dzke33GeTm6zqznofUN5JqVJvxWbpaAl1OCwhNh0XzDQBVu1uNivj4NFAFc5owj7
aGw01mnEpGoaOpHL74rzwGR6vU1HnS9/z/iLuY+PCs2SZY0sdExFFQAGp7aQdY5jWkG3JrsMmcra
QpJConFdYL+RlqQVAY/a7ZmZgOWU2li+zxsI7/UzlM53GjU4+5uD6UfKbjMQgLj6YES9oLI3D2S5
RpFQmg21jEQgUzVEjMH8MEaBd0ps+p6D6OrYXNoPhGoaEnIaq5/fhvLDzPq6bRn8SVB7w81LN8x8
Hh8bwRlfgT6PtAuwt3QutrNGr57ndXja/qXsXm6ng13L+KDhi2VmrYViRRhnSLSDQoEr7k5poz/d
IyM3puHi6dsEF47IQvh1fvs7p1khYgiiBhrvltM5PcrTPU5D8tJF6LUsMM+cBa06qadKiQSGylHh
95tSscpkPBqlRgph8zN8xFMyeVO9advgehA6ZSh01CesR4Azp8ljRpaaud+RVz89k/spyr84OeFr
qCzAdLzMM1UNPIpLvvqRZKio6rG56ur02FEqINedVwNZP2q/hDMlTvfTAhSqNWc4sMWspQRv7VA/
+QPadcVI8vZJgOVqpDhD+PdokyxpGw/sDAAFn4vRGYxHzFlFrFlZHCAD56OMYjXAngfdO5vtWS08
+yUbJahSLn8qogJN0S0pRc4k0+cGvCssiAzmjhB3N7S/f2Z9AB3VQE9KMyNYRLa906PJrpXssriV
CzZtDNFVzniM+8UKQRbCZO+i3C8eLhD+/cgyL4mD8egU6PShpwsCPsuzUgXMmWeiIoMJlPPAiG1Z
A3MGOiC4tY8WCcH+6vumnx6Hqg9XTs9WAubS8zChWC2LEQJHonA6E9DdYJbcqvlYDMgozE7loCeV
TQWerLFPuNEuopVjORKl/diRdec/t8J08TC/w6Qxgyyz787r5210pd7FRPJ87CkRoRHkQYSgucXo
kET0CqY/2U+MaellWl90q3KTe2vfANcixTHgu1tdIfYsSBjg6CIHK+1Ux6xkPACwAqzMg3xy8+T3
jkaH2IF6ZVjVgWVxwidyURqOot6kkpfKXs7uaRNKReKNo3bPMG3XvkezifU6dgi6zqRDkJvTYt6K
eXW677KtQsKTvsveImVq+Rvp04HWCwlL7YC7brNe2dRD7tUa8JTjBf0Np36n/ZbF+3mSR11qAKj0
F9DG4kRo3x0d2LoIHSlaTIQ7eQs99R6TuYEGjfCputUvgmYzPlMHYlk15aggHcaGI8l6ma3xjKvj
r4q0FLiOCj15Sh7ReMHuKs4AxQKMTO4hVZcKHlLcytzvkeV/ObKS2Wp9sKUVBUtNOxKFNzfv9cDK
lKJV1rd+N1w/IUf10B/O3Ny6Vg+zLf+r2n7cmaDFQgXuHzZz0/ITZC+cc0lTj+FscGHpE5675d9+
VPv1TXoIDmZJGYDb/EfPlDzO1AbDxb37d+ppCZjMQDHrFy0HVZ92LgxTylpSYr/FZJb5u3OGPCQY
cBCA8K5orRDDyaLnx/I29r52hL/xkjVO/59QCa0zwBMNCLvoWP0DNfmPqTv49yVxITstUbZ1TgvJ
GP79gtTsb9rp3m2LSPuMO/0/QCTG8iP6OKu/NkR37tXn7ft3KHhHr5ZRocRdZlbJn2IvGkDD9Eeh
njtHQ1Ev7Y5rFhA0ziL62nJTQre36yW7vzkICqMb68QATTpoGsjl9ajABS3Pmr2BrCa9Zk43TSXj
PJCvAe8GO0RmOuhMJ9WT0C7sZJBaSXwJ1YvtgE+kOdU1GXVGQwYyECGn+rY1KoXKs2SN0AmLoZPq
aCD/9UfjA41s5fHvkgqE8Axra/KidkJZ2JDB/Zk+Hji1SQZTm/puYQq778Oh78+/u616m6JplqUg
orAPhTdnZNHym6YmQPVD0elRDnBHnWhTupd5EMPyAwTigjclEknlZSS9tmenWm7aZlezG5FQaUKl
PQ1r/rIG1daq3YLQIonl2BEpkSYRpNFoI3HW5RRi7vKjZMPljM8NeNskT+8NrhfrAAbykYu+zhxI
8GWnrse8l5PD6avw9tWnH7CuRISHmrGD1KyJQPWNIGxFeBM8lGFOiENxIsDvOmDAi4SSUZMN1AlJ
r6Wn0TCeA3WCgIxyEHYsULs462eMUTlA+HcJIeYmKyCV4O8SkkvuFy+YueKOc8AARzd62PYkB7kU
qmFLG9h1NR+Gjxmof2BkGMGj0MwZWKCzXcMtfF2dd39xDTSNpgbjvKgEcTGNcNkmOA/avDev6m0Z
bsUk5ucGVSVrgRGryfd3ZROIjVGx65QcKGmWmHTdptD9HY3GQAl668xTRZ/OgEr4Fyezok7G4m+J
MBTPBrsqI1hHXS/RUQnViqrehKfHRqKX0l2p3IL/UvI+dTryYf3iyMg5F2yXEkqrq8b88L/4QqxE
oOk+9QVpZBc7w8BOYZ8CKKeLjLTrU4QyeW2fo4lfpiJhv6Aqdl1Ehn+ccnvuHXeQwdQCpoqVmkBQ
PrPgqvv/m6AamPsFaQeauO18+wmlg+o1bD+vKpW8dxkZLIRyxgIDryyDeYLohM+ssU0y8IPPjkX3
Bk8oeTOCoSltcaqWmIeZ3xMlwXU8dpgAfUpB5E5KRgySJsvsvyLtJqKUGSL9JURgMiGAcDHgdVdn
d6DhxT3PUXK6Y3du79L06yecOga/fReHnjbZi4V49nzP9CFKgnQyaT+5ERyfgk+MGOj+aE4EhGUG
yZWsBC1iYxZatlCfMcGNHCzae7uHnuRe/GZivvWFVkQAHIuUp7aiwidsRMuNxm6dNncFqLLoUPiW
NrvFW7vaDwfbayiqAELuFpadXnQnkR4rvWQkDbsdi9ZOGK8s8aoxeDiDCXmuKI0Bo+B2MDaO0Gus
IDBNo5CA852+j4c4Ga4ILbwSZvnWLLI6n4rpDBX+d87ByWctZD67TXNWBN/uQBjcUVFNeOaTQN/Y
6R4VaTiiQIEj9U5TtykSaBTcW3Abc+vFAeN52r7W84psTVKjeyYrklXCdpeacXuodWHkSq59pgxn
kvrYbNEWSor+KRsW6G7DniYgaf6KluXOzXlSOWGy1o35wNqqDA+5f9/cXapC0YvWdJ9UajpmboY+
1eehtXznZBlXBibzFQks7YT/xv2bnN0KNQdGjktKA/tQp1rc1VU+yLatyeiOgQSbB4e4/LnKEdLH
Q00sftLVuZrhb1juvvY+EpgIrunIQ27T8EVtQvyaG9qXqejJLUpjItXFdEiK7nMB/ChAJO0m0XKQ
lwqIuIv0+m4B4WopPSMa73MeyJLopAf+y4LgV3c32+fml2gY1q1B76r1kURBmxWIHF0U7JrVZQ+i
YwuWvtCHpcwGVCyB9HxVMbbpkJ22GotIFp6CrrmzbuCa7Kgld/lONODJVKF4CBXFlGXgXHtPbYbZ
iOOG4Stq4bHJiv0znSCCDI26MTdNJsKVnXdF/Ms9DZB1VD5Lhpg2W79P6vOH5UsdMeVkO5GsuwdQ
aaxBZi3BBkqlQ9BY/G0WzFkylZKfcEX1GZ9PorV+H1vEAmrjjze9kTfKZYNPbsm1gCiFm0n0BoQz
otR+zGfJKfMqYrkLMSDh/wNhKWDy4Kon7gAJ2zS3IR7/adaqnlgLwAGIEBc2/ODTKFkOdThlECSE
lWuVyMB4BQfgTwQXOjgQS/MsXHSN3j0nQ5LYt+3W3frezUv2oc6xIpLg0s4koNRvahrBV1R6vo8A
oWiEzcqvruQy0mKVxSHIhHLgar8UzVTzT3mt46qIDRQSOO7WJYPnkTTL8D5GnSe/89DZQnBQsGMf
i8rJWA8ff2DufJ6caIrAlNy4oqJVmhCt5B2ufanlwLZiVTztNaiUvS93GzZ8vqPOsHRjwzi+D+xA
gt/dEzVK+zYEWoPeGUEtUditfzVxXAdiytkPdQRl7sFlCTmea4+iXLx6l9RycIKFhHc+BRnHWt54
c1Zez+cmuzJDxDhwZ1iDm7zhFkxPeUTxA0tzSDtRP3EBuFqvX0JPaK7aYRqXTVDzyucAcCtUK77W
WYsYiqZE+sWdYV7boG5s+pG4dCqG+oAnYa0jN5JsMYh1hGnuaVpp1EUOWo7u/GPc/sMhQ/4xF11b
5rStIPAdM98YAaBVFSBX2chselIrZsDsQ/My0qIz4hTB2MTzPJsqU2czCV6QVCQa/UAvNqQp/Jf4
yPKVtIe51Eodr+rZ4tvb4TpcRFnJFKLd6Jz2wznHyeePOCepZLwKSI15clHqWbcCk22ySW62wnL2
pki1jsTnaLmkOmkxjQLyTisRKM7BhqkPeeTxC+7hXkx632lH+r0EPww2MgzBhnSYZrLXyXxFUjXN
V6TBbwgmVyy6cce9FxModwBHLIzrT8IZp7dY0QQfznfBQ8tqtn0Jd01IWrhvQc3s8Fu41SKIvFUN
asCQY7aZ16i/Ng4rKL+h/lLjktEVfhyjsWsQwRj2fu9YfAfsHc8fSUTX7Ny7SjJ4nWS3zt3Au5TK
TTGRtum4lJmeImtUxkIvb8lKGQBHIU6oww3OnvJO0wp46HWZPp0bJerBs9ACMM3oG8wDoO5zMPaw
Ey47gefr4vyJYQzD97kIJ7BN9AoFPL6RX1Y75p+mnXiAEOB3W+cXKH9vP4LyIYTxigVDumiZnyRE
5gNd0Vgbb9QrvzU5JOTaHBckOK4G+tGIt0VZymiDcOyKdxarJaaIyCwthcvFwM9xPclZYmrs9D/5
xqpU1bRBOEk1n90+nLKdUnqI5HNl5zgBcr26khYEVNdezsQrMA+U5c1zWCnjE9TwYKz4uWw9b4RW
+zngMPOXK+BYF0v7azPCoo2B0LqtrE5KSJN88m/sm1lv9T49JZDSaYq+sZBKSPjUjOWIz5OtEG4x
oCDtX9J6tcQEh151zVnCcljAugwitvxjQmqw2a+iSg0HeZevhyWXPtUrBQo2awS2KSAhSwVI06og
A1Z80UXaMRimnql4nl8hRrb8G+fuZclRiDLYMfFeg/bU3gecNjOoXFORVYUQ1KspZc+RLmOG5TC3
tYI9TptuuIvMSA+v7MBT5KzZFo1xlUc/6ZfIhDZxkqTvKn/dMCJHbWDTM+DqhsOVXV4RFGDx8wiw
qwMLMxHdmHNwjOcI2Q1fRLW7vg/MLbw2RfSZzuRSIyvaFSIcO59ws6GqyIHobmznNt9u9+AB+1zK
lhHSCSKAkKcgrw/VavVjnaGOUYc9VhE2x1DO2Nb7XMWAYsd7IeZndR0upfvo9YQsyfTfFNDJ4p8s
mhJtvjR37WcLHoeGCMnk3Y/W5MV6G/LV/veuLxCYMrYL9Ta3soswuGVKhUiVzWHD+lTc5Yxo6nhj
ciPyqNURFb5FzHyJLfuo7VdBz8yFA5p1Cb5rw7vQ64gZ4X6GMNSA5MODXs4BPBELbkhHRTs8m2CP
YS2ievleM6Ium6fm9DEeT6q2odDwWztNPe5qv0+rH0aLx0KGrf5POFWv/E/OFTGm4Qnt+bPNDLUk
IlByvVnEvV6KlJbxD+tHTwECjuM5CENQbmCyhIp9VxGtZ9M4fENhfyp5OXvBDA9LVjgnhEzwq3oC
Cr0FNMzieI2WgpMgEm3D3vvhZtG+lM7Bx0PE49YsfnHV6J72YYVZ7GPT8su0Kjd30iPM+yP9etxv
Nk/QToDKECJ2epruJrdo0UhSeChcRc5Zs0xQALmLa3BwGQyAq+UxKe86OHVtik8GTRarSVvJcQvo
VkRXpEGLb0NcPgl2UukGUljlBYsHrt8i5+PkW4e4RIXfrOvpW4L8KPnRxShxN7DGScjqSDmf3a7t
ynAFmZvapF3fjJ71Lj3GUx5FzC3KnpergM1+E32WT6v9sa/ucHRAXNwJQpHgKAhlrnP8U9EFLHw8
zEQyF4buAQuXSaKE1v7PuD8/ryHcuNiA7ug6FHhU6wy2aD3+GXlVHO4N4XvZGRq4fvbwjCgCaetS
+b61uPCjVdKbHaPcYM0cdlZe87PjauHKsCLtp7p+L2V1i98KwTItTB7m8wf0gSLW4xT42xGuC1lo
70kfRQSpx1crl1wMCzcFmeVUISbDeWCiAkDJIET+Zl6E4+kzAC2hXl6AG5OBNAETbgcADwBx1YS4
gJPG2yfUbR6NL/T3ANEhhQvxCcVHV/00UzbDHYYk1/FNap4oUto6ytuKu8hx7FtXKpG1A79tRMsF
nmrX13gQrGBQ09eqtzV+mto5MZGC4Xh/SoF3OwBGDc3j1YfMJGx5JUFcrAW6ycOdd3L13nyECXdm
CxJm92nVkyI/xuG7NRMtKt9fBfiEq3GaeuIDW1ERBK+6fKzjtdGBjDxCx3VTcDO46EFaT8oWYRTN
rITfniMr8SBxpBu87pQUHl1/Y1yTpTrMmrHUjiBIFUo6C6XU5x7lMYOwfl6tQrZ33y0aeZ0hrX6B
yjKNY9dxU1rPMeGZvE8DNoyl+ScpzQK4L1Wr40tm4+DeOau8Sq3MIyAFbOo0sVnjsXXHFhL9wOoo
jmc0rJVfkdyV7bDp29G1GV8nkUZamGuxZOaUmX1oPjxj8Mk9nsm5hWjolhaPDW5CbFA5CegQy84t
Y128LqbPuXu3unqp8vSsyW41HFb6pXoO5FCILXvWtnoqaAYjhsxiyM2rAnc/iZ5w16Ak1ttJCJKE
RIV4tFLYNJn5uK8oEDyxBhrtO4J52f7F8vYBOwkopjf5+F/6cTUbNWsLybQzq0A77NHJSWtmrOMl
wRobuu4Trh3wV7yL8b4tMxFMQWIwmnORcfiGBE5NsFk9d5ifc2yKhFaLYv/eM31e0FGz5N7HYVR8
MpCcX3Tuu9LkJ+OinddfbfMI9KreqH+ZCNusa2QSvTdVXtseweiyAO3LLINm3BT2804hF8EnssLS
0La+/4on6tdreNhXQnTwnb77biTSTjz1QdpvECiQ9K0wlA5ChpIcQQe1QSgMNJek9M/J9p+nshCI
7dasrkd7RuvAjuD8KFpNhE/FOIMrvKWvPomRxfgDV3Q7c7+jqzG/yf8jKM+jpl0PY8shmw1ZOvSK
TE2lbtrrxev8tbOhJ0YNjhGfmteL5BvFzgMNeczwtQ6/vkt59bxDRsaHKh+Nc1Ci4h0SlfeyOBdN
tl/IWy3vidwASbG77UvgO7Rc8XEKS8Qyqp2R+/PMnC3pr6SoPWXNInfhyzeDHZ3WqO41f7lnY8kU
iNXFYhLYxxDYnQvAvv4cG/tUqdimedSzYRExdOevHjwgHCw6DRte7nqbbv68Qe2J4+1zMEjUY5PL
fsrTsJWMhyC3OyCLDVfOjwiUgBzpEu/I6oc22TbZ5qMatC8hjaRIQlrWVtG7A2QfzZUF5tOtJfcv
jihVafxOdMKwCdTzBGzHjyUTY2TJbbUGhhw6GgJkDcfzdPCJTxEKIYgMcrBOAC4FAHwuTgCzeaoP
ltQV7CTMqgr7YYod5SC+Qry8nYZ33TBwCmgLu3Rxx0qPS2BnbA4lL1fJ3hrnQ7LYZ2ihMnb93ypr
BS1bi2+6JH2TIZsEX0nLQOPZychEs7SXzZ+skee0mB1y2DeleEnifS99zsTCP2lfCiRI0rVgSjKd
JQdDxw8Ke9M0iab8SbpD2LyzshinzmNgsMUGvcnBAQsh58ds8dAgky0CkvZykS7iue+gqjSSSvUk
sTF+DA8nNkSdCJkvQPQHx9hFjJOabFAmiIWjOoEeT4XBaU9SIH30xbE7FtBnJB9s9vzY4c8LiLhz
ksRCXT6W+5xsgEC7epP3IxBH19hsfU+9v+LGZt/TCWjtnT/3HxIg1dZ2ktPpUJ5P7x2OYwWG2+4b
ZG0OpJwtp66Lyp1mNdmFYWb2c4v3GNdbbWM77EIJfC39PBg+zQLh7lsU0M6WUHYFz8XEsCpUoRvc
KorOQIt6Y3EX9UIWKvetcCmNN6+rbsWnjUvjdYlyD358hBxpTW2e7wiTsE8F1qWEEjJQNgDfgaP6
UOcnvlvMU7g4KL9usKymnV3e4SLNTFMFUQQhvH5hnl2kMIg8rfaDfsM1oMqkts83ZKG8uSptIbUb
xEDzXP3m4JBmLq1HKIoInUNtxyH/QvrriujXGEnX9ioOkZkKB/m40CAcl82UX1L4Fw1hPZdk212l
mmhNpbeEa14HeMsv8ot5CEEpVWUU/aXJTgrQAI+a8Tf6LEaDo5AmizoyZ3IcEIy3HJGXdTOPG5ZM
87aN/26xYxSvc22OYEzTU+wqr1fM1nlnHeLxV5qUjbrqnRdohLgU6gXdd2m29gUGKehVJSAfNhm2
4jBRxxvxtI+u01UHEqZ19ahsJG5fZAuWtufOvxqf4xB+q7rL/ilWhTkw++yqBXYuQjrkGQ4Ln1B/
STk2VDzuh1RqQwxBXNlhi/+6VzDTPAAPBpAGVNQX6eaIGmYYoavevw3PRsgYwauCSf6ZUMb5cRJ1
aycKcyDUerhs84mCU6OJrXKBeIds3Ieqtz7YD1YxIHB6R69aHsWHDPqFgUVT3YJCQzfO+Op6Hc8i
skto9kNZohkmm8E16AEIbPXcbRfUUBwjbGUmtqCV+4zNbZz2TNSWq1/q4lqDo9NJEqjKW718ahvT
9JBcQXHDS2KEckAIlzJ2xWqmdCQIWVArE/yOaXttxPx/eH1bXW9jjezMsDp14b6NkMuZHtNdy78V
JMBpSBkqEr8eYG7e0+uLQ7ch6pCysnYmQ8e003Fh3XCvKGoqf0Hvmh3UwRNeUWJ4uMcxR9EVWVcs
vfGx+F6p9l88vrlj403QZ5Eyl60QUhWu975goFB31lgMZBUMU1Zm7mkz6UYdzfgqouqePjFa+3/T
wFbq0qxTYWZNWBX4IcshIHQ2Um9+POLf+Va9xUtvnTHeO3UE6F/GOmUpsBwGH5pOSIhYl1HYWyfo
iU3YqKsHrAQs0/aG1ulwA/30pBBowADE0/TpLZ0S1lXg06SpBNRKckgpCCgOCELlFXIDEKjXcYrS
HT0q6NJj5UY7Y2MlVsM2TKLth8le9oMfEEeYIlpV0COcDokGdsPfw029ksBIfRMScsBVbrAyhhDU
8KLwINW/PewlNduo1Z0bX6xIwbmN9VBIol/Yhz/KVd1bFUdAay5rcFMJxANdct4yn/ddv7kA1tK6
yDGg48LWiilS56ibsr2QNHdf4Le5YEsRDzAXl7jNAUHKmXzVeOtyXiHw+TkJVe/zVdwAWeU/ewbZ
48lCY6laQSYSYjpaMImffn59PwOLaAOlchMdW1R3LLcKHzjmPx7cn2gqTJ0nxNv2jz56zFQswqzc
xjweMD4FDl3GmniR8bkDmjitCPG8XbC+EF9nCZ9pK0+olkCGRTp9NLdEjYSPVTeeNc9gtFgUPiLq
HyB1mkBKT0Vnpj4re6Gdr4R3C75TLGtVt8+FjEn5m4e+aRjssllq2x44AIY3woAb0Sd2e0KaQql1
B+AdpNV0QRE0BIY/zzOwMfGFavv/EingErYKOf8cBxe0vOpMY4xjNIbsOIx872i/EyN2kNeWsyl4
4JrGpjVPdPQfJ3RxTlViFQuXaDAW4zo3B+K7QsKWzYXTJ2LLPswfycMJvUIjnsnk/YhHE/DhMOcL
V09UUHVpCtcuZ6ZuCbhmYYa06POZEUh2ggOST5OnpdW5DG+HK9uUTiVb1v51gXZ5Dmb4eukAyoPw
uTq8CaUm4b2sS6NlODLKk/7u+Y/RZFGaLHdTK1CPiAj1FOqvviuywVcYJYRduXrhZMSVpSm1TONI
XNYIQK7xKpcc2b5ZfMYHVTxViXzrAjV6Eu8tnUxFcpK8iLQLrv738w5NzATGeUQ4Ksytmsd4Fjj+
MUjFrVvAl1mpIgoK8qzsKUCuu8BgGhVeASXcvVI486xpIYHjr9BNYCdctAKZ+FYzRw634BLvh0Mv
1o7p3igPd9bolye4wMUJHfYOgnjQiLRzvO8rV7w5p9Bp/jjbyWTaEm7RNfe2P2BYKClvEqaLeGmO
bHj0Siua64riGtQxfhkuJR5tEOvPHPvgCwB1Mw0XyyBBN8pVo/qXFc7czunx+Q/9/R0eyGFi+5PN
tGjJzMgmdf9kin/sMkomp3OG8Bs2kYQi0EjNalxcq6PwWunU3mybmTbK94ootAdGFJY4EgWxsje7
hd0moUnJdGiVV9JWtlpAWSA7AMyWogx3uajCrdPObvjOukE/ct9RsMADL+oocJWHABcoal41Hk+l
9tkN6tehVFRSvU2OgoAa0z8QFBU4a9nRNTF9u8MgTvWfu0PjUQbzyY3ivuFxEGmkGCF/ek2cJT0n
jdMikEEO2+9vCh8mwMNNzJmIbUEUIqNuPjhEguuD6B3x9viGkSbvzsGhq9E5zG01ZhzlcgUcBt5o
hCkC8YUujns9/uxGKZZ8lvgSUYiNZEtQXBdbteOKB4sd4liJed2ZylJ58YRccHWj2YRuUbCq+PQc
5ePDmMlyW4Lc/CBdBsNDTwdp94sTN2JcF2b0U1hid4Clg/1Pui7g8OqiLwlcF5cZX+aW6ChLgIr/
q+qOfcCwbzJO5wjUoK3bMmkDreiPi2tKlTCXD0A/ckkTqADg4FJAcWcm3Lbhn18nBI5x+8xpaCcL
sWd+nHqlxaT/N295Jzr+kfMcSWmIjgVPPcxLWQwn27z/pKI+qZXDaAsgLDdWuwbeW7xgvxu/nzsW
1GC0YhHt8jJtEUyGS8gYwBmh85D6EU+B75IBHkmm5DNQiU+24Q4vjN3bJYp75mR/2ciHQ+SM3iEP
v2X526tN7FttT6MkuodlZgoROVA8cwMB8I7ee7T0LdXxoG43xl+yh1AIOLnpHK/pK/IVpHegAJSW
KpgfLZSiUaLie7/zWc6HXrfYTDRw9qEWqsf4lXDQmjdFUBenUznSanAR/gaOpvM5EYsoV1al/hW8
kUFvVIGsyyKk28YfbzpE9LpTehgO23WM/6isL9hAeKx8StJkjNrMfDnxMUy7glIOPRtRAVTgzPwv
2+iwmzkQ8P5qlhTSs0i2QfpVKAiyqIqdYLyBbjL3nnIbk174yRqQe6BSCfTfHRQ27w8vcJj0IZXs
igFbPVG73VzsFOBq72w45q+gej/rU0PJ9JI4NuXmC4vCmw68A5HP3jI4/LQ+E4VPwl/kCJGQPmzy
3wy4AD5kdTrzjuRmu12WhIJuxjtcSkC17tdNLGXzYLTb7mGLJ1YriYHZWMtgvPvqFxVwHM+O1Fhu
efn73P36d+PUpO2AEinw3JtE7Z0ts9yjMQiUA2n/MpeuFy+DiiuTLfED2QHYOXoEINJx+w69TKjU
g5GvOi97x2olp+Z34dzPm/z2etxRqyVAatx4dfPhpSor899Rg0E++VHiDvo8p17OmyYMpzROLjp4
RT6ZprzUqybct2eVGgTLJc8sqw/Px/hm48DuuPBP++LciGggJ7mo7Q04xsg4EgdBNs804wxysWNd
JcCLDkILw+UD6sElHIwZPGrEzlQBGLHucS2ODuXSYU7JPiiY2Q3b11PAAwSE8oP48Bx3uQL3nOOg
fvMq0676XlqzIfW/2vgxb19xBF7Ub/N86K5t+TXEKTrR8VV1xf0Ps2mNNzOYErC8Y1PTxu7fT8cx
zYUK5w56eVKGF+NZv/IFCLVyNXb87rvR5zVNDnZkeioLkSzLCOTnumsZbE3o7+th5HYhZ7xRFaeO
99n33zkvrRtITVP7B3xbzbGAvivWZjNrkyO81ilKqFXyKsJZDsEeTGYeuFXTgGZ9/YCk6My7N2I7
VHLJRIu0SzDITevbunSCg+hXJtY8YEXMq3RuF6/IGoRhMjfVfJmK5cDmeAy1pCayNeVGsJ6r82zI
OGHWXgWOMjP7JjC/zpzJZlxWMexQlin+ewEv/8I0KUa+Kkirge+VdcD1VVdzNyGBOZTsl+sJICfl
SogIcY0SREb4koajn9TIdrs2CrSkoMLuezpcJdaL+yXMGtbNelaJI2jJ2J4YjxtbcrnBAPOCEljp
YkiSsdBuRbLR2zc1a3m8G7nE8KzmiVG+Id8Lywn8T35JjhixxSSNy+3CpeO2fEkgt56gu3Ogh9Lv
9Q13vNuGWV3nZlAPVPZIiZZMHFHpHygWDvAQCLwksCgfjibIYJbBRnaCSgaZ53/rVBUSE3qvlXOz
97dD3cYsJjUkFFyNlxdeoEZvmrnZOscPQU+RLKPBntg8DixCV8ja2+rjOfwnBd/uFxqKE8XV2C2P
6AgexR00Z3J+SsTwjtCEew52MrQVb7yaBzpJMO16wmqrgleqQFj5XGKESVTc/fte78MjuES+1LYI
+C1RYNf2BxB7dKHvJJWrqUas6EUd75samQGkG20bUdZUh5DUB2xBjz+51jDhPM12XMu1t7Q8h9yY
mIOboSGd09Lzp4+4ehmyYuD2QKySSgZxvP75Jr+3w0+yElQ88Yc8Xjq98ZFwmvY6piRRrXDhRWdC
ekFcTl+mFATi2d6GAIxT7o7fXH9pt5QdILjZd64p3qe9NgdgJg0NXgYNVbP02QDtmbP4r1KBnY/J
3HSjlqdRMGiUc2fDkpFuukZXMl2MYfuThTjeJXRY2aQo2yYaJSlpMZADaWvWJzjnUG+RYUzss6qv
Fdzz9W7aXyHbC2SpZKSKQVV2YcFz0GMYhUHWfdw35/WN4l9gvMxaSu1IVrTmC7yJZZuk2ynlK3Mc
LxXM/6k0omWlIVeAVplzqUc4Or6n0fm3lvvWtQPYY7hd22WyxbL0q6D/yL6uqf3Au2M2uCOOkr4d
O6u2krWa6ZsWyYEfAy2hcP/ZJLD4Ae1G4E3SeSMDdpiuTuwFMMxgodn5V97kZjuXoUEXcRZGRYJr
RMuBJCf+1mTk9lBk9cC8EX1xJUfPbTwnoYIjZDhZ02kVv41g6alOtHTP6W9NDlIFVFgpmdRMqE0C
7+IzQWnVtvwkmPiHklwDQeEnot6qIEHmVSaLTOxvxAfS5heMSaWwrzroT3DhflTwBLJm9nwopyMx
FHtmrXB0CvyV3ldiMTgHxmtRJXRedFSOrQt38PK97HT3pKnTL2/5f0vivBv0/qPUIu+XTXOfOrx3
+9iEY/hrQHiaYoLv+l1vbeA9OooCvxwN+iKnQ9l/1jl+EwDUDWJjRdldV0STOYI4ujIv7o+cm0Xf
cspLBjcq7JdPVdFlg0VB+P7o/BZIQpFV/i9C2iEezN68uS5F2Vftyaxwxe2yBpEqQPSlBbKZXgR8
xlnI62fvAm/IjmPEbF3g4xtfp+CIuRczYM3CfDVw3fZ7n+Dwt5iHaQ5iiOyu6TnVIxMD1IODyU7c
14XbFHhMucWfUomb2PJG+ZGwwj3+/QJEwlNdOSsKIoD1bOLy7mAu3LXVoPZBpGvTqdJ6MSCfVVxA
C6Cwk3ViJmvhBY0q6AzAslwu2+SVEka4NDBul7PU0ss1OJF4RnoRc5hW1BKBbNfXbCxPGmPbfvhu
gThK7R8yPYPf26wwB4cMPy64GVzQYkKHQZ3zKZufCcepSX98X5zT5Q1KIfL1tLkjR2trYyk0RWfk
Tv+yISsBVUlLnJt0BDC2OXvhdg/SD3+wfl9AmlZPQ6KkWXZueoNgz/b7zGIYWXwP7clONVGNcJm9
r4qDEWtes9vOfc0MOacoodki3d7peaRJuBMdK1n2nciZKhlb0dbCwI2Rce/3e+eguqsPrylCvobV
9Nrjpn0J1Tfy7aul+mbGrmP5tS6CNZNNS0K2rZXRv2I9Nu1pi6HhCooht71lYrQ9fEHMYsBA2gr4
rPMqMs5znqY71lBmhXe4aBfVuklMIeYiDm8zM+Q5C7oQ+GGQn7mDaChEDsqu1L7wTHwv9OaIIkII
n/Q5FV7pbQTQEjfO++iTKvOgtwkgjRfkn+VyXwEo0AO7OtELagsk3mdLlZvJAqWFaMXY4YvsWkkR
vT/0LEFw6MIf496IcYcd80dMveZmr2KmoNXtPog0XGaLKq7E7GxMkU0+9EAJqkme0jWGo1+NsrkZ
Vv3zG//nut9A0xOQBqONvhud3KYWlf35mA56y+D6RG/NxQxnoCutHDPKTKp8c+Cn7p1GmDxmlMTR
xU6paRRzv1NJhGT2xtCVjEzoLMHubZCPEVd11AaJDoOwqoN4v9o2Ya7XpieMh4vbCmWQBXIxEVPN
8JKx7u1mqTET3iTVlFD3eOMectAU6fexCqr6uSm5s5zZ7acrkaiAkK5pUcYhklDyWki/DS3/YxtE
3Q623RQYTM1EmZRyfbeuuhu2k/SZH7wxWHCv4OnX12mpCaZABbiP9jXBG7uihMwZbJDLEsOfeKpr
oemAq7Bex2Y8vj5qPOb2jJlj7rfSSKLNIChWRkG6jt7AwWmJS2L1VlE0+75RzaZSEmfd9bj/3sfF
xyxicbQJIaRH32fS3jsKP9qFlpQk61GpJb2YQFYfMpH54RFn/Yog7AVSc0tXwQPezPsEk4Cimexp
29XRf7QYUjzzigci2rHdOujUNX0Znb+/PAE80H2a9yZWBrzqdi7w9oTGsx0Dm0F2II36EQv542QQ
pD2TNVqprqScjcmnnqkyNroF9NKg3qPyRUdPrNqr3fwmb4er3HerK9Myf2SlLsTAzoyZHeCgK8e9
uTHjIKS1fZDvNlKkJbPwUQunPYL9hyRen8hCcFJrvQTMv5g0puemZEAPWlYEwUtiDPkxbm5IWsct
NYgHqgxe1kbB91eJFrFEdi9WaREx10StgPljZXus6cPVX9HBtNNGk6oF1LWU0xcUjO67ZtY9ONet
FUb8xWxzDakFsRPcKEgJ8eP5RXGWR7jkptWEEgBFVAPaCK+Doraduj12s7HATALGK4KLCop4NNSS
V+E+G1nL7XGokHQOtwpcwWS8scSsR50LuxIqSzCEfLOV5zqCtxds6RqvuH+XMrxPmIKRPkz31dMb
lfHMJz9APfsQ/pfemkGn57D8XPQy7IUjHY/0siA5HaIzM//xMQ7Xu5lxzWUW/QDnUsGDlGF+TI9H
NZEzqpMe111+2FqTKH2gEpwXuZYOF42nSYmaCFNgjuRK6lENaWqU7yjCTuOhHFtvIqfusokib/FT
UEzgRVb0QkJ0/aYUYsMu735dGuRMsafgOMuWb6Yv4ZQ1gK5LQ4bwUue88cTiOw+3iYtioDK9VKfk
TAsl9yVb0R1Dzqf13Ci9ql5X3Tcfduu0NZYYNuKufidlm+JlHNqOQouIRHzhSBVbEkl20qurGonh
E353ZoGDcbRJGnnha1UHgXTwODjo7rZ1LdMeXCuPneKY3jL/QgNhkcY25+Bgpo3SULx+ONjO7+EU
PDXOwod3JcXdnClyPfiyogQ7GqZs09S7Fl3SVkxf/ccl4+/6MoXEWRXl/p9duM9HlaitpJweFtFO
wwolOtaMe9St4ZdtBLn1vBSUgI6bQvkL3MrCxtAPJuoPp7d28s/nx1xgulR91ruTmi63t15Rc4py
Mu7DlYIWSj4qhbaea4za/lFvELkCd6lt/JJv8ESkJ9nJjEjNz5VaILzz2Cn7WcJ3U3Qs4+DPCJE2
F/JcTHAQmHTYTZ3hgYXu7VYCeMX9zi68cdr7Cq37voAQa/vfEMSi6lbl6wh5sat9uEIluIk/NdvY
eeGCKFWNXp4XsMFjhHRG31RWJx2Z1odwGNuabtEyV1MGcYbACh3iXkUtNZ5qiTuwZcpE7oR9+NIo
sk9o0Oic5QuE8PSJtBwSHEP0dbj/u2zHMO/1ozuMHj4nYmiwIox0PX8KeGyyVS7ip25sNYh/c0WH
c9qWNRrNrLOtrNGLR92+XcUw5Fl1/KITq7uR7RLp3WyCQbZH2/aChh/+x3gYquRef5huGK+AB6iB
h/0Tk4MiSZV9kF8kDsQ3auk8O+FyXT+33qxub5T3tPP5EFP6UuDjlit8OzehdhYIkgYNcBcrty+o
dhoE+GZ8QG3n6xC4qTdHqm40Y2+dUgqL3e2jXqju11HCrLxGg4GQln5qGzO7IPCCdrxHbH9f7ezE
c7GAC8EMAUh3CZNQnkHKNyVo88MVK9NMDe0kZ7/x/z0q/pto/H581E1543sJYIxg9r/DfPGjdNAN
lkGWMWUMFIr0o1X/HM39xaf/BQzDhGF8mkFzw8COcMUpm8NgTK7dENskPK0jeDIR+4OzH5Fb9gG6
kyWK/hfFf6CMxxnpBejagk3XZ/RGHwXvpO8O0ecq5j3dkEbiRUt/VPfsgrRQQHCud7sTsIQCU2Im
D2Tf4XvBsWUL+Pijs+8IFPqL0vz9ZK+d0lo9Sl6nB7pE36sc+bdxk1xRWGZD4S5hwnlVMnO8ik4f
ynsvTPwS+R5e00j42KF6Y7C5hX4F75Ba98ZenwHZU7PTJegfmzubrQ4X6xNXoWJFVonhnW1zLz0E
cmRA6k6dLNCE7gDT1SQlXDcV4CUjDKopc5KXVJfAus46QQp5ame42dJnXoX2g3tk/OwOlB+ielKZ
IFdIh67iOylZmWr9RnfT5lMKt+Dwus4+lRGPw3EvAILUG3KWV2kZEkg6t/s/kZkKjONhm0llgD2d
5z55aKRN/55Ln+Ae5WzPenl0axE/j73dt4sl/otDK+uHTIxkoInAfryDKtVRlW23c/7B185g6bzR
GjxD86HPznKe292iAfWJV/oYgfspjFTtJ4eknw0VcJWfUMDLN3Q1iw9u3doJYLRnleyc1JqX8imZ
IEni4xIVzwC6PXJtCOUGIoKb1aLg2AwD/7+ITXlnNJ7sPY3V5ISkDpzUKFSBXklndmhg+GWvtl4j
C44wPB5FDRulC5NtXFf2tGT6rubGfCsuiCmi5aPOvriuCRMCjLJWRAPWR+D9esqr4wOaIjf1jlkG
jRIwlLXQnKKdh3ds2ovD71ugOlWAVpaKnG6rGJ8nYbzJRSCs7wnYfYwmz6qHibJp36NuzvqKkPPr
/18jbeWJzpDJC+G7DsbSKGQXiny1ZPzzpV8ZFUYUZB+5VpSuC2tOr2aZ8ULBgykcJ6rrMpKT0kJ+
D0VCmSFIc++aO/shdBQxXzZ+LuP1TajQ/0YO6xzO3hTg57BsajEdPcmPFcTXmGb4n1mFi8xbZgMw
GLedQIPyOAoTjujSoORLo0g5xSHxY0i87pymfklgUApVEr21xk6oG0uoZdcvium8bwo9tyLudbO0
b7chpZ3U+tWE+Yal0XHY8ZJfYoQa5FY07e7vTsj1cMr0M0UGlY5eiOGtl7f+lHdkos6Af84O20JR
Pn4qO+opYsjVVsknb2i1I+JzsfHG33LhcgQIfaki+9uwPHeS2SeW5zn4hqtcgSuvMx5OBgNOcfsj
GAX6JbNXtD/+APHCG2pPGZj3zqAJEBn7yLKMISkY2fNw6bKF+m1gQE1Lc2PjoayHVnyKfWBSjMaN
rkt9Esy71eJkv96fwtyfWOv+mYDSg+6sH+1EysyiefMW19T6pGkDCbEguuUscd9XH3odC9SdxKdJ
vaYjmTPVj5A/8B6kJIVm8e/k4RKoEA+eZZ05bkxpO5lbPmYKFNaaGVPScUQ8Kle4O1G4FtUjvd0p
LO7SPZVuW3P8mMWWlDib7pgUjvfFIAs+IpVCOGanFJH6f3BlxJv6qcggJeitDeeLq6roMoN8TeCH
WNe1zF+opas5Wre8IPgNZIJk+F7H9sfoAl50RIlBkRCJHleA6lqLMhN8Aj/3WVJuKFsTtjHjWpcf
gtdzp6SVbVlauWHL/Lb/5mo73EKStkD9FvW8g0UANuBJt/YvHy5GvylHok5AixhRb/KIg6dSNKw/
Xt3kvrZgO+nLFpkRY3ftIaciDjS3P7OvO9KZj0YNqooxufVx/1m7+qGiGweaLX7aw3/DYXffZAaY
pEylQkSoArnX5i/eCjsmFDuccstmou7n896znynoeBo+HGrV6o9RS7Nf5LHIG0B+vphs3xd2zhYo
cOoSjsth1q//Cp4fa+VYzRMbeiZxLtq4QoglE1AuERGu7OaJO2qHBv1lSLbsoxn1ybr8qAUF83Xs
K2FB731r20DEDIfZ9qJAZzvgFC+WCYOGqgwzbq5lIydCybQfSkM3IRpoixEYgX6jhvkvwAIJn8tD
Nx+ZGiJBNMwAbZVnFM/JlesuECDG5T9aJNztcY8GYbTFfLcaDpPtyVIm2J4J4294mtiZIogo5KzK
sC/XXnZ2p4i3nDntI0IPohgsQBbSOncSsvwsu6r1j6+L2cRkBrIYoOj6oUWQTV8qLjjHUfU+o/pj
PCAd7XyaWCq/NtslKnPoXguvTX2dTqC1+MXsVUgt/N01ZvTK0ERthiBPiElrriWOFxQEhcCg9X4t
PPhCQ1cGXNRKq06QWomFyeKAxdEwzxZzl61U4pH2QBdZFIDNUc/ptDYBBKrAQuvJKG+ocGTICjnx
MKdOESg7uuieAK8vxFk/7vFBwBAaHu4TSait0f/Nha98Juc6pWK4bLX6nl+tbj+O9LUvi5bIsxBd
W3q4Z6rruFEf9019YJKsz6ZFbE/N4VUpBZtqUTEk+T7Gs0Q3BOZyhtxhGV074JhZjdhU49Vea41p
36c1b3KjZB4vqEaAoyl46I4A4zcpHxXiu/FU8PoidTDnOpNLP8fsbN6CS6MSpaphZcac9xoPxPhD
8vQwwR4xzEfYjDJxc/BKpAI6xELQ9kXjFP1F9ZbmN3hk6yK8O0MUVCJfFsxddZoB47jNZnKNt3cZ
jG6IQt1F6kw4A+zRnP+MAfw4AHyUcRpj8Rarq4i+wZVmeNZKrztnkpANuJtPSKwZb+efp3LN0/P0
lvK58wb17c9cxy1AxEcl68sMS23W7hy0fPuJCIj/lzS91bCopi5IqZ565ry2//hCQmthTFuhaas6
fHGFsh2ylojex89yUZnV9COqVAKkMPAJMSn1PTCMbPt8rn7DllUvOzj4PLC6CftHVsH/+DDL0s+8
hpoB+BOkS3UMlRLc14ZrlUfXVI4gYKiDDQRbpDIopJvxhtMr7K3lsfp7DKk9oIh9LSbsJbyRKOwE
srGdFCyZxvxpmm3788ODXxYIDi1z8QkpniN/XDfRMqGLFMhwFo4UyGFaak9TRYA1u6EO1ofapiuZ
a7N0DoFt924RWOkBZYqWLQrwBAa5KBKrH+bzTnESorJsNs/EyxLewhw24sID56TQNnGOZYIiyEg2
h637o4KjCVMZbJL6UvlaR9PjK4EHzoFjvxv1qFWAnTnzcIs7yI0BrkiQjk0gBkGfmNTABhMQPbm+
601zbdHbOYGfGewr1bpSmtO6+mvs3zhJEkNSwAdJ2SjWX45oCBuad9O1wgCCiQHxp1Aze5MVsmeU
4V6Fxtj1j7Xi2uXhRwm2GayTNoqJc7NsvMKtS65Z4y2CohqY0DslXBtSkhbcvmLX/suAoOwV6SSN
P3lAo75Dj5UMUSJEN23EXwbN2ZZiisR8nspRk6GlxntnFjVK5KJP4dIU1TZALvHWbRclCgR+CQjU
edmnFr672K9XXLMCU7XYRQrHSeOXR8WSo40FAtrnQVGDx4YrEyqrbB6zX11WEIpmR/V9m+AK6dkA
Tj/L3fexb8GVG1qj2xIVpx3jfLW5pirffd69MncxHCmhStvso77pUOQ9nBylH6VI265hipBYzx8a
Fqn7tbNS5e4IFd1bMNttoCzHgbLSZqcq/meIUCtY8SX259Q+EiTfnXNCJQZbys0o0JG3m6OXVzoA
aJzV5t+q2exG0c3BUWsm4jP0EM2F6ukBkH6i76vKKV+3tuXRPWVHwMRZPMtFbXkCOBwj5MK4pY/A
1Wrm2PU7VRGAgOgG+YySIGX8Q6guCwWwXwamzLQcrqzuc436L3e9tIipdu4H907o7uTmMFp/dhO2
rBHhPFhYDCBdI6l4zX1h467ny2rZbznTWIXBIzYSdIAg4EIv7zsLgXy3n0I7FKzL9t0Af43uKHEF
AJDw+itFyPhxGhK4UNMwRFKSGFCCyRiDURr0So/YOOVPNet4YWY8KIG+yNKxCgxeh8R7Nx3nLIIZ
l2UWldG8QIXpRJXANIRf3Ngb5SGorJFQN8rO3TTqqR8dwm/YYITerUSlze2b1zcC0UP2iPIOwQ2Q
OkyiM8mddLPIh/8uSx/d+/eR1613QB06nMzknwD4Mp945ZKVYzOd1kzDcjH1FxhMzH3w75YGk1T8
Aw17EeR5lOEKuyFoFD8ykdy3hT+nWfAaYfMylnvPgOAtnSfSEO2bBW/hN231okcCbA69mNj4fjCZ
dlI1I8P8HDtbpjc4TAPqqpmutSTJz/rdEKttCIsCiQiCnkvZUixeXfn0eP7B9FUWv1WuKUOBv4me
YjjYE+8w2vHB8e9Eg9y0QM3RKg2LveXbj3M3T3hbGcalHgoh4M3hUv2wMvs2JMgor0x2Ck+NENp2
513Kp4Vo+jgBEFglja0rzgvlTr+ZFIvpCG8rTZcOhpQVGyhY2qI/mqojwyvKlG12LjFM/0tfFlxi
KIoy5ki5jvWggM6LMOf20bAqvFLAX5UwoN2Xwrph/pDOyU4Gvv6vXPxMHQp3m/I2g+jo14DEVOZw
gvNZM03j22p12pXZITIqq8IU1v9mR5W5JJ9WH/UbOxUX6SnV1qVA3KLCsd0MYu8hIOAYchTXPv6g
nNV6P9auHBePb6PB5ASN+upFF1ps7WY9JeqnptqjsZBujd8ioehZS+5qvaj8mBvNc9USljEzB0PW
N2YK2ipwYaeWbNTCwxvnVAE7a7dlVuZ1H7w2jUpVjiGjFDFtS+T9Zb+W4u7dP1TIylqUBuL7WpZc
082AjFvXj7qvNvjYbV8jTfodyPWHu/11RBBjkrET4h14D3aYjzr52R86lBcGsnO0JXXCd/+Q7nyb
VoBnaw+r4dH3R4MCpUaXuRIxtuzfjgS6YZdnxQC3u6AKf/j617D5ts5tEaic18gZHSjHtRF2k/Yl
XKI7QfSj4LblUGdyUKZf4ebB2Qa1MqNAKQ64twx399cNi53JWdImmuKjLp/hF9KmQIxbK9gibuT1
6U6YftedyYH/XFErFlJk7elYpN5RnWQFSNu8P/905zW0jiG9MlnJOr4xMRfiJZyR3ugL//uWEeWB
uzLG/pZUriFWcx6lSYISdb0jw5V9w++MOoOUIlH2DQDlEDkN3nqAmqU/W9DXUo9yU3HiIsEiy1QO
f119W0sOdRI3YYmatD2K5Kwdc4WTV4Gs1iMGpPWjqL5ZJW6lOgNmN2Wj032I2GvlqAibvEgJ1H6p
CSpR+ZLafHnOEQZksUaziU/X0O/wn1MeGmilcyf8V1OhNFRG/t6SK88JDh7ryBpBYW/B0AVnfjRT
9gp4O3osQwH+T+5xNS2wVmu9EYBvQjaLbHP+nj50UmrdO2uCId1Ig/PH4KEojLqtkuSahUa/Tcrn
nIHnkZoAjK/kCHHUjUxOz5mfxTNfUYeezzVmfbXmWXMnPqsq4r1BcpBpMYeW56sA357IZGQhApyW
rOjn7xabdlUNxedLpJdkEiWuH4bkCQHQUO9hOMDlOyGTpyjUk31sIUdN5eLl/EqtyCLRC02JPI29
tF0rbdXEI8EnDPTtXPrUrj3Y/9Av6J7aRLzoJOZoUFt0/FV1ux9K3tDdrrtWCcJtm/D7Lq2lkxD4
wo6hmCZ358K8QzGnGV5klq30bWiPW5+A0suxsHgtudT2neSyEP4Apw04qe6DEjRQJfppG5DFyvuS
fGC3DNKlh7uG3poSRnpLz7YyCw5uiyb6A2Sp7wQeirW3ethrqlvMNjMSYJ/nD3KIt0Eftg7dNgDH
7pFDTA9g4Wmv0XZtsuV/qs9GTIhhYa3in3XN0Z0WsnhynSnnDaUiyc1c5wTXQn1/r9rb283IolcK
/bA1g/i9GybM2jPEAbnwokXbRW0oSjhMS8gx7ymJ2ffcqlkja7soovIN64OKy2UZTeNfEh3oC+We
MzI9Q83XwF7eXcJejxqTk8zpvgJBwSL/OYwwvXpXqk8hSM2iciNzI9h60nBGv63Ukt0EheSxmGJT
XN9/H1SKYS1BpHYd1LbGDBFUrOqBLI9Dx40Wo491kyouY5DUPmc9OQ52lwysLNdO+UZB6R5p+L8w
yjra2nFJEagDjcN3I/n1QHZoV1yav7YneM3ACbWsXaUKsNrb1agPkk1QJHKIxF+bpBV9NIpZrGpS
nuqglVru1G1Y2dIW/+IT98MX5PVz+ueo2FJqI7Z87QDDGGybH/vGjf2wX4m8wNNupz7nzszPZ9aN
5sXvMRE6/O1R9ZuyrzWVIlU4YsnSMgjAw8tPt4fePqd0F9aa41GH7JfWvjSMvxgyDNAAynZvL/qU
fiHluBynjc26qvApgmeSLQ4L8vuar4m2L/tAxB0ybxPAEpTJecIHI1wE7kpz0HKCBUzN2pjFqXqX
sLAdJbGEEd5ZUrXzRb0y7D46U29AS3HgRht+uE45pXCJprmbL0YdZDx0wD91SQMeJCuSohRZ5N9c
xlEXrQS6gXypiNSzpZ5iPkerleg3tz2XT0nhhH3DLvN4Znm++6Y24jyzP0/sqrB3JHkK9+KeS8Gx
b1XLDZjLyp965rgEerAinUKCGgZHY1EalLbgYGI0sCEHuVLRRnASAKbjvknFt9ijOH3aAhFNoPBB
6t6m1+9nPlIjhWMSqnQD4rfy9ASV8XFp1ocvRLI2SKLz1ObQ6g0f5sQukMuoAtQe3Jid0TIWZs8k
DXf0N/0RdsgVyh1XJtM7rAdhQn/yB0lqZXN9/h/v+gHPxJ4qJYFAW1Qt0kaXKBObMdnvC/lftIsb
OesMC7JCqJWgplAoM8drSw3soT7yKgEp5J7M+m/VA6YaoEUDtKZUxWKBWqYwYyin/TSyL182hRbZ
BPRzq+lR1yEowPwIRPAgFyEA/Z/7fv1hq1qnDrQ0223V/yeLJRhFPEfPcPa+9AxZcCg5X3M1cKYB
furfbRsuK4W5nJvbFmvbQQ2DAqE3skeKoPBVG5Dl4LJ+Zkc22rD3tidesQGlY3tEXPSmZ5KLpS0+
8PTK5+HgNCJwb6cfGDj2k2AVYkx/PrqhAA36iMzWRIBEkRWKucEhN50GXzqwZbRuEMfMQTnVAyss
bWj+aWSkhkJ1r+Y+q8fnLMFsOnGzDKSudWfJwvfakKaexR9ggZDgflpxmgRbESAIJnvG5S+2sAAJ
I+xetaOzV9NaLsAraA1fktA8r5cw0aQeWz++/gkDuoVG93bsNzaljsa/7yvb8tTmJSUmuyP1HTAC
BilvpP52ka6IxpEJwb4Tq9OK9LQFH9LPHwQZXBm8CBpH+P+SIp544yB4S9bQmo2biTumcAYEnALr
ktHorNYnuvO0Au3HI2V31oHrRLr33cZNd+roIJqznfpypvrDC9iS7iafpXdyFp+vufh3M9vyzalU
w1JfSW4Swz6ZByStXNE+3ulufERuAsWDTLL87f9coqJypDBT7N4nnCGdf9TfX9qSu8OlvY3eCNva
qrQUp2IkTA1QR2K4YHa4g3V9U7AIw8dYdbFW5DDQuz10iqg7fgd9sxV29y9d3duV8hy2cPSFlqRx
tvTubOywcVrvUaW1yQXE3uVZYkXSS3wJJOTb1vAArhaa/tcb6DAfHXgvli+5eUKCBqHM3+LzsPgx
S5qhh24Zi+51dB6fUWSrkCJVrgkUXZWWbwun/m+HhJAIcbU7mMhL0aMYG5TjNhqwyzgccxrbVLOL
HiTQp9pVPX9FBFgRhi6YLyUwXMDtWiU7JXNnf8Y5aHyUNc8R2YvlTiJ73hMQYr64guA+m4jBIYdL
g9Q2MWgyQDDaQM9Ok98VW9wiulUYDXG4IVCZit2NeI4rjyELmlYxA36JO1SBy+4bGr41kei2Nygj
ir5A3Mclk++0c2ph8Ua7u4kclvU6aQVbHzdIa4uubV791tfBxE0skUr6GQttvSmYokxDCV1hDFqp
UhbcfMxos0bU9lzjEvhNj+gAaTDSkf4Ohe231CVAi58SQJtiZoCsdsiO3eqFVHX7kuxDtbrKb5Pn
7rHQBYxYvTDCOxhDbED9LpIN+44vloVJ7+Uq8uRG0avR+5M8InMzW8woEBGoKnrtn/VJNeCVE9K6
5/vZXbsrN3xNFylg9VVbefGb5BZPJYRPJO+hLzmJ1AjWKtDctm4Jmvv2HrvEZNBlrfjJ4QaeaP9Y
5LYw1OH9YMyhWicOSiZ5wxgUskaXaW2TRBxFoGQSLBsJ8hsPQK74Q1qJcyyY0qjNyigjE1VW93q9
xZgV7sFtz0OKWdXeOf6dNTmuFuy5oGjZU4XOmZ/cq7xoDfkodSD3p06Bg2EzEbmflf3IwkFeKAQu
cEbw1twPofXUCHQMwaibV+CE23TpPu8cIiWCSjPFYowcyw3CldNlZSNB1UP7ILzdC94spVmz5oQZ
m3qHqU5wDfZ9+dQM1MP1T53lDLqV9qnxMFjEfXqfTKTnUplx9KoTFfoijYz+3RbZCpef0BjBM6l3
TpPRdjSFtXSDJnLQ50ypwX4YfvrhnZtxD2qUknk5tiltZJs6/UnzGS7h1aGHkq7DSk7/Ng24ka9A
kRHenH1y1ROoBe9NgVAs+mYWJV8lV+mAzbZ+a8vz2J5RMROnSBnzKMcUGSwYxp885blUMpFrqKmu
JAGNTXFgQlbDZqDmHGehW3jtT+TPbGMD9QZX/rWncMliUzLwrRrRZZRTR4eqsSQUauvSGaA414hQ
94f4d2oH4chvgoEmeXNi3WfG4Yt77Vp/TAp7TbiQGjFXOKjNhOiXlKy+GibWi3IqRP5REVsm03X1
2I/0/HupZclrLVn7LCuLthR1OH6LU94rDw9KPnVPf7gsT28GxXQ4yQ0flfsQS7tLtadMxLdqS0EU
vLVNmJ47m8Wq5vhjs7hiijhOcLDsfChcH3LKLz04vA3t9CqdgDydeyXIEbJbJHYoS4veCydXtEIw
3va6owQUjY8EtEE7k2piqMl/+FeT+z7AVwBPSQfvMEut2SPYW+AAtCzhPsp/P4uxJo++t5OOZkI2
RTNZZkhFVzH+gLh1Pt0Z4y9jbxiBR/Kkorwz6qJNRvbwGFnsvgFnaEJYWv6duSO0h/HHnj7cogOn
mVKFIoGjpGKIYK6NnT16aHUgNoNzbldAFM9OgiEKNfB1IVO08gMrbTGk/iuS80lUqeO1Mxg+erzc
GhpFjC/Va26CH3ZhYYAFC+0o8rw6z7auJJNEjGmt+Tzsn0WIa0b6g90ANhdgpkhjElr0uvHbmwIf
FI5A1CEHwVSsm5N4JIZRTdbWo5beYShjhWQWcjWggpxYeCS3KIlBA99g0/qQ2OBF2BJYqJL2ajke
wTUtejmCRulAiF8cNHYS1aCexX7pWiE7WjCo7yKZhUGZUfzOHkyljezd+lOY+cEXsfZY39OH6jGO
iz4Fzn4UuhwShKqCRzXfc6XZ2KHagTfz03rJ0QlRS5E2SOzrnd47O9k6nPRw4qESE3yOjHfPMfcI
Ww6/M+QhwIOb0y9geWxHOa7EmQOJaF7/e/GjFY2Z1Recc84ejjJu6C9aC19iXM6VBmz190DujaKQ
oWM4Wx2OVs89srTm6F/co2yfhdd5oZctWf62V+gveLlY+Wpj0Qjdx/75hRKl3Ocbacx8HGuT3hI5
o4j90keGNBYRVMhg8uU6tpl/DAlUNr+ZNIzF23lOHfXkUul7CEKcjRpldMSVkfTouIx3Xxj2cpp/
OKcyKAISJ4tisfJX6iqa2S99ry5qT5IWKqydvnwHIy4VHEv4OH3IAYlRfpJoFYzaOPPajMl0xGPs
opZbxT/jTu0NQK2sSYdZiD5jwCrY1ey4Ta76k0AW9X6dhATH1XxVOvyth6IbDrtUBa+VAQjCi6LF
FDdLbgt7FYMyObQ6ySC9qzjxHqOQBtmj8o/HD5Z5DKPwMtiInxgAaNCAFmn547EpU0Q7cV9ZjNMK
8HCOcT875uLTuCF6IepFA8U4Ry44+WXEnUBYwjNahsDxUsP0a68RzJAggPdPvN9Box424hN+O1eS
pq1aPbdvYOjhhNDJKBt2XbJ0kO2c2m8/yFeQiOafdIHyWjZot3o8nBX24MtP3+ObCMPGIa0AuSv7
V0lDg3lc46Cp7hLgDgnr+89tPdFwf2muOKL4JJlWVrmWdnA0j3PKNAdmQyyRBD/OBX3xp2yGiTOV
gpLzeFkOsBFCXFVNgim1vZj72pVj+0VHg5AUweNuvjWhUl3x6X+KdEc8KzlMm5rIjCDK+pKvFmXL
b0r+AjpzDLgaBCFVuj3ci0zMaZKeHMitaKyhasVkRqWzDjPVM/9RsqQhJtapBhS1b9s2EHQ35lhA
RwlISNlN2kVGI5gFlOBIAVN5oVOIjhdXPPVHtSJ44v+JEMc2smhKKhXateCdnsfLIVw2q7+jmRfY
mLyWdn0jKUMRnBPFuFfIxkednKOQeXHAKahCbccFNsxXcdN3IOuTgbhDQoNnRTMBT0KMRY44OFUF
awALHtaUUOcatsWXhMfUcLt6qFLIlAj3cqjmDrmKTPxPlxsJrsbUyMhU2Z+I202yH1U5FxWANN2/
ti8Ziimb5YO6tmddbf+cemB5bw/AIhR1rKbBiUqu7txgMt1oOlBe1PpvEQn16qDzx22q+djaZlyJ
IbHfYTU5YI9sNUmEQNueQHir1KrKYdfX20BsyZ248VU6kUWFKUH5YrNyawa8AL3U33GNTms9oTpO
UoIC+1ougOqang8V3QEbjhbW/S+Gj658osngZD0wOMlxtprK/oJ+ezFs0J/4ycxqweRRgD8z373p
IuALArOoxU3tCx8xo8iTA40bFvaRu2lm2B+vB5UshwQRSfYakZgHgjAvjWD862yBOsEztIWrZ8hE
Q3e7rQPmXPI8VYyuWANmfkJQU/Xa6M2gicaSRcK/SDVO0cwTQVm5M4lxYR3vtKFK9+I7hGxr8LPe
HtLRueftdxa+lpMHVvHhv9HlnCExBP6lwvy71BtG7NaJUqeAUe8C1PVEubalVDFtV7WWDs3n6ZgZ
WD7Wxdfy4rSjGPpGl4k9V2cQU8RBoJWHs+v3uRT6jjplGDdskuNLsyYlJxRZvapal+C9ZBCxqfEn
vbpf9rX0UDv3ehieEAMp5zcZK6TVbR+tEaFUKnEsaDVcd9oCGAL4VqyYglL6U5ff6ux4BJhwtnH0
TiNVxgTgGe9sFBws2gArzNUbE7qHte6Fj3Kd9JAjInlS/e11VAtWEVh8GG8dfVytBLjMQrTaFO6V
velJIuTVIVYSWBw9GjPgPseBsNevfY6yVrq+YYwFYdNhwGTaCtNXC+IvtPm5vaTanJtwxPGn0Ddx
5fgxqf49qOaqlxkkfJLZAg3Lx7Jen3dB+xhkHC29Dn39oI3/L11g5ZLCd1AuuIcY4LprUIdpmUzD
5+YydnTtMwAWR7ZhfYOwYAxELLh1n30W+cH2eE2gBPFuLanHiOg5VATUT6+wf/fwPq1mOAjEOy9Q
SyESNAgM1++OO4jHkGcAcsJ6SGc0rrbY+hGrlnc8qSzInbEfR+wBpu+QeUVB5C5x5HIjnnfit7co
0Pl/s3Ai0enPGRKkdqEZVNpJvXr4JoMLcqiIjyI/23M/zluRjjH18rsdZvu6jJc052GBKYCYGfGV
mVwwiQAspui0HA4aAkBjnUuKRzNec3juraZnkz6Pq01FKXI2n0kKG70oh2qNDZoCyVlJwtRmyxRx
5GtSdJchJPWAVxGghh48A2DZuBBJDUd4QJ2DNi2D4CONFyp1lKkBG2fiSrLpQtZacO4iQ4G0qiu0
oXWoBNO1/oFOfzmoY0rvEm5EMTsZpx+OpIccWxiyQT9vBnEoVwR8RfudXQt1YJeGe8fQHIkDG0BT
+jksnWV2ogZlMb9Fp2b6HKlMpQkquGzeGzObAG/ToxZmahcaOc5KDjG5C/Ebzu2HaD5sZEA4rreY
R5bazqCEELU6Pxp6TX4D3agHOT9oKXybxfjCL2QtULuL62eSfyf4thK/skZ77obVIk/L4V0pyD5P
VeRInbBImk0tMLrM86Tp4oIKOoZCM6NUN7tNBW79wLI9Cz/fpN956NWP+MoeZYTXhCllXCJU6hgs
4F7E14TBXWPsfFREVItIoS17OIbNhWkj126YOZrbZTzxfnp2AfZNwbQjV+q0kFkGfO9jo3bnKu9I
s+0bDGzt3qVpwAt+C8EH6Yu/UCdJLxcbzk+dig8ijYxGiBoPr26k5H495UX2BOm+9Wp3fm4+hnck
DcIVA3kIkYg0xeSlH+yCEtdaoJsLSVClQql11iJ3KV4sF1FerGpSN9T8I/i9TuHXbvInKEeQnco8
KCcw7kKf3fNsPI0mV0k1AvxLaVzmWv7IFylVAnL/cDma0SPqhwMEB5aJJ03SxAbegpTTIUwAl4p0
GvhOhbVs8zNAmcoCk7kuT/3135w7XiDOd6yKhXIVhVF5tMzC/5w+44rIXU9zwL8sDOgnyeatxbCk
xrdsQQzcTEtNk6LtO3hp96GNZRl28PW7EP3YtphsHtUUWILXJH0mf7X8175JBBx6ZYJUHjy3SH7C
Sm81ffYr63LfXZbFMWRifCzudy9x9FrpiS2nO8CTEYUlQIDZhPA7b1xIxiI0Mb54G9GgRNfJfZlN
q/nIE+aMIi/cROodI66H7QFv2mHjpilE9wsqwfYGXmQl7kgdTh/4OGTenMxK5Gz/qFCdcCtL12OJ
PBEr+abuy1T78X7X/WrJKUkTDFrh3kD5htiSuaDvsM1uHmUOxceh4VTKvUIVdMvdy1gL+LHWXoxa
z9Qeb2r4DacF8zuAQfwgX7ESupmno/4p/GfVaTjmBzmDAimlyRVx6E4Y80bdTrsz3P/0Z6R0PRVU
yggSXXrAPty6PccIrkjFqOzigFVqhy8wafNbQy8J+FAb/ThU0gWhIiBjq1z2AipooG+TuzX7eW3P
Np7aXzEEFhaiaLWGdP7nQLLzhWq6zPz72wkMRxSdbp0KXu7khEYcj7OP7JRnFt9P59WtkbE9rmtw
71JYdHdJZofmzvE2CwiadvCjSTM1lCj7r6YB38ZBNZKZCsgC82Cwr6PWixS8xhKQI+3e+3vNS1Vn
0S9TGgZTuYlb5N46RuV/nEouHKA5sU/Nsk3aGpnj1pgWl6Sm2MiSdQWkfdCAsOGmTe8hAVrhQOHi
FSBuqLcVXEhD6/kCx8kz9jWDOUwV5eivDPbDjw3f0SeWdkvC+KjbupLIDbxBzutwIPROoB6WkAzZ
lmYxye4GLDaNzZhoAz1k/2B6tpcv7ABghjC0GS+9Z86F9LaS7sVOBScZek8UV84zvmxl34pMsxv+
bojE3DPBtNUXiHm1ES2pW3ugKBjBkZYhVnXxMtQ3wYvRp9zaYoMlkSG2kif8IS4iIeYWrAtnnJKd
AQdB8SPQzAFcz6orU6JxcXYxRO45NY0Y7PlH4LaN+pBW3vEWkHp/08M3yquixv3hIr9kV2NKkKSe
nXI7u5IIuwBBlvbLdd71OU+0Tmelo4WYLMIVEZDqpl4hd/JUeCYPrZxKu1JX7y4uB1tT5KSffGdm
WM7yGszLJ66w91ZUgPlD6VdNlmxoAv66aHQnECq+43ozFWXrzBP02cjCRKS34l9nHl/0/aq2hWrG
yxpHsA75hI9CEwxhYfKjv9X3fhO0fRWDaJoLTcQYUE0eQKoN2l8hMTs7qUsElDn0xyI6UMbAV+rU
g3sDkJshtCy8nUw88nsqDNKuMtr04HeOLEQyIUMDCtODSKEDmihPayWZft2hfqQt6TZU0mJtNBGv
EdKoUliIBGaeQqS+uloJV9nAdsJsLfR/h5JzZ1zYjlRn8AyMu4FhylYnG9x1d/CZk7pb4YoLYG//
oFdnIs3Kx5t3Kqw5ZHj2DIN9w/pmiKttStDeeEl2jHM68AYOt7vdy55ifIsCR8qXLlnKvHBDPc4O
vIqbLz25A4uLAFwGH6Qe8hD6hYPJuw2QaQLp/nJYlZpv7ExkVnM0Q3XAJm02yOXfCzScvzWtj62x
WtkMQTL7R6xmdlq36DlkWV997ut6lR39wReY1c2sD6HqVV6VsfGX9TEpLibdoGGdDU+O76QGmyH/
X2JeLhJGJi2X9fuSJMtPunXrAk1ochOs3qWCPQBA4kt2tg7No9lGhZe/+zyavPApLPHUrUsPYLvj
k6GA1oPOUBdRHSnWYhm7P2+KSq699cVL364kw0lOQ1BRCRUauHEZ6tE/rZElNNxbN8SAbDyDsnJ2
ss7h9lHbchIpaymWkxfzMvO9d09LIPo6Syuvg34QZPKFy2foQgSGDyQ8L5xJAuT4sqQd2q9jdUBb
QcNE0/j4l+hi+Q9DB3f5EU+R8A9tSZEeunwzqaszmi+4lJ8B3HtLpIedE654XK0rQlYN6c5Muy8N
d5R0+qQhbiN+kLt4N4AxjubkEOWtP/spSuLaj8zCUQ6oLfQv/9EcSYhqn4BSLb7WiJqR5MWsYysb
41RlGStMQZ47XbO1/8p+Hz+fUIojzVGf+wH/QBU9nzjfbsLuGFBKSRVJifyMtoTFouhq/aRKRX5O
mzrHH9A8ghRYf5hpy7q5OoHIP8g5Oa0+yE/f8+Fo5CaEbcD7QQyURxz3bKIboODLyKGM4uYci38l
KarSFxgYEm3sKU0bWbaU+P4uNAwMQFQUdOorsk93k3RT2qRh5Wpb+a+V7Rp/teg0Ql68KbtDVxoJ
ilnZblfE8ZK+ps14ZIH8epNxfVhbM5cJ1JLif0ELgKtTe0SIcqru9btfc3TncYCvj9WqeOl2A6yP
qs7loi0cNfQwBaswjBJfOY71sqC3C39Z9s+dytdqK71voKJ+Q4t7Jheb3CIj+BBxgBhSLloA6d7o
V1Rhux0xr7gfKoWAGNKu5sOmgRojo+Bb/m3Erp5Dg4b6yZLk5rQmqSbZVPghjp35b30WlIkSjRln
9vP2bOcBn10eTOVZkETwDPyrc+WEKnRCoVy9IrYicVD3Q28MyV9nrKnQ/BCOA1G6XpWofGX+IEqb
WGc87Ndk9iKDSgfL9Y8/X8ypxdEE/CLVZOgtiaA79reyIIDCGMKoUopffylCV1Fou5hFbDnd/iCi
gbJBdux7OqKXneZDWumpNMaFN9jrxq+c/rf85nXl233jw7ZgMHAQnRYZwwp5gFpioVqb/4W3wLiV
w58Up9Y3YRDeSsdz7Pu7zghrDc4ogXmTmMpZ7m1tZOGl24amughloZ7tTQOo2IR/aTCr2cGUA+gg
/GTIiKpnxdckCyaStyF6ILP607aSPZbvQW78uCix2Jk1EOcKp7frcsXqqm55KK2bOCD/Rgxumlh0
Py/zLZe0pAT5EOc7+IY88gSlZwFZXEeq06xFjH6QoqwCGyTpjAQWC52elBi1qWwIIeYFReGu8uBX
FZSOJg4N+pNT6wc8IBO1wONXTXWWYb0YOWlwFhPqCLJHnjqAYzmOJUiV4B3LxjvVq+5UERCQm/TB
2ulMr5sigdsLgngBFfEkTUdpD1VDFPlOxA6JlCCnHPuU067D5gDipcyKFh0ErnJkNHGItvchkBFo
C60gF2rzM4DNa66G950Tf/9aah8huhe78tTmSmoEaQrZNBfiBKKCwRVAL21asYFXwE7/ARc5V94i
VmEsWd4jl4D9xJvEh2ut5unNfN4GPUPG27RL/jBWaUQxNmlpc61F5XbMkbUhWl7ezxfXX5x9LcDV
Qd0HkgvSCLIdmWvyVaVeWBkQFVrOvU459/sWnB6cMUIr4wJybCWHKd54WmCOO23Jr21Ii4qITW6K
87n6VizcsTlUl5YOyioTT2Ns6aNtzVFrNyleZiJQuJ2z+siXPEsv3s86Xy2ot/C5ypz1DHtv1pSe
NtGVBoFpE6nNcB+Xru5FA+Wi1/M8AZM5KwGMsElmFWXNT+FOlmJ4XWpooVG3OqNsWuEChyLzzWjZ
XVeuWpUtGafwkLUVwSHMBrf6c7pEd8H6UDasifFowGuNOSAt5ISTaJjWZCitBvpVQr604ISH3UcB
zLgPiMr7mMpU4cqyZfFcXeJ7XztohMIiK5FcOiC6j23Jw+ED+2JBeHjbItvsjR+H4EgfQwGfObnf
FbTEzebUgpJn+8kSPz6bLJO6qWkOQdZ7gz4qi2Ey4pWA4nSvZd5SDkEHWQMz9BgA3orJr5dTGVQw
HYILBpENxejav4QUejvxCbzEYQRfzFUSpd4KQ2OC0Jr/4KMhrMnWZQ5XvOwC5qqq/o0rbJaFBdzj
BNOTZGTP0xwE4SNnwZYOkF/veHvymNOA67thyHe4TGQuDI6PKEhcQl/IFd1FZP38c0V+iY4NqqRP
tkg+BRD86YFlRsny8iOI58IBkksrKbtTfTnOiMI3n1xW1R7tzxYWebmvGljzYcCiBUl6kNQc/zDZ
IqER4NGhiD/eQlqTHXmsiMXAFxicW8FN++fAW5IcRETPsUHTjHvXIUKfxV7kTUQgHEPb6eP2ukTI
+puO4lzelNvyMVygn2ZDGk9BjQgtH0UlYlSRpSqQKYxacHA+rKMlOpOg59iTJYNXXicghwzDXrl/
ai8f7JypYMfvxOk6lwlo9w+FBqrCIHqLbLAFDqlz/woEDzuMmpTnvItQCKjsBJeP1LfpqsDW+On3
cagwF7XRaBo2KFH3a7nvHJbVYbXDY9M/aQ86A9O0m18EXVVRFvmQG3CN7ud4gBMcOb3choZtM52L
5JvD+9kXVdCJwX+9lOm2Eu2XylmaPng0WTdk+chv3kSnelVNMBj0WNxqPHEdER4MFmvSDv2J3N7Q
7r4Whgz9vVVQrVpDnrbenevu0MYVuPuf+9iopaegwLgfofu/5E2+22kU/NZ6NampDN1H4Ow/y68i
63SJjpcFeTiCMJy950dFcDed7ZKmpnWmVj7JRvEhbZfi4JnUuvj6Wu1hL5jIGyIceiQn7LsCLQPK
M5U+GrnQp6G1MVbM+6ZzYgN3maIcWe16LT7NGzqpg4/5DIvWh+Mc5UdIcXKM4g2WjEDm11cFcoyo
5X3jkDN4psw68GoZ4ln66YGSMmx7wHCGF69S3NfRtGjhM3XBo0sLXb5f2GFRFOy06THu5vTC4eDF
Xil1V4Jo1UNWFw2St2/BJTAHeIZk7ufoLKXUk/zEpPBA91rIAgN6A09XlDP1kcdbMQ918iGvZgob
LYO0kUSOCTPBPN29FfZ3atQ1RlvvyeeDzzAjrVGX2ReopKWmOQR4DxycZQ7mDNy6xqDaparsjczI
CJ4sPmEOqqGz1uKmox8LwWckx6bHK+5kuvSSxsGG/UtHBFZ4NwPdKWtIx7uOSPEi191FRJI5rjFs
GUzblxvv4QwWyHzk8l+oZYphNuorcacBm9j6IU1GZIhHPLfeJGLhaHmU0WLr4+jT3d2jEfGebZVE
HLIaZ/rcnmoEtsPLU6G6j61hIk3mpJymaXj2q8y+m48ZtN9Q5pVFhBb7yZK8gohQ1RewmC8a1a9+
IdOvUplK0FRsZlI6KS/sBhY6gUiUocxTccdm2yFiBbMm/jkh/pf401m9KsgySfYWqZKGYjxbNUDQ
7aeSSqxUShyqSDTJF9TQfUvyCmolaxjEUAFAgpedenmk6ino79TJbn5aNWzstqNc45+TTYRp1vv7
YIVgv+4lpLms87mtku3+X/MZbxeOfh96j+Dv0yUTjH+qEXaMx1U9kJTSVSTZe25upD7wH+6EnpOa
I/46lS+miOx6t0wNULNzXox6E5beVgvXctZFsvASiUsS4xNvqE3GekrbyOSmoaLBTjcqVfU1fY4z
usKa9vq0zikLIirPK132d9iLC4SMwNODYKaF5SoQqbHwPAZ2Q33zo1Ip+K8GzVTIz5mhUbL9c3Oe
VB6BNDOrqVXmu2JzSZmSi3lNjImflJJD+j0XFfyf4gtxiWN98LL6CCt9QYaur262XHe3kaBAf84H
o8toNbV2xewV2jvy0DUOvaFqalbtaOiPERRnfbHAFAH+HpJhw0R+6Ef3+Zj+WE4q5U9zQZxFcaQI
dYkLiy70ySrW8qfD6vAMm6isHeGMsdeQprcnGqqX3ccJT5QvZkcCbc45zWV9K18XZrYXv2pYlago
Q7OAyzBy2uyEhSfnnp6rzgFAPh5lVw9WrXiwoQPuPzNj/vnqTOzPXcF4dUEXxMdx5kuryeDqNeat
7tTOxy1u3i4PVcTOcwlkhD8owILrSBYgnHngmwrsyPz9nivZtFPMSE3k0fEIjz8jmJhPjNDndYyI
kktj/LV5pCtuaMMPRVN3HtJC48jDxAxk3fkuilEq61Y6RB7XJKTM7UeDHssWSXUHRycOM8fTSX0S
ioix3crKuqfR5fsdfwkT0KzbqNfROzxlIZfJQSUYfYvjGhB+9zCt616CdEHcPC6GW3cdcB5SxWTs
0tqKJaR6/PvCAtQs7O4Zp62jTwKPjx+5zfXpu4hy2M2Xo7Z8bvuMdVia/kuHz20YL9aZhdRloUAA
PcCAgxeh6psZzWRut/WLtPviBnQxpeK+OnepqiDjmQi9VUmk3OGf1J+OQt/iQdxygtldCPEBLkFa
s80zkf/uoqUD5rFtwc5T0Uop1c2yRNpblMOFb99Ymv81kcmV9DC/jPYcsjud48ezf9s8M3w9eks7
RliwzIna8LCfyKqZH76WG6QsWoD5Op7CmGwlZzFy42AbKCgK37Hi9rbwr4K1ZAxXQboZnjcbVnHB
DvBIYZWhIggt5fJ0Gog0KqDOcTEqI/JYVYnIMjOyFF4e9O3GnS/O1KtnUimdizHBiP1C0xo4Y+1K
WusbZOmLliphyZ34nWOXo2pdstGO0eplqzUwXvMKvmCzMK5Prj+9u7WvIPY1SmgfEUKldnCj6NBx
xsLuxhJO6oMu5CIehTzjdQU0e8F0qcz5vSYW+OtHUBu40J2q7XfMX8FFs8s7M/RqLTOP9K3WIook
YDQu8D3ptCuy20cA+oTI9jXIk98rlSEy58PFITXNEGK5a8peOgqqS51gGDhzLxosMqEvhujyPZ2J
00GBsDJuexc7oWsuLR68LEVJjElpOtx0temVUxPLtPjySpMtD0/S6z98KurYCczJfzuW2SjQOgdq
GCFMvABgPAEzwJXkdfZKDpnDBTWyHYTg68sS7u70uUo4vE9pDkc5yBnK7LayEse4g61uu1vspa1K
HcL41gHvfhE01/i/Lq/IQ3egRlR7wRpXbW2z3L/4F139FvphAZVR0v1tguHVzid9bhYttrL3+pwr
mBWRMu9M3AIAR3H7YSHp4mH8GiH4PlsYh52wS+hgT84zZRkbzpn1YuMvjlo3EuVSUpZZMLktFwVJ
F3t45murJDxlYp4dEV6DuLqgdI02Qtj7zJ903frP3r9tsmfFAh4hP6EgPfod2ISqPeP0qf5wP6zA
Zhk4zyF2l3rATxnbnsFmu+OCpIaFRtFEuw1/Mu8X5OBA8FxuoolfU8f+5h5twrrka/SkbYFJU/Ku
PN0q1vpFJRN2qT1/Gym3b89PlwJIt27cGVp3wWBpwhTOfNAa+rOD0D30el97/PKzO2GOqm6BW8F3
Dfl8a+6VRUQGLUHc5SDgCah8eMHFO+/frjkd609s3ptRRQ07iJJ+fpR9EbPrl48sfQKlZ5Zjv943
dubjZpBaOKsrckeMZbtOzL2eBUHNm2GF93mAdLMQ2Wbb8W6vTBY+QqSf9/ALcKFLWKbKSdwfA4ED
UkBTrGKISOuZDl5qI8x/itBKhYY5J/eNZuu+iMCzUt03J6vYIBh6F1AdzXeZtjzDfgazmJ+0nOhA
2jwjpmVKf1cKU9//Q2UW2ilqfTBEl9md1itHQdQJXx7GNZVHV9ssB46imb/x+knC4WypoO8bIhtq
76hnwebAKu87oBWr4CFBrpI8aVFvqyrPV0wi8YeKg2vmgP+Jcg/54LE2hZaSMl2ue+H9Gw1Lh9gL
/FNe/Svxpr+jE5n6y2sZJm36Dty+CuhAD2NX1EFan9jGyIgN/AJtjWOCDZL3XGpheFvcEqO4v7lz
F3WtHWGvUAwsKhPN8OMyxOkX+5FmYKonWcTWrEcy0heTtBa1BYp+pBUe38niy8iKXbAcjDTohe4x
h9HufGc7D9O9Cdwkikyn75LLXOChBVZWAUMgF4MvPEe5ZmpcDcCV7Ue/iFnp5uPViX0DSZi98hCN
MvSosv3GXDLFblhERvdKtDEO9p1r+l0JDQfgP34BXVvcWWYwJ1j7a/3demr/8JZyqBeAYZImvEBN
1V9sw6DjrwqjF/Qk+t0gMxN4VbO7qpse06Kbcdc499i6vS2M5heV5O2ogBNyN0fvd1coHn8ffYj3
3mVmmCsJU7cTq4JSDmZaFaFoqOYUh/uoCnKEcOCbREe9DzBnmUtQuRVfSwYfE3WsgaepFMj96e0p
JP14ZUPkqGrS39AKrVNT8oCC9PSWMfQUlDdr6huGny7WNciG2ImvGOHO13xIdWY+zBL0Bo3r54UU
9emHYT9fImqsImjUz3tIcIwNDv4YAzZu7Gqv7a1hzJUZJ9igb3U13ZVjW+8JoW6dHK5n7LiVKQ9g
La9i4lf2VKXfRZKFzDecBmGYT7RDaz/uZKCQosZqLOZqMFHuUf6V0alJYJQS+oOcDW3GyiWA9Pk3
b9L7MZkcjM4AFobIEifETYsUdMIDStyv+c/7EUGfPqee6A+eOgNF7+jRhPXqsNeeZSLkyAwF2PsU
4bUPlfaefFetIkrVt2Sl5Q8rTsFdy3EOgttOEHiacUzLVJlh55o01aRRWgPxTQfYYvc9e8NKKE0a
n/1wCHqDLHbltquLgn/yhnmnj1wfudZWRpd8ie/HFUAaHzhgY2D1pIbfqe11IFzoQx34ScnxHn59
L6M/1lK8r8E656dVOsLK9W/jyaKxwpgoDmFwVrM41SW+QvJWG9Q9GvbsqZxYfvCxNcjth+fG6WTo
+MWpWrjhO17KPjoT7qERWNxLVEIErbpFHjVwN3YOKB8uCgPuy6Wg65IyftvH92MgkBwiDgKu+oqt
5TPQoTJd/TXqfIAy0P+45CYnbB37vyvEMMV1uvrepG2Dx+SiFXSUiNJRF69GpX6fVngwxnlz4Cf/
Fvr7KhO4SVV2IFQLB49yx7kz2ykWZy5CU38gZA6Xcay+NwIbDDBTMu4ZeFoOdwVXcKSLaJYUOuKT
O7RrK5t12yw2uLuu18uWhxdG6vmCmcFbgun0RqqnYxoRRCrtbvmANIKP5KMZppevkqkvLd/DJ35s
d3hP6w9qattnViQJuX550jn2TCRt0ADpayQpqzATVYJyyQ5yRrYG5setV1uBG7BWsIBvMyb0L5xw
l1Qc4EhozFYYDRtHfm4V/fFL37AKdI6FvCTuJjFEGPQpmesPY7BMhP9NHWkNm/KUDK24D5AI/1P+
VzRHbOQfYWRnC7tBv5MdXs3GXt27ZZkK1kl0nXvDVGW86GAxsqs+bZhqu4mfkT7zismWyfRvdHWF
8dFYVeMqXXEjYpmVLxj/Zh77HEEJo+gFpoix2JZLBDGuitdBmwmIUirQjg9ZWgqypRAy8RzTr4Di
ggxxb6+scn0dL9zQnjOD5gz6R0Q0PnzaOaAqDDs61DAgydZVBtrA92JkRpRqGhYVSl0p+4g1FRPd
KDSP2jyukvM7V4jtPoPAnCYODbM2B09Ui8fZOIFJfTdJudmU1KcfvzDlw+HNmovd8RzKu1MjzR2a
1wjG0Q64X99PH5DiegdTVhVaZn/TKWeIknKA7XKqyolBmz5jrvWSkKV2tPolS46bLIWnnsD7Uz9A
aqLcqGN64ptqMGQe2p8ptdCH/ayZBQon9AJ9m/UGA+ElNupQOI9HvEvSxtcjl9PUShYtJsBMbAYD
8XZUeYdSfyPkWXjOw7SSmF7fPwrHrba3vQQBmI9yNJCXdqrh0ZpTWyA1DtymkYAwuCp3jgF5szfv
rGJ/w/4l95dlW+nE/9NU36tp7W78jLstaeje6w7gegkuji3+bNLoNE2wRcTNzoQf+1CFfxVi3jm8
ucPqB1pZuVKX69+6k/qsfpvFwiy00dUuJwBcw1Lj7ILp4qU/NzzkLClL5DiaNciS8074R/nTIYIw
CyqKD9itoT+2lH/iBkgPudcUdPE32xBClsh0GccQIKaKxeUtkWCyu4o+9QUzNYbAFQhrE15k1Z7y
2ZoF65JrvAWmY4Hh/q9Laqa/UxaO61HQAjOo/vB2CsPloPXZfcuj7+wruPLXSqgLBWJ7YH1Cyqqt
TEaAyruMNzT6r/2T+tlpHKjW2yRITNSlcP7q0h47KP/CYcEyyx/3isxZG48XxLCTTPU3Gu8ivv1N
lJ7Gup4CadQushA6OcBmWk3FONpxMPAGXEPEFeeRsNQzxi4G8MGEPTg9Bd1HQ+/ZRpSA3jdi2EUO
UeU7LA8m4hJVEHROXwruzBAZou10/2Nk6+gNyv2OHzIm/WTa+cVhCFcoAttPljNN/KqT/rtG9Jft
TCGjhbVFgEyfx33W6gSEo2IdBH8Em/9rbIej4hkeFaaI9EHXz1EGY99rWe4sssZFDRqkEQ2YRPZt
O3s2ZNjcGPIY4VFJ8OYRLTW6mEaYyG4MWrEHiJRpz82coJd4KZTKnbPnm2wWjqdR/taaZUccD2P0
zL/rzxJDvQgiSq636kmGB3qYLWltYAHODqW0iwOPEhC45+pN/Ecsf/OJcJ30RUQyvt+APvc9UZ7g
Inte0OplCsn2F3gotmXAqvLVdd8o74XYbokb52LkDZSbmCGjYGuvRwJhFAm4JcaB2uRp2u7d5bDO
Wai6KKGYd+0qNobC23N2Q/4oPsnTPcs57Rvl2DcLmRD3cmwjmwsNuWsnh75dkNqE4VTPE8cd4dA2
POD75xOplqXcAycCEAa4MZWBlLU8F5wd1qjmYy0chIZDRByLRhk/i1nadxCL/1eXN6O3pqmncRHA
mzRTEHTS06RkevKTiqR4k8GzUuAKtsDmntiV0V02JUH/lozljCJ7dcj8VoBEh64E0aU4iBb0QT3z
QIQvDJRW5avO6Et5WZo2S8P6xfwkrnwKgd1ssUrxjLtURpDwTKKSkUBC0XoAPlH7FTlIdGzSEe2N
mCmnIGUxKFW/anOidaFyVkOH5h+Z6yXFGJA9CtWYClP8CZMzpdpx5zqIULZOJd4xeqMLTYDqoOWX
V4qMqUSmhbob0kAWSjnoZ1gWWMaizbnS4j5FblZF7mTbpytg5gV1WaLEk/FUjA7VuxFuJs+Je4iY
SJjJ2+9oVG9w1y2Ssvhpw8FtNQuCI1zmD9R5+Qx8JD+Bh0zpDq/B3RFLerYqMY2a0rMiQwJkxd8f
kVmSR7Z5ERfAiQoCPAKRudg9TotFpy67IQ2IiA9zbyxQhP8n2K/4UsSoSbtEvpDsEIIkSTRMsbm7
UuaAAgXiUXBb8bCdiiLToCodaegIAerna8z9coVk8zB2udtrbeUpvSTbPpUVTe4LTcA5mDGTzcd1
99gXvsj0UU+6Q4Eqi4ThchE3IfreZBCAIK+QIgasbtg1NpwPxqpI8D7OG5NSaBfLktEw/clO8s8p
NFuz3Q2wt5LzpFDlgXZZliT352nYpaxEH10Orz6wRM9iPi5l837zt7LBAkZ8FcxjzFAUNi6YvtGE
FGbaf5j3g+JcTFCRjRJlML4S7YoR0N0FERAai/wZhiXOA4NarfsS7nFuaK76R44lAjimp/4Q6ym3
/64e+K4KqPzJz8J1zCkqKr5HmJSzTeohy9Vj2MwVNwV92tZv+YRAxV6rSz7dG+etaPq8rjNo2OOY
nNqpvseM743aF7BGNlhhRm+jw9tInK0A1nZoaaJcYHcJxzSdqbeHkGa6HZRoGOolyrCgWP6wIcrr
7TmGs16v0udzvbs1E9bBckkz5cUeUrXgeHGvnVBp7xQAVMyfTBRgtICx/WcPLSFL6TvOEaM3gaJ+
csUHZvjxCpRqdzjB+MwEzcF5DPFsAxyIK5NH5X39A1nqlWiHxMTsfb1vHxx/ccsqMBAI656SoIpj
VllPHZE+b6u1Slecv0NCwDZtBagrPePt10gFJ8LrI4/fUmEpfCUE92XlxzgVU0YBYXyNbxvg5wI8
3f/aL84XJ+iYFpztGBfD+XfW3nnIXC+fYV+oY0KAeRv5MICm+EOw1nOfU3NSy3ZcRLXi2rwLE+C0
LKhluGQHoBEhdAaJDius2Rm1ha94Ep+Hrycu+bKWW2du5ZHhg5lhk+JVVE39ZfFvEpNRHwhFub6d
lYaIQXwZ7Y2wcb51FE5MA3HX9Y60dZu+n7RrVfTQceEGcjZrkqZNv1OYi7ZkD+7HBkINWrVE16hb
9PqdKFyC6veexlrJ2Sl4rAYAcPNZGvM4JAGHCNVp5rhw+Ubaj34zGAQRRUZYHwK2QAAQyNvref4b
vitHV02+ZeirK5pJJIHiZwpQkPKJs0Yh144SFWfH4WBsbdVOQMxxcb+BmXb1hbIbIpMG8qEGvZJ3
WDmgraqqNu+1axi26EP1TUAMCflveQq72cTWX0BgEJ1pfmtpy4V++YlgvmI79B2dN/ktWiQHc52e
W93KsD13nSJc3LI1/yQVkBqNOtf7z9KQJmqnO5hIcQb9grjBIsVyzSODAmzW7ShEwgychI0vIKQk
roFJTElrNbgmIpLJIIoTwfHR1tmUD94pMprfmPvu83mNK+tFbVvsRqB2FxCxGtuFJZmJFHOvgmJt
Yft/POtusmhW2U2qUHkXId/HufZAE3GrJJ9larZ6YpvT+MKmAmnVp5auKXPMIvJRrohvF6+FY+Et
v3yS6guG9wa2aqgypQDOnuqNe7eaj6M4bO33Bd+KSdhYYg5ws//LkNZuIgzI2ckE1rkQ8atEsrbd
GKWvKESTom5XPcKiB0nHZNOU8dDjms7ijpNFE/JbchMqxbKXh+0I52WvsdXFWtwnvtGYuTZt8uI0
ljN6wSTEBo9fJdDQVBvFokOKkzs6nu3c8hQGIeJ2v2Abkp4FVUgGGrp4K4l6K5AasqM2UIqQuTAV
UoR0M2LMESVxfbDYig94YDG+1SOQ8mb5LpJrQZnYcwdIb+DFLqtlu2k+ATFL2y5K5AAi/V3VilzZ
17yJxhhVtMvl79OHA8KTbGwjKF+yjrwqgNnmfy+YVX3YE7PVDNAG7CMABYnAIo9Ckvk8pxaV8yjB
sYGl9i4lw9uxi7JFo2QKxwHrgdQy4NyQ30RKvtcEPqSyY82nPo69J43dZhGn85Qw6mLWRCIVK7IZ
GGc63lRkeOrJqRL2TeXieagyVPYzwdylwZL4cFgcRhsV7Vfs7l0HYke8KeTFmn6T0JjPkdsIbv8o
6vBqsgviuJzKAQgNkvrXqrX+zj7e31DCb+dIxmWSnC+QdBcuhY/YUpHLJUnXG8edPW2mETxGSz2u
FH+8/Ccpgq887WPf3w25YlRcazrT1KSBaP7kww/+wXtJkC8ivBqvh6lA4TaOOTDYmii9tznex/AT
2N5MCbG1qlqxcWXAR77+bZcZAmXr7Oz9u+eeaP8R9b10L3QK2dmeVTRjXofRWcfgs3+WaKA1v/wh
2Vdq1RCCNbv4GMPwmLyNhkMk498ybEmYvPwa3AKUlcLXN5keJ5vWdCSQN32HtFA8wnblzBIcQUZX
p6/tiCOJ9LiGBmv6PHr/1ezzYgHq3XUfVYDKEWbcEKAeEvb3nQAFxZJz4nMuAsTVnphH/csUoz6d
7djl82LlO+emVrOZKr07+FuYVGKF3JWM8NPgR2Qtg4WcwADsML1bS7nS6lMxy9h4FkmSHiAD5qly
AL1xjmsdvkID5T6chOZn6qeFVmxcZovXQcDcuQFAiCDJoBD4JLE2qS43KGa3rJ2JejmNf9rh1+0a
auG18ZyXoka7vBsYXJoQbShwRZtA8yBpSlrMLKz9n8A8BkH1+8Og1TIspMoZ1ZNkl9X0xx0M2nS+
rifmwzFI0fCJ3vmjd/g/U2s0QnAbDpM9C5t++kGQAUHZZnY4mRFD8A6hTS8M8Tpif1pxMULLSWJw
qj/Zry1WVMwenu0l1/1tfrYzHt/GX6GvTAAHeP+jbmvftG5009JSRDZ/KAa6kkeiraq2h9Tfolpu
BIiZv0/5NLiWAmBCdOMfjfOeoY1yygNZ4MbSMxpgLFa5oa9zFD8hbWG0aBPWoPJOFLzjgT5bW3X6
zKOdN3BVWNA29PTjc7Hs1bTKlRWAtvBeDx/fzSdr5Yh8DOCZpho88oow1fGLXaBZj7vTcGPC2z4t
mGnGPa9u3s15i4UgIfJP8HPQPjaAQubk/beyEQbO6f1Jmqnf3kQv4EcnBsLixGo1T8aP6iVvt1pG
F3OCMHWNSd+yp2E8VhoYFb8PQovCCfWlynEU5kPgm52dTi+or/Z/D5GPYWvl2OqnUmPUbPA5+QdF
Qr8F/uJ1WgkQ+98kDjK2n4uYncNkHlyqzxz2LuQoBUpTNMo5zlVci25D+JrgDoq3nzELqWwj3vCJ
7P+Axmy8J+XqslJ0pOduk+WV1jFfxRfHYtM3m4QJs0N30LtVgyc6t6RosAeIInoyoR/tMEJuKAQu
/mtRczQZenunCGCOFi85HJ/dpN9iPVf2FEjwe6d+HaOqFdifG9iORuPwriFwgNbaPbt7IsjcgZ1o
vPNLqYGsSIl4Lh7wG47BE5gBJOKSPk5qmnz4WLhDjEPv9XtuFcpQNDEnlP9XdyYQKtzxFKTn1DRP
1lUSJQaLKerzcl17iOKGd2ne9L/hkYzjdTYCGK0fFSP3rqcavdB+AJUi13HadxhiO7BO/KPnL3CY
Ju28D4O1G6VteMlliJnEujIahTr38pc9e907QfUhjq/NCjz0H4Hek/GA/i4CTczk/aFhRV+67Rwb
YJCxZ/V5UGIGXy9rFHgiDhJNfHzLVhNwzc5a1fKxvBHIChBdbtOPirN1dj8SZvzYpCoXRXLILWRL
aHTc1gZ3bIjaFpQL0+WQ5508WUDWBFuioZV7dV7h77khLw7tNaq8PWV0WFDismeL1WQdSRNb3aIu
Ary4TBwCj45i27xqF0XR6W60Bowu42JUe5Fd0HOd3sJIO+rgmJBxFhwb1TZUbDRH1F/LG3eeMdVj
MVr0H2ivmazDUnotGO7lRGWw6i/oQ8ODDknROkGEt6wo67fvskWbb/5oav8JP6GkXw/iFDAA7r7B
7JSnWILc/eLXk/3SRyGmyeJ4TIqc98QAp0nPLfAtgUWbPGuiYpIF09EnzjF9Nnpv0R+GFbzPJG+J
4/iMT8qEU/b4tmWPqmbxQEcMJTEMi7q69me19zZFB+zWY5u4+hX5sMxtwfiHZPldFvZkMqntRnp7
u5KhPe/fSeLLG0db4ueI7njmGHdzvU3kr+Q9EbFLmZfpO5HfC+wZ4knD+4NGMQh4VYhDS8Ei0FGI
jTU4DruDAz2a9lb/JLFb5yc6uPn/shvYt133MhT+gPJXGYD3gkp3+124+a3lKPFU0e05I2R4C7bL
hLWX/vnDIn/ntX3iV+OArI5XTbiPVKR+fjEd/6dGQv5JWt0nHB/gK0qrb0iKcx8l0+oNXvUx6iYC
9ckJTFXG0Satp/vS5R2TRdu/gfVJpqCuw1Inm8BtZbJ/rYxnOQOQt3pc8xjwhHHwwN7EBaxLQU0d
KH6EKVZBCaw+PHQI2uPbuB9L++UeRczeUm/Th2BVkpvIhD1esQH2rXrFL4+25YJC7QgDg+bDT4pq
1IdbVVrfwPPDS8PIQhtsFLbHKvKbfFkZGLG/ykDPtXQL7XOOpKMpiY8bqfBTg7VIHB30kaOvrrgu
fh/dm9SWTtMvMYEHUyX+0Z8GQLLz+yOSKCE0OQ/lHxrWMeoWylPgoNoVYNphUywF6bKFP1SJlLe2
UbnqQzVGaNbsHHsEhX8zTlfUYYLAkw5+UFnWRvFpxJ9gP2OxtEYT8tRnLaN3xifGnWB51beJG0R4
9zdmS3akejGLwWMyKIngOk/TZlm2wnihNj3QrCRevBZUveHHd7xjpcHCnBMFHjPYfyzGKX5Eo9cX
Jj3voEg8yf0jDX4SEiVH6ONz2jb4Xw/Icy0WcCIqYtzRHiGSDzfuUSxkeB27z4KBpiBxivtWsod4
4DWFURRMqCkaxDKz6nHZOwWHW9YeYEEl8vSooNVeZYRIagcy/8GNVW/oHOqwYdLi0uyUsCkYuCbq
IwGqdpCKV5+E0baaQm4o5r26QQ4UXVQURdAWp64lLASrnxJKBpdq2XwQRA6rdUCZyjPHV7pw0Mdp
WNLgcThJwTaHQ2fnqWOp+x6QFBEcf9xMYa7FswU/1ijgvS7O9RzhYaQO2ZAumBCP3J4ZqoHI16M9
xwSGoL27gXEhfSUgBL2Giv6psxEHcM0YXcRIXRKHft6xghbLoSfjljjwMzTnE52YEwS2oUazHlhf
OjJRm9u91zz08M0CSca5Bj2wpvcPZAWa5XCsaAvACZ8YpErIJkv2dvmjcRWMgNR5l3lkkPBJxtkH
EeSUzpjhUMGRinoeAeqeTDlglLBPeYa5Hv11qos0TlsWNaHAPUWe3huu3OvORBxQW3FMtUZMkEug
Nb6NUbqFBNb3IWYuPshAe/NXVjsGKwwPe/jhisDav2QXz//Ufkhg/cKu0wRPIp6Sr+mhpvXsarI3
WfF3hBG4R18Bd9/JZQDUd8UkoyoabVXJexBWSAJbwuMa54/YrLarzmjtBNeqVuukMczBqk5F1/in
wH8LYoJSEngf5qn3r0/TrTtDSijVMJm4GyRuq9wdOeozOdBu7wpwT6Jq7tBX7gOkz+OrpV0M5ETY
1pvJKr1gjFNvY8llsQJGCefOIwOHWMEfOVe+LCuoWqrTUWgzGI6loj9SNCSMpFLAI4SuGluiwRPj
3snHQo6tDP3PLq3S4wrFGLPTXwtbI+kvtD3/iHFShJJSwos6AF58V0iMIkqpfouCc3oRQgO1ZOlc
yEHNGHQDTE43rXdYKpXXbaANR3Pn7BUFB0qS/8zDwka89XiAUHp7XU/wqU8ApxOWD61LHc4MR4n7
wK8e/bnh4fk3GdX1+ygtak2GgRkxt4eAYk9cp4BCKVG3z5gFQEQ2kUB1db6QxC2g3oNGE+Jouyr4
7v+EDDgBu0G8qkbJNNh6zWtmteRuejRJg4aBYcuE41pYPh24XoyfhcUM1iSXZ0X/W+h9OhIxkNxZ
QaUpNW663BtZC4rBrYT30h1DY07XGGqgD9oq35aKlLalzwnAe/Mg6FnxBN0i1LtwWq5sO4sncAiP
0NflJra3uYOhPRIjFEGIF/tq+DBEtyEjHI1R1qjdzy4O5FxDBZrej89+43QD4uS3sg3iiic8w3ab
4Ayevw3pitovPGbM5sIuJr6HVXh1QOQ89+E9Ah6YKfMSv4RCKU+wfpyocPsv1f9IfIHnjZecyuTW
vSQu8mEE4xDvG2rRWiCIRCRM9PW4L7zLk1NeyZCI1vc0kwsvrOuemfjOY4cMynEpC9q1uhTTlYCz
NZN9Dey0/9GmvKru1xyIRMjno1u93MXvEqGxXvCc5k10S2PbB8IIIet2iYGh6MZIQLGNoJ7qPx4K
AbcHnotb3IrwinAifmsDlSmFWIfsYREbZt0+UcSIObVLrWEEzAu9VgHipCI3a1dUCKUKcTgJu+0f
BQyfOwC4D2Rk8TSmyNlyIAPf0NxM+OScTMWw5nwb2sCHthBRL8pZZPF/n67e7qMjeamZ+pPw7Cfb
SfteTI02o5HHnHttNpvRuBEvN3PQzAx+MIBD8aNlOeFLy4d667BaegWLKuaIlu6Sjuo6uJmTRv8p
wV0muReLzCD9At2+DuobZnZOSLBrVnswo0RgPpQ9tdrcQoX0PZysPql54XkkYHJeCbg1wQpvawSS
3eNJZ0uW/b7ce8b1y7xUBIiYtVNMEdsBV+0OBq7ApzG0440V+l0+6wloswYItmQIGjRYVdt9hQ+w
o17v9NX0ua0HwmTYvnD6gLSCOfUjqyAvfRLthLnmwpZmydF+JB71FEBqabEMlNdKek4Rtd4baVsa
1h+omyl2TXlMSoEepW7p5vnwHFjZpzUEkvCrgr814iTXdfT1Zd0aGtit73nOVmgQVpRaD78akR04
qY5/oOeZMlMpZ+sHMRkKl8sC4D9q3t7cxOscxcx1G/MCT6C56gpYwibUf/wmz5uxOH1UnWyA1gVn
5JpzR4pbfuIcPd/QZkPYzo41E1FlPcP252ZslysNNgoGAzbrz3zTnWYTFuBQBFckmALBzxYKdA7+
pMAtRA7atT7bnLu2KVGi3FiUSaYo74Pf+fvpGw4CtpsBcE6os4G0q6DjDLWWJinY1CWxwoCCLpx0
6WbFjlqCWHGnLM9dn0tHlUapqDWVvF4wnYMptjVpU2sP+o8dZjq9dDnrKoqr1TYR8d5MfzuaMMPg
rlEySsoDhUdrRM0Ng4UwezgEBBgocRrkhDxGcZnGzTjqaeV7K9jt8dN857A52a30gVntk6MVSFtF
+OSjFTTTIKhbIceK0BITUoKO1IgJKAa1aJYn6fguqH8E6krxOcgoWCB2VWGEMLxE6VV/1D8FkRn3
67K36bZwq/TvhsfBJ1CPnhFChnMSIf6aFoYTBUhhhX+KfnT2c3DlhbffQw3pauSX0r2fIOr/V5uW
Yy+tZ8Uk4UgCzQOVNqCfMc0p5jHVF+Hr4XU/5uTHBYcy1o4AaghxZ/HzyNWOZFnUM68YPDZdAWDk
kCDWgmN5YYXTzj9DM+ako3stf73ZiSbOa2Lq8wyllD4T0F9K9CGx943peOV8qoSchDMXGM67z4/a
Abm8oXLSD0+Sb0pm5+ukfBye7/IoAhfVIut6MLvQKAtBccMpso+vgB+LfMh/Y7bSztmkLSR0es7K
SDE3k2oPmmR7CgQzRJetjZMXb/YL//I4acZt+5Mua1xcOhCYPxZchjpPJa2ZFb7zHgvnU3NR3Lkz
zka+0JD7xG2CNuFW1FfHjS4yRXMCGnl5032smc5vPALVLOUFIBMjl0ijVBo+f5I7SfErrvJR3OpX
eaPY6xSGLYgDKPf21hwmYPxDHx0NtoNhoUnBnicjK0EFJPAn+uGrlA+eTWDZXqDXgN2iCqv9VdgK
OnHuXEzetNw9LmPwgfROm6mXVzIbh+nZSN6JiC9R0UA/Eh3hsDMMzIAjaMdgGRhQlZMJt5H6hGhZ
k70TGEKK5Vv9l7MpwVuarR84RJ+aamRBEHAoprgxzgoTw0YqiYBqgLXO99hJRXX47So7LgA6NCjI
J+oUIzVjknAXUs7j+O2qajnML7UqnFPJ9nAwf4V9CxzF2HQ/SqG03E2eV5NFkSJLawwATUhx5X8h
2kJTjTBqMrknIbnw0MdhPHpJGCWKdGRtcG34urk8Q/TLcp5Bk1cO8BLh14EILb/Mh6zE6W81bnLw
yZnuBxNH+F7KhinCsk+H7LNKZsWVr4WwHim1DsCnuXITGGfVfm2qevEx01LPLjb7pfkcMV0PiWGi
e5yAGjvqGk4Wg0roCFkf7R9auXWvlpFlyIRiyjcqHTSLD0TrA23K02Vje88JeH708YSxqP2mvOSK
yrdVtAw/DdC2r/UaqkAyNy/MeCmQwt3LSj7pcjQIKsGpYoUCuiUJ4Iqfys6xz4/qtPkuXl0BeXBH
iZRQ6UYRjf924HnvbBQO2YiztA89Da4UQ1CDVMDznhkCw6XLrl/Z3F0aJptr5Rqg1taBorIRfIFd
jWUUXAI4x3O4HdI2mdOiTrGq8cenJjZuSID92Rqtbu1ZbrTGKYIhjWA665vy/QRzKhst+ZNZpCF9
12yx5drB3WSHwxISmDB4xKCLiscFWu1IxrIN/SP0U6hxcCdfisCMyAYxP/76+tCrW2ofUDWDjEbm
Yp9Zfk9MzsSw6sItiOZClgzuop9UrYr/9rZ9pzwQ+Pcz/iem6k0mCEznYGpo6sVNYCj9oxt1tIM2
nmZfoa/EB6EFgwRpd0ooASa+xOdOAJEDhQlXKGHlK//lBn//F6FL27gIy3G58OL+maL1DyjkUrnk
y/Uo6mPzrm4ul9NOJWeWzS6VDQZLqmssA/FnLrli/UFnBXnQ2ZHJZrMfArZmY7PngLsFIT7gRT1b
PusK9Jc7rFcMa5d0UjqDb5bHhXURmXHawu7Zb9+IiPmp2PfcdIpWw3S9QOjIpCVgkfxIAL8kQS7m
nhYZHTRDXwLKNYuqpipjlR2dx2wjLJ2qJV6kTrTFLW/Vcwh5JABwogJQzPQ/CXl1CUEOy/KusQY0
gCWcfMQNqzgFXlElDc25/Pn/buiNIaIeATeuD4p0dyspUyLT7WTbc13AGvjVOMXm3phEZr+HVSdR
5VW1XNM5UYTvIMihnNGzdwHu4lqyYEUGR+0GAWOvSScDEEBONeUXlM/BXnJf503V0WW0FgMs5QlN
Xb2pXC1C9n7PQLkhJLd/C4AfVrpBoMNLthedzqZk1cqnkjNfI4oYRAu2IOA0NY5k/NCN6QonUf+W
oik6KIZTPXF7C9Y5RmppXyFtjhpy+JyfDyEneH9XxACjudC1WHdlTdhNbMHBB1ZaYRwPJrfAfcpn
uP6Kea4KIGXWaO/FHCl1cSUpfliGcSD4bHQnijz+gQeESqQOvy7s+G7u4REDfOmFZFmaPTpgxzuh
yu0QNj91ZjVmZYbntlAAJAd6drLV1CH5CwpdI4CfdzbWQjjt7C1AAH8dRabsgPhHchJYMp+E32Tb
GtTcEq7TM/h3MVxdTucJerFgtgIgBWsAlyuDYtPSrGg5RJBLt+n+uSCHya+qEzo9Ru3c5c48YE8T
1hBJZQLx8yRIJocHI9ck22A++bNmnEE3FYIeXbgnM0NhJwB6lOP5nhdIqJgjqYXZLEOFRPSWjUza
zhkQjvo27tfrPAJFy7OkEN157/0kTXdcwpS8DdPpo11KpNSQakJuLtHMhMB9ndpNbSA2d4Fh06Ja
6aHApMOzzklOZE4zPM1BdtQpGN1PXANZtEmNTc5yDovv+pCjvUAewL0dfM2b7jwHgzZa3LW7KWq7
B3if4tRzX214KY0ln+0s8pQmuB5dp5aUaupPp4ZJz+Prl3UQyp16qAArg+pf0zGK1z2Ozj3Y0jf8
+ms4Nn6Ut02zd1Uu0Xm1/5//p/xSuPvagWLMnIHEMVX5H2RJ9X1Xy8CGGz4PF22ftL3oj+tuzNEH
DDXX73A1Fu9jodJVZub1RBY8dS4olgMNNCoJQlgBeA7ylAMLSTqV7/R3OxauQeLmOvgFiqtxa7id
Zd5H6L3bEBY85wPPDbqzSDN8dAA5I41kj7xIWoW4NE5W1iNggirREOCLOsWmS7jHlVgqecdrJbLE
N7u0QrWwFKIgQ4VkTWm9EaySANePbf4EQVamY3909h1Hx9vSt1V04JqM8eveseZfSZywuuGk/AMV
ns9CpBzwLnD7n2krU1GpklCgTEo7JW10VNr5kz2h/HYyzVJ5z5ajCPilxXwpPNOhn0VOZVFnE3wV
CoiGH/ukvlgw013GIiLaoZDEHna3+15v3aPuzGRGhjsclJew+FztmcG57InjfYljHFYAhfvXxclf
IguVKi+EyzIP99mfZinC25Q9jTOwEW2w6fI02pGrIU8jiODG0HM2vKWz442hGgHG6GVnx1yVurnD
iuwRicy0+LdHhwrnvEofR7LnjJT+EmZdctPnUF8KSaLzhaYZuV+MjmGwZNhs9/Ivy1R1JKgh9qL8
2UowYuTHHhejCYyvRRJJtaXFumIcDYoSEDZxhAJl3rWObAFVDRvU4J3All1Ac7J/tJT9uand5vwb
NpQPRo88dUb+6MsvwpcrL6wERAhLzFyOD/SzuYq4QrL8yQ7qMR/iDDq9vk0XhqczpZ1NY4PQvvYD
a4+AM/3eKRHrwOpH86UI2e/CAHoVz//sNI8hN+D8DUIZr9yhNW2zmYfBUn9L/XUq6/4d/VjuGr4W
d/N31HfLuuWkTMXO7kfcJpXrn2TAEl0QsGQ4OSw/aw300u+Qsn7zlblPBBkLN6sp8xoLqS/xnK8/
W0yllrZiz2QZGQLgimprHqpoMIzqfDy7YO6Q1ZZuGgIMQqwugXcuHlB2W6baRAVmMYUvQnvWggia
6FkbEiiJdMN719FhV4EMpdkp9RCc5UVyEX22s7hcuFt57Lu9eN/UTU7YoX6JGADnIM7uw+LNz4H6
Z/Ua1fG2P2g8hhWEBdIi/NmiPAzFR6WHo/dTQLRCRmsxXr+Lc/raba2xQGaSPJ/E5b8an1L7gryF
OyKBigVmjUXLiESyaoV5FPfFjU225PZ+ygq2q+IFnD9Ct/wsoNuQDia+TAPz/db+zJTyGKfF46zm
dMTrS7/wCSD0Wvnv4uuj4hrjx6qofgRyeaWSI4n+h2wJlrP7B1lwSoIH/7Pxu02EOEWS9ZKF4F8r
VsAucyWRSDWh6FL9K1DYwL18mbt7UEdo325yWoli5z6wKOKgQv4sCVKa/9rb2UxYxu/2Q0yjGaud
KokeoZbYkbxGXd1oC/ONv2rqOoLWtUv+ObC9HKA2Vh5eSxqUq6cktrHyR2ilVOv9HjiQ8xlFd0mX
teEAtd8fEknUMeZy03hsNc21BZzLTShHOiuNVpu5VPH2+H0xxibuXvgl2fGTH6dOsYWT8fl5Gg2n
eYUDYW7qWj9EPJmq337UYJ+33fCHm2rqpHWP25ELE/PQQUima54tnXULM8QepvNCNzrZHTwdsrmX
cG5D9MyGgbcGBl6aqvJJBwbI+cXzxIIe3wPREy6bGhC53YEFDkfBpeew20DWhRtCvNdJC8cFFisB
Nd3ePTzQsOR/FtmcU6mG0mmmntx96MsvPvzsb4OB9Dc3kWQZS809wpwGsyrAkv6dts98vGqQTRZc
AGW9XbQoAv2rQ45/cWi/fZ5Ty6BDR5oEVyNwS8FsF1YmX89ArKgjAXi5aW2vndV4IMh+rKWehmky
E7T3j1QjqNz4sC6s1JnEXZbUB7EC6VwAXb8DyaGqAQp6bLgJuvDKsusAQgtEaTW7+XctraxFlKje
Q9Xs40B3BfV2pxXgkHAMHQzYcRk72K3UlMW79sds3fFeYJeCMVj24vUYOLyGUtvFr0E6xOsq04UG
JbtGWGvS+yBrHLnlwx4Yu+Bfay+ilGZRdpGV0mPqvzzPNTiwuFCwEMR9/gBulHXYOcbZRE1XpLUN
nWyB3+WwoAoiajHa/qgCTWvLQVk15uCo4ClT+rQfhHYZqTq9VPBoWB6esbQL5lGEYO1vYkRtJQmF
2aoE+5vH3qW+ZebUu+RZyaV12FyjZxchT9NRgkLZjqfwHpOL7Q8PqMo/XRFv+xSoYE7keLZDC2zs
hEizHHSyCP2J4eO1Hch9m94jwj5qAlAbQ5gxpJrHxWJrUvbtiHavAdkvp+YgaS7RrrdWzZ14nhG8
wxBKdT2snKcRNj5xEM/WtvO8LDvqS8j+lI/AgBdWsruFKF9Jr7m5I+OIgAOi5gswRUFVFCQAKmtP
qEtqXnMFNl89mXVEPVV7Jevc/axX6xaMFxDtgK3E1Io0jWpm78O9Ozlb5MV7PK4DwpKBKLSv+Kdt
WIj0U3O17vMjbnsw3mef289lBEClFvLIlAIujgvKHLyrLWrfWx1m12ECXr5Hkyml5xnKuS9cklKs
IIhH4zv9bRR2QJw06iq6ZLI2QYe6EnF9GZBd0Wn7C51L+nT9mIJOCo4HHtdVLdRknlGwD7CGAwj3
Trl5MQNwmloQOUveskp1/poE/AaEV5JqTIr9NJzLSa05ErzXQWQv+S9h/MC98Dtms88lsIUXZf9s
Wc6b5DQGuJJU8j+5LRTzyq57APJcuxIWdu+O6JnOJkvxbVihP0af9yCXfPK7VKE7t+TYcTPH5AOl
9BYFu94+mCX5kqmHHgwemGQleF8D5VUccYHWZzv1+oGnYYgGso6RpWeg41CiGstQ2Ia+VLsGTJvA
lv9byVtulXgDfPNMf6ddDpp8u5No30klZHZtGBxTBP0QfAe5+kLPhy+5GT2FpPIGIJkUH/eoz4Uw
41I69Sm48K2wH21wbVjtwn4HCOZpa+wNOHuUhYFqWxrf64y3c+vl4htrOl+xKWkPxDN25e4Ocz4u
p5J039XGmT6kWZHw1/N4doQKxz5UfquFZjSgUa8hrR5vSMNOTAFAfcuDRJNMGkaWnLfyl8vdKbfU
lqT/JrY14SRPoXE+mtAkJhKsdhv6KMDXKQgE4H9G3+oQAH6LnR7Jwu2jzo8epyxzmi1aVhfGwlKW
I8XxmLtbf6WMc0YDb7bJeiELLhzvCLhCFIDalrMvoMnoOQhLRNob9ZRRczGihskWvA/iUFOp92XB
vqy9w7WEqZTdrMfe7Ef74rJZwWcAkiUYHV3E9nUQvT3iJjzjd62dndeEJQgRK/uA33zB/gTDLuiH
pwYg+4Lnh4uQHXgNsXrfFpeJH88befRh3LX930D+5p8posX1INyz68FpqdWZF4dBY0JT9Z8+UQSa
vs51yelcTUJ6JkNY47g4JcBYh6e6jaRsZ0jK4GNSc2CUDBjfN5G5FUXnZC8iT9wOORm38EEC+Rwn
qqUU81vngVu3yZqHA5UQAgvBvBQTCdYYcOjQ5gVa0KUONO66yHmMcSuh5xucGF06VGR+1cuydcZz
6U8o55cEiTReEpgOAHs4GHpT/Ays/9OrVYorcAljdbpRJvviBExRh7e0k8zMsIKjbpONixUhfS7Y
vHs8lrID2/nDBKaq2pv9cjQMse61+YdaXtmUovWSa/vUeeBUNATVqqm7dXI7lEE8fc2MOEAUgoqd
RBuGTogH0cqVbgrbxbDhW83k9OZiFsU6ObHVdP1KuVMiqaiqzRTfTFwAlOKDRczz6ZAUsWxAuw8T
p7Iyh9PcAdAejPGIoFmVOg4+VWWGaGR3P/VLrVLZBQTHLZZpHcABVD1zcvp6b5VY1BhCvBRNEch8
XoVYP+oMbBcQ9JD2yLhArh1dsIMWuJPYXTadSnQkpSt9X9nWRAKb46cFh8WMsvY1fhkDlFHBu+IG
xSPXXARPb/cISdaTeKHntkYnS+p9mn6podLgTgQkXDruAyQs0rQg0Tje9fJRw8ItZViuYUaEZpR7
29moHDAegAK5mo1vcs8vn1Ndz4K7JfBL6AjUePJE02uc4IET5Y3LwRpbhSYrC6jKIUZADfOztpVc
DiqN/6Jhum7eJUuLfPF9ZxUrV5FRdTm+ZGrFt9jQBa0c05Th2llw/y2sxlPVXyWWWrfyf2xpAroe
joGFENNA03e0EGwYkZPLTdLILTo+Nc/zA8D+gYjqtnCmAVYuCfJvECf/GEWEU65Vssn11IxNRK4w
d9/IH8dhO4GqFL+e9a/+Tv5PueJMjY7xW/Pjocyb6bI+h1VjmiURH1uP0+FlOrQub2pZje61wa6u
/JUsOuTfYfUse4fS7srXmUfI4BGiLXhssDkP3Clf613WqS4UKPRH8xXxtB308d/aqpWtthRGkAOu
OzW+l74oGojiRt6owYHNFpejhE35gxlZ5QEe1zs0hvrdC4ZJ6R8EpWHot509oeQFZOCEt2+zCt4p
23xd4sE2Hfl2mcvr1ObGuXTD+V8XzhosehLTYp2r8/eceVeBEkwh1yKu45kiCF4dxKwkUOevGSeu
d5QLk4N1AuHGy5h17NL1dANFEvZCfCKXtUGRMbMlUK95tMWsIDnElL5KiizJhUKMhTL2JEPowmKd
4HlxWAMOsRJZW4rJdXqqWsSL3dCxwzLWvvRi2f8dsva3OFDZiSrACU+Cmp119j7ZZgX6KIYuo+5Q
JhNlb2JrsxDSvvIM8sFVqfctNswqY1RlVzbto/Umal+EK3F3YtQQE2DtPR1h4SeBiioyMr0gPn7h
1v6N6rXQbWLrSHi1RrWl9KMdJ/c53zGRvYMnuKeQ99U+wqvQduV2HujRjiXXNjAZhBMmlTBoiiUA
JhJwxV7ZXRR/rNPT1Z/+bePgSzCiN8U/rdVkndQZep2GRhlXPME+86jpUglQ0O7m/t/5G+l4MU/y
8sUDeSVJJA3PrvyLDjyAqOXjSsJ8sx2GhkWNPyFmWuMGQBtbbliEUk5A4cMLlEZ+5IPBLovf8YKh
hwj3Vk5tLeOLX1fgFFvMoGbpilxBpJjZDCFnmQHOUBuR57DkssaPvzdA3tu72363oj8o5R7VoqpZ
2oA3UxrcLCMb+Q6hA62oTdk7MelalQxjDYZjU9DWC9IqeeC6sPbyGh+/eUbMa9ZRMy0SrVjopiEF
8OJxEvDYXv4Au0d5rVT6QsJkaqiVrtaXHFKelNJiGclyGvm1u7HtSn4RqjhqwIMBtpSbIHScekRw
KgfbpkMfFm3EuMm9m2SmOVB9sff6nw0PNkSbDFrDAgGxEVHzqc2chfXpfrSU3i0r76Ky8CR0izag
PC583Eenk9qf3CYwG3eeRYq0TvOYzEMkFK6bnqMqXzSwPgQ5dsT4PDHOD1s2hShqclOc/Cn9XXbz
QOlV7jgP5tb60YU8CHmNCPQIoNbWrmU0WnIS+XAG3XNitJh41kggGQ0CvStiqDrpBbUkLlbvMDIT
x2H9ZSBNmEW8Djlo+uvGIEAtaKOB0WSxQC6CqafUbtjYvwojcGoyRHwt/F+baJ1xSGO8rP+1/Eny
bv2T4rL0uEEyrNOyG8sMqg+DzPKYdMTbq3nwh38ct3d5R2bFHbca1kE0nehFiIfq0H8mpgrsvZib
j7iwzYp5ow1GfU6MSnjx0Ni1IDpI75e+59OvKT28owB2zdRnBYOdtDmsL3GUhY4NBcIJyftqgaiX
+VKpdDm2a0dEaXzTqVpnqxbTZmjk8ajSGibV+86FoVayR1YFUiCZA7le5hZJ6TAGsQHelz0SL/0e
AySg65puZz3fNin67P4Av60BQPHQodC+H5IC6ZbBTUhlNpon+glVB3F/4lBxpXfLqkJD1NWsVzYw
fhMS1CLY+1wqlRjZWJI4WIhOXNLCDWGr84TwJYc9Jf0r3wxJsRSuR3DZAj/4qskdohTiJBHhmblf
0th3VjQMVLcbfJzAG8s852fAVzX65GksRVh6Toq4UeIx08UiarHxn4G6QhrSgnrka95Rwg2GI4Bi
xyK4oqOMBVXedHzEG2fVaC5Unc1KvJL12B/JEB1BrLKOyNE0+O+gasV5Omwt4ZeTo04oMygNOsOX
VD/SmZk9ckiBoKlqvio3cQXfNLLmqf1eLTOf5hiJ8oELWM0eaYWuYwbVJ7KATypX537a4zrBzQfB
DpLKPusAA0OO3jKrILjBiMteQ+OeTBqliWeCSeW9ZUltWrIQpMpAG+PDEtmIkuG845CRnYp8HdMw
G8DBqqe5uc0byFeGH6SlnicXy+mFIF10MdVJRf2Vaumu2vQtS/Jxg/zFCFugy7GxSRHmjowbcRMQ
LEo8oVAcjtjPOYrYoU67sEybeBnwhFACY81Q9DCxkvcsJ5yr3hrjIH57t8EelW/GaZpKQ444yyPG
nB9lReK9Uvss7YpVsZWAxQy9KLKmpsrjnf/ijXVBZsw/JTsLGOhKFSdYSTJe4K7Km12eocBwQXUh
+jwnMwiqhKIsmPCuhJQVGkmbZwBe/Yf1Ztv2u3Cg3WgXRzlCdr4YcaO7VR4OZlDVREVGu2VFHXYC
4IppI+7CHq0QUFqYKW/roBI+1H+/6toVUIpeUA9ZZNMNR5L1y4Yl5o3uAI1xaBQ3lWUCDf9VW3G5
PqsA42yhfwOXzkR+RtSFASh31IBSEJytgOIeEuOitWDkJpwnrAoq0cDc8SCwqILdln1p8C265US/
AY8y9X3kQkXvAaODT/nD4sHiwH1qRBBQVa2xevZx91aCLaJKSO7jQHQkSWqcV8UUS3vq+vjP2S+a
H0NwjNxIgP44FbT6SKHK4KJ4TQPnpoylw5UZKLxYC+7n7URl7wauRc2YSTwoRQI+ilFIF2vEGdWY
Xaam/ocqRWBvFutiFEYy+7RK4f6Zcyrb5WgFMqQx0+G2BS2/njm0lUolOZRvHF5qxlYvNhWB93ZF
4c+tnif5wxC0kPwpxNmjpkgiH/nMU28D/TGqNkRwrC8PwYNmLR67nXEzAiJm6cwoerV8UpNfM7XB
2XO11rWfEW5RWVgm5+hFsU5tc3tFnHvc77ht39Qq3zQeMSQ9b9Q6ZVYqsE6pTpUREOocAccq/XnS
lCOBpCm1jNSU8tRq1fCfCYz+6s1SobXyys1iTBt22BTJ/iN4J4FixNHBvbgVva7jThQz2lBJyK6V
D3V1NGw3uJ2eboHfY2zdPJZBRkKQkZd4KZN2Nk6k+GBPw7MkGvHPEy3VXtN4Tqg2L6MwLrVIMGVs
casfylxVa16u9NHGYaquavQeKcoHkMsQXxGs1Ezr6kyprOFtUsvCiEv8355MZFlkZbzwxrzBbtTt
450XthjucCZzOKW7SjuykmcbWgLPQwYSrZ1K9+zGNONz1rTZQA5fWucujybqENFC3OOIqXGImM50
aIEmkpb1ugCiBJ9+Rut+BzEtUUozy4rmehgMZC/dflxi0qKOOniLGiWyV8hkJZ7wf7EIZP9l8B+Y
89Y+yUnWvDYNuRKY3WEzjCpzru5Sk7OjL6Yi1mT/kRZHk/Znh7JYwFQ92CauLRKOPQNotTL0TpMX
3dLK3xF5aJAX2bfy1iM8+4LCIoX49/0kehkyVd4N1twJKPWHFJY972mYYxVs5ktxSP6A4WZVHRn/
qFgVESgqGksuZoDvW7ibdEAd9Ld6YlQiSxkXgTIZJjPrVI9NUMbokuRs+iF+wCZkRzHV2kM52SNC
kj1nmxW9u3x9D9PBt/MhOdDc1cp2496iE3eux1SVv4hE/sH2x2X0EHVZBra2YPmEOGs/UHyAyM5m
Sg+Ji0tI2ctyqYAvRWGGMzQ0oWV92lpTSMeT0Al3/UU/OoMH5Kphzao0A9vvxSi/lwESMsJnBg08
U1Gv4A+dxMvlfVWAHtlVnrypvxPX0GAmCC4rSahmoKsNxsCv0GmJbFKt78dgnxCYNWyZSQ5qYd6g
z89kScBBNzkXnO7OZM6wwRgUcRqvfPmU/hKFAvJqCQPmRVO4TFlBfqa+Wx4JTew4/vs6ZrVmeJla
VEN2/Ls5Mt7uW7CSSqahu3qy4PbRbjp8mMqmAaxyGAelHqY1EXUfjwGrwTBHsdoxnc5j8hMdJe8p
G/40wYK75Jp95PnvujWKt/kKP0UoHMCbMUP38vKhpwEFUQSRvQoVcAxb5jDXK/piKT/IsA73oif3
39nSEDf2mMnbBEJ9ejU22Ij4KZ0SceO4bIP45rlZ3vJD54ocRPRPYw6BsQraHZlvb5FD1n+havVt
BvlPq1OEAoW6e5uk7REyu+zavfa8lqN9n/o99vLj6H6FZnwqrI0uybGLqOnZoYErQ/wGrEFaJQpp
M1Mgpjd7CqA6hTYHmX06HV5vpvDltRT/9BoXDvuYSZrWkigiaA42UZqdTvC9aRJurjiGbEgE85iy
pH7QhWXcHwwrU7xXFW2/lSCSPLr6iK0vueKUezA/OcxnQvvq8js2NoMoawPVQGto+Ngmze6Jn8XD
0t1GcTYyci0TsQAIEi9dfYES6XffJdiRouDTIw2suagG6UQUYnUiuTdZxrMjYk8eso9Pt4zS9wnV
0BMSu17HoQ4rz5RXBbbbi7hIpvP4iwaWPrGaIiyXsBlbHd8g4+bYJYXXDv2DxpiBND064DWlagvu
B2NHQtl46JMj2HIUHLlfj9RNLok29U6SGRgt3PXL3byhQVuV26SLOLbFe/H+Gjv0cjYgyvAaip5/
M+txSyZ8SgDadxvJIIav9PWc4y83bnCuk+4DtC69G65VNx8jSgW24JnJ179wuQBxc0pmwiPNRQ9J
/8+cbiIehSp0of+0yAVcY8T7QSHMs5+dS2A5cvn+HcJ2kNUXb9tMpSzWI7kfSmEpOXRlJUyS3eGP
TDQBLCnF4Tk5KS61jYRJ4MVpnqKA6SPkQJWDRleivZtWgOB1xaMZpXdoomFEGqsr0HJ0B367Qw4J
UEeuKzwVTk/idrrWlU7kkriHBG3ka6bwM1+bzOyWFFiUFhzmVBzzkZ7q5NawuZ3IP7Pgl49j5/oH
HuQg2rZbVoggfIVmDycgjfhLddDBzReJ0e9vGXJB5OPDB7s/5r+GcE58YX3Szzvz6vbzMTo0GArv
k9qzucr5qGmlfqA1Xd0ug4r44z5G55sbRqh+0rQpbOzOhjRTLdnPmqczKE24aGSOhIoevWTihKus
o1e48rPMRjXQpRUhKBaEmerxpMS0niqLIN78YBJx5S1zviCuSAkQkrrnYaCkK6rQavgVSkNeAC32
AZyusgQBLNX050tbgM8aPjyo/d9qvJEMTsR5gjWEb+fI2UrhauelWPrh+L2lyXrsSAHrVHXdSS+y
Js0lFEzktdvi7q1Me1jdh2QCwjJLFRZw9UVoCL1+A+Ra9JXECm7F689iUiEeGxmt6+o+WTEVmCay
FhdTluE+q3jrkjO4puGW3U9kKsKxDC64S0X76QJcqKUzqyTv6JmhLRQ72Y/uAqK3HAICku/ldKY8
gq0JCJIACiK5zyBop2MdjroU4tQLBbHDGdl02o0AzfgBoYOm9p0x3Q3gFF3FrqEVMNN6u6/HDUp5
YSyKK6OwWI8M214RvNhJcmaP15+i9EMuHlwQrC8Xe/i8S2Ix86kkqnrgk4dY2T9C8cwX+qDXmTYf
2y3oAC7lNodNahJB1teqeedP8DS4i4jteI61qUFePYIMySFEKNVWTQaRUjEJt3RuJmtDiFXR8elv
hDNM/9XZZPXqXdpNsaIPM8swI06hbsygERsExIrz5gFsawbdohCKBZaQ9IzrFUlatMNqtsdtip7W
OCpwok4pso1drSJTn0z9ZaR7tN+3anQ46mlYAARblzCafbgHkCLtC20xszCakuaEd2zpj11S52CM
eTNQuC91g6FkdFQmbRXckT6ShEBOzkXvAdsizAlnWn41go9+Q2aaRGUsYJIOTSvtQP2qrJLQUK93
QXYSxLFjG+CUmiS97HCbPXdyseeqC7cvOOfVr3jtPDwuFoZO2dePPiTR9GOMiS19nkAzOqcaXFR5
c4nXvtnMDaeESl1F/Xdqgg9N3L/qq3KkDia+EcG9M+IRx1TtaeNUqf5K0suC1RWu/weIDzb3+3Rf
8U6DqlBWzlFgJfa6AupUi64gXHKY3cve+zanRGdqy6dYIZzkdwtXyyujlR/fGvGn+9LlTGYiQGO6
vVv7A+o5ZkAbRdyFyg3joR+9Z7qWf0JMn7TEGe093SQghm1+vDuBVhRdvLqe6ofI01wKx05QTtVW
kzlwuMQhDR6NipxyMrd5+k97Ohu8k0laldcTtwqlo9n7XdAN24aW5Yu63QlwD5kPnlRTZLL7X1gb
JT1a6ebgCdYDyTr8R5PtC84KSmXJI+CL6uEBZeLX408EllyBbbtxeTZFYFxqAIPrYHoPmdumj/AM
InYPmIpw74ldER8tDj8VB9hXRCT9hDdYMvHdWvU25YK4B8NdvfhXN2jXEMoTBi/NXiRPM0RX6kIi
erOzgRqri+YlsHMk7M8KCmzjvgnzCToXkZfQo3cDN8srQzNETSHjreBAg27CVa7maIt7wfrTUlBV
BGzpqPw3GmTguSdSPOvZPGpT6vbdOFAEoexbmSqbwisoO3n2RidADrX7lr6m5MwMVu4j82kcK4lx
SiqyOKYCCqT4FGxI31KGWD5l4bH1zQ1ClD5lna06ZEeFf7bJB+75xFJcd6HAKv1W4B3hWDMiMfmZ
wmO/kk8H5lvhBOhElPJKnn3ac/qt6M8+RBAaUhXf6m8vSkoWILPvgry5oo81urC9JkTc2v8pA/kV
Y2ySN0/a6lBOt/kzWJEOt27fjBY27CFVw0YRmS7g8QRDBHGxTVdkzuwPlVL8V+Tusgx3KUNPVxxq
L1mFAsIpC2vp9VeTQj13Am3KcX6fDvH2CjCn7pC93ZDAI0R+wwzqrLXsjPcW7YDYdlLClsVEzixP
qayzt3k5D/Ugo15niTV1bL+E/i51ZpCK/uq3Nc1LILkTX4b8zxHo3X0477Nrp8IF9Md/Hk5A4Q1b
Vsph6gz1PPZjNNIOPg8RvlQFGUveGnC5obT3FhIfwVBkvE94AA6bcMjuASULLx0xy/15cPe4SDTX
U3QZqlLYLis8CEt7pa+Gl6EQvCmDGKsuIr/rD95nh/L33DybNMH/A4ouAc+J2fhgqxC8n6xd8fdB
F8JpVK2tcGqdTUFwrPk6uEuhVEwRTOTjtgt9d9vWv7jBaXMJAbZt2zFmkRrdZrHH4WPTz0FcyDta
dI0CXUg7Si1mTfF6BL9apahjTGdvlLe8+1BhU7Q8cBODHrjnCrkLdKtCJABV/0qKIMnW5HCBM8iD
XN04gZtouMnGjUph6kGtSTBA56Pgf1jWRVWFquvsWs2+AUQJOZy2BizjQVJ6gKKGSNOO540+tu0A
VLPMXvYK77/SOQ/mvHxZaAFLu+2K0zp/s+P5c6OkkLzUoISOwoa0DlBa3ffdCzplU3KJXawS5lml
WfRY4DiMec9DPcXm+fM4Bw5zjIW9N6l+NYzsNjDgrnPvXLHS6NEIoRtqQvEMvHdmL331FeiQNgvQ
pjsAU91edYNJ8c/Z72dZlR7dhlD9NFvMtRX6wsRfP7JPSNw4uaQYoT1etDr/G03YhDyyJqcdXpnv
7kbE/ZLSuw++Lgzk9IXdNT3pbwwPTSfVCFazKBCchqQJ8d6Hwf1oFlPJVjWy+8lbs1gGyoUpXN6v
QIo49cujHqb0HVRCeIaK+2eaD2O+UjZUwfhQ5jYP87avTPOiV8l2mnRBuTCzim6q0lq/BuvaMNG5
W2yrj5sHWFC0RqTdngSg0A33vuuN35ekNJ9PN3YkhS20stjrxJ1a7RbxzKlHIIodAhwJ1hfcHikL
w7WWuha3WhIaJRPMSh59N4tTmZdFJOLahhM1kqh7ssitdXIE2DzK4SaQgOM8BPgzHfxD5Yt+ztmr
hsOeFu0QV3f/qV3ECeYn+bfiXBwBO4SdWZrgoSDkzYHA8u0w2qloAKulm6tIwq6vJ7u5E48YpMeM
jMKs3l9sEnWv2Tv1fK8LEy0dZ9lxXwGpvwTCkRxxKrBPO322rrZHxrVDFE+tafgpEeCfpqxW0PLM
gRcPWxF0/n9gD/pbKPBh1a1ql4P9TemrVgGp1yU4S4hmJORn3X9rHh5Xz6PYgZi6xg0P+MvwmsgY
R96JwFsXjub6Ad27H2DDNVeGClxVqERk06zBjUBxhv8R3G2pawJFe5G7LuvrDUEo/tr3IMXkxlUQ
RsIrk4IfoCOZyy3NT+K2TSDd3tq2LL/e3+n5El/LlwAWPiAm59sP1TY1arvPr7+11H8o9PSUgILF
H3ZRlCnqyH87oycDa1zqCxbnio6GKZzivXbqOLLlTaFje4d14+/7XekE3PH6QPmx6SXWk8fxyCxn
KMTC3vZuQ5MvGysaXOgF8c2D/TGMm+3ytwXKtoGvJYKE/uNihRW9lBgNPr599oFIdaOQAUQWPeWE
TsqS9DCVebl38dV27bR51MWWI+EFyNxg2bOxoWqWy8EQPSbVFxKAs6bappRNqvuYC/qNahDc2RIh
kiOFqG9Cqg0oJGUeKlwSy9rsOXd1mlZ5FMDl55bnK4Ha0/rphKBKuQiFoBDYsBjO/MFWf3PUPt/m
kuHa9IBqYhDtduQ/FOwRQr4SRdmEKW+QHpa1DUr5h/SlxeRI8+C3Xv320IbfmF+EET1ygKpBNJ5J
a0qoDzlzcWPHCk+uNqQ3GlcIz+LF0m1ehZReSEUSHjhgk6mMMSZVfbYVKVVCvAp/4nNwWvn5nBgk
FG4XPCAmkaSuPFNYalzJjXEZ3CHYw5oIPwg06dVHBLhCQ8MMqgK2rojy8t5I2KdwlFUcHxDb40kB
KAaJ1tPc3eemiYOW0SWrwhI9riLbUVhDlt8YOpZc6wyPFykKYZpXsPM+MfooS8JL+ExePP0hnohP
QOW7P7bYs9n9uaXv7v3auUC7BaI76cI0uT4BA1XX84b1qsoi797hDd9E4I32n/KyeN1NGcBN7VJi
BEzDNeCgJtMLLcftsbRXD9BZfsSdlVBMsvN5gIkyUQ8bzbaUn5GawsEoZgEXBSKeMQVTKtdvv/aC
LToe5IM0L6ypk5VY4OJllR0jPuDJz/itb8zKqeFDQRdz/SoDt/9jDXSVOtf5ieZAyhKLDFUV4S8g
kKVcalIb1W2OnRSJHlAFYc4J1QECLJxYHETBz9tSXW9GQLGYlniZdMHk2vOOuqfH1ltJAQp38hPc
WG8zLjanucu4om1XzqMo0ebIQmH3lecuaJFIyy45TsQb9orRrDpirfRDKg8KFNR1fh3gdTlMYT5g
sPLNdFbh+QmoxbWe/kjjWD6LsC5+uKoUCgzkql5WB1rsuXGQ4CctlhSpvEK6CDIQ1DLcKYTfB9zR
lezNGUbDrgsNgJWhMKPOmiuBs7z+IIv4izVUpAsaK4YwGgxVrtljV8KQnrBrjF/7Xw2jRO43Kq5l
kaIhcYjjKiehGmE83CoouiwRkwIkyDZ//+xHWuCS+QZrE8FUhFE9T7ogj2Kl19DDOvd2OzCetJ6c
t99D9ayCOADVvIGVdbBl7OSD7px+kjErPdJQdefavk5Xe2gI5JV9tji74790nzA1ns63+4jx9oLP
iLCDsXCeMwIJ298HfyxclmHTjZaTfNWL224WJdgMln0FXb4jyib8W0uxn6gYcDQ9rbAiP4+AqH4S
AOmtoNQQyo9x8G/d96rbuJoH3F/7NCR21jQalv7QlTOTVlk9NIDJ+hHl95U1f6i18H823/gLWetS
3PgkpZvOj/rNDuIfDi3DUo4PDx3h53ToF7dhM2nDHwNFckIm2AZ2hVI7pJlhc3Xp9qN1410ipI/X
Oe1kOgimrMdkrP/SSDhnAjjpFlp48w2ILKEDtEnSNTt1Rs3NFlih1WUVE3jXP2sPKm9uvfogM23Q
ZKgz+0T8Mo/oEtYc/utFfKYLRxCjasRU493CtKiFFuT1YIf321j5Pmv6itADhvaieFmPzUvSGuuh
AvlMPUVm9S0fEyTZProa/l/xHPXjtOSd5eKGWGD/rpMig30uFR1hNKHBVyZKRKIDysAQXw9bNTzN
D4KyieG4CRI+7gnXUn4mHJipRqtr+5mPIHyV0p5i2068Vl9b2lXU1hfOe97MB+P1Rwu7Xrnzzdxk
MlMwzLn7J3fU9v7/ccCXvTlZKyuKzIRZVFduGTI1JohOK1YmwZhonZHgJ52CoLe+KuoJafR8tpvo
KWAOAH5Ag0k84Dy7T+H9YUA+ExIx5hbtkB9fmjC6q9Gy9pF5Ew+Vrg+oOF7RfmMnP04IvNc1UfSD
xlHEI+RejqOLl08OPf6ZUMwnS+ITLdZcXUvveqAp124LSUMD3TxMkzW5uSWWEVLhf0TIwYRiPTaa
NPZ3VBBFEtVIC/BJLzJNZtLFOGb0szm3F04stArSW+uep0Jw1mG+2Ek53hyWu7Co1i6Ns19N0fqW
fjeRmTtbPCMDa+RvCyX4kjBKrHOCFiv13l8j7SLNo/KX4nZkNgjuzJbn6+m5+MtTasiDwdJ+jMsB
h0EJL3jOxfym6xB6IgtVEVbBnEHfQnYW47RzVtgV27IhuOttW1RqAZZ5uoTAfklerelbPwyhZXGL
forRjCymxk/8+wFst2yCii2SK6AwX1JtXKsstqsVKiSgaAV10gQT5yR7GMfNB+ua3FNChSr4yjM8
EpiHW65SAK4fxYs6ePHDT1/v98afT5mhGLbK7S8RmzwQw3azgw9HzS3rL7UcKeQu03Pu7olwV9z/
EQ6ZdoH8lxFQePaWxPqbFIhxrdOY12Wf06z7KZ28Mt70INdzi+P0pwYI0DKpY2MQFDq9ij0lF6Sp
iWJSg1+ORYAloGdmfyXIIPatN+/ylBMD03Sb7A5BpSFlQ3lm/cMcQQ72tSxyrLvx1ntHoGJHk6mb
GbmF3jELovIgOj0Wop75UaucEF7NjXRmG8oDHNCN6cCh7ro9mivOBwyXiSTtAYQ17cN8Pk+cYwx6
nv3cm85YdLJM6OHL1PGNfMWmVzn0APNhUeMDdHjTpI6x8rSfdZ15w6oseEhxfeHS7ntqHpbbVl2U
E3gUPs1HpwHb7eNwxEAfEkp37j5BFCsOHr+q3R/CBZa5kdRNSOJWIrXhih+B9yoDPmBVmiO03N6v
HQ+58LDkPOL/kjDuvUXlCmBCDfL5ZUmbvyZwbFFBMOpvdxr6S7oT+4DW/jR2zlbDSJwY7sdaPj3t
ensrlbZF2888qImVlegARaAfUs48t72MXqVKrLrbwp48s3UQByDjao9GDSbu0iwaijYDDyoyVAUf
bhUu7+sXqb5j5NKK3slWyeRNQ4TGu7oP6Um6f1p8Vk74EdecHqV1Kk9T1mMV+CGrYqZv5KAXYFOq
SXOsd5EQQLqjhJEUXunuWz4FcBqTrIlHQ7HmTv7w4HdELmrmFjmfJxumATpKl6Bs9YQ4SfIvEFjw
qCAaBQF5HnGtFvP1Yj8KZ5kt3FHXY/ahjzJ9h+RRt7XQ0NJMaKUMHhIQIrHLX2RRWVsxCXs9ydoF
B/1DNBwpW6QNo4DvTgacLPj1HGFUhgWZnIffvkGbcFGjNGkHpXSz0dRP8z8oUuF8NXPKnmZzg4Lc
zU2clmTA7n5G9Uzf09i0pX/S94cyMMchYvgOQPgjscE2xEjgV2ghLXs5PGAYo5/FOq6qaQnDHXKD
dYQXE1duAmxCJiEViBlxyQg3nFrVAf7O+zMcI3y9wtTSHsrRt8KUJffnjT0dEPa2iRXUHVRW9imF
krw+HCzDjhXo+wshgLw28WNkFUsyp5UvxJLmDTuTzCVSPOB+/erJUGVbIFnFWUTQ7Xa+UQMdHH1S
kiE6P54LJAypusfANZv+mNTqBaKVtiLc/BPP/8sBibJdH6rPyhqqK7mwb17MX4KJuQ7/AFIKlpJJ
W7+vsSi1WPH87WIeJcWiik+/nEo82755/irnr1xaliZ1JvdwAeIFmyTdLOazTp2WNvBT9yVKDFCH
fcBsSxjjNz/dYAdMnwe0UgtXd0rEipW7JCV3a9uTc0/Dh79xW9knw6amvZ7tPkui+RFHsHHCUlh7
FB5YP5pA6iARZk5DowlfNFIqN0Z01Fp+iurTFpy0gNdXg/Afhradk2tQg2kKPKwfsO3DldPFbVeO
OMRRtpLHtOdGquwDKoKGGdugSrF+g3XSIo1hswXZT+sFARZT8vdQZ3GCDfrcmg4HuFNBuI/kATmA
WPBzW+nWA/zwOwq9TxsttWqNZq1cSqva9XFnSQQPixwW6mP2owiOgCU3rziubfVkYBRpI6KTbg3h
Y0KmBKgtCWKe65Y1ZLvs6k1U0rD1yupNgs9vBE93fV0OMOswGZg9Dj4NzrN/AN6lLvcfvMRANBp9
M2dVjg3JWGHNNuQNAY8K3EBvQKdCQko6meUbq56AnEASCK8u/RsLKrH0xbu+pLq+Nv2rL3ZnrAER
IeYFsQGSyY4egs1gwIWfaKdrS62S7dVyzbfIfBneHxZ1ifuAl/XdnuJ1Jg5OLlLGnG6Oz5yuAmeF
J9LBz3ebJnaBX6ZHKElXyZ5pFJnetw4oUtPK6tLVwjIywLu8ArV+pdpGorM+T8koJzktQnf6El0R
J3Dq6iB07XFUgidy9co4iEnqAP58NsjpYbK+hmui/ZK6djS6Tcl1Qk2HR2NPmtbYvUwFjDqKNJ9+
HpvDQMkP7NnHHjgYR0dcI2NV5rA31psdPQhg+TFVHMl8qus0qZryn3nLTEi7iofk9cWNVqvh9UAQ
Xho+worCQXNp68WXsMRqI0yJL5rk23Ec07E59y8jIF/b8SyJbbQwjNfCyk71T4ugHC0Xhm3l9v2P
X/ZsmUssuurt+T5tGbdnghRZ+BcKCbA/GlZctWvxCoo+OsVgRLneI4z7fjt8hfWzZp4rOMKTWliE
0ElnGZJ3ZgLtRMeKnLdP3WrTGuBThltzH5sZfe4XHNDctg4S7LaQO32aVhq+uR39JglEktbo+4jP
z93nfwn4aNTsfezIM3tax+h7DXPsgjJzbVo2pReht4/UdYtkJ7pYhZU2Ca5M1a270fZ2oncmbj5c
4dglGdblVZUPOe4kruxqI9oJzXSCDSfBuPvLMRfAqvCbZoDQlOqmNTfFIifHl34mh+l4fQg62V4v
E9yU+51o3c4SjLydBYMVpO/sCPYg+F5pFX21l8VVfZHQuFuxOhrj1jEIsvKTI3p6v8kLEpHPaR2q
fVJyRMXXm4B9F6mHxjUUjszRto8UsxDKTEC6AZ2SnDIMTdeaKoYz8WmuChbpWgx0n0/6x+hWomTW
HrZKM4RPuIUy2NZ9BvAU7Kb6kjVdISJ4oY9hbnGN2CN2YtbAwvxOX8v3PvsmexjT5Jg09pDjtDa4
dabypP54jz2IDD6V38jnvJWaAyGo9tAQfwXm83rvAD/P/d5cj3ezLsnZjPx162BLyMW1k0uTm3Fa
MCosVNql7QezbzmP7pKWtNZSxHtGQTx2J1PapaFVkJnFVfzYpSj3EQS5z3NaM1TmCZMKr/XS+TUb
VyopPpyi9Yu0c/r1S2jJJJaQ8WGNw627pxIgUS/Hfvj6QO2qEy+WynMOb/W9HdENW9bmzCZKWD19
lsLGZ1WJl5cFTRE4waBiXIYMrUkjFWCAo8f3nuIUwNwCW/l0nWxFKuQKB/u9cfUWc6ImRCzScJsD
biw1XgUdYf6l4sYl0TKekR0uOWIigRR6j4bHONvXnNedndc1KUxnTL4v63cKIhhkPuhyVcE80SED
nfoB7iDi3gCuijW2m/fWt7Ccp0A7mVM/0eBdEw/OVcENEElI8dkxjDguppBDD5gJ2r3UWC1txo14
RRPeI8toU3+baa9uAVFUl9NP+r8meuZTiKM3j5NpcAH3WJ8C7ZkC1xi0zHRSXR62mn070Kqzgzrx
IkRG9RrRNWMBLFEL0KaBl5BTfmQNjoAfUOlIbdBoJ439merXAUmjVW8rAtUiTIFbXdA7kZbSpNZC
7KL/vkAtNu4KoGjStB1asXC11vF0prrRJ8MqfeD6XHi6zSxG//vtbS+c4Yk2lo4Cs6tQjVYRKypN
9SZtk/89wFSLfdCRyQs8JX5CIJ6ezl79jmMl0+Ey8ybDH73r2+HiPJYv33iAaV6bEH8ZjJWBxqiP
kIS0FlwSEm3ggs8E81q1Q3FNc4T24qlw2XmMCmLFxnqhtVDoRMCXKmMnMywjzCA0g3cjPpy2H3dw
L93bPi11eRD40zqd0e2WZNlR/+/aib4YmHtjyc3WKlZ+BAfrxbKbKwLwTkv2DxWOs+yQNzRbE5jH
PJUNhmGtT4fVIf60/+b3oS89drvU6OGSy19CZtmwrnEaMwB9nKac2fCs13q3dwNVZO34O/Onzyvh
tuxrBOtfo4CyEeZFfNV6oGw6FrD/tciZc0efcWX1x5Uk7/G2s7I8aidBG4or1rGX6LlSFfbm1BLu
nkprFDvmfMnCXU52GPVJX5hdMUqch9KG7BfX8UiNIx40u+y2Y/vmc25mSlRSPIi6gqpbB6Bd3Iw6
LCZoZzy412AoQg0jQvE0/4eTelNWcBZ0CDRhknwlYZY6GdsEr/mNsQ3U7sNI8UwV5TNCLDHO8U3v
CA/dN569a0L8BoZMWJUMk9/9uck4pz+DOS8/QwuaTnOEd5wQHeQwGWONwKZvnZEp8N61n3aN5dXQ
nXZHVqfKM51ashKJtN6k1dXDM6SZk/F7SZteLTSZlFE4va3cUNgho/HrBhzw3oy+xu2umAnEXI4K
XlVSxbINBwe9FVarczTNW/LVtQrH9+VEpL81jJgmgD3ZFfYcmwRfklPpoX5RFCUIR0xEqj6Z8zVJ
OEhbZlQIYENA2rb8WbSZSUqeSu3ZLAoaWCP5HaHB4Blh7I50MChQCJ9cleDxxTD9voENhVQP36o2
guD8NTjOxAuaZS4GJyzCan4hGL9TwrkYobFkttjBkijxdoTeG1URKBXqX6wSQRWM0pGfx1fHKlsM
zLhvWIjJ/opdJgvJBX6CsE41SPv0GbW6uyL+bL0SPdMNQGn5qQwW9pFf4RpYko/Dr4+gur5gYGX0
I1R03mwo2EmBg7xl+a9jeKscVhvlVx4H+uMlMd1Nof6Iu9M6bJsrmxVoga6ftfg9BnT6cPQOCIPE
Pt/Zpa5EwtBTBAreN8YKuIezXC+34SO2fVe3aitCSnypZnUc0r6FRBYyyJmZdqr/tse1w1Ng3y0e
AejiP96IaK5bpz5KB73kOQKN+4tEv9/ouaCcg0S9CYPxC6ehxDRd29MSYnXoM3nudEQGg2zCjgHV
rA5OhL2a2G0snFxv1NpmkWmxchi5tufAKyOycnVul0yXwe9aLl5MvkMcVVRJFHM2tqgzh5tGIpfe
hb91mnwbtfqx4Vx5SFc8wZVKsUozLdVsi7/Oher8p7CYulB2hRvvJgGIgfe6u0fV73C1vqUwiPEb
eGsc23G7JAXubSa5zWr4J7dRKWPa6GNqoJXYra/zvm+uYE5JwMWCc7tse22jKGIRYT0Ho/oqOXdE
orHXlGr/ohsf3qubJOJYYKw55De2OgprxrIoT8ceAUpqbdMjfNeJY3VGUPVFT0iN7O7/2Z7S6MYf
pXPQQGzcxXX8NPkiJ3QkVLgsfYgIqBIOaF9IWJ1KMrRBUCwe0BalkEh3UHXITX78un44UCUWPjO2
+Eo0GxQJnaVbAErTHzHXTgbCXo52h5DT+AOGq3DRNkCZW9mZZLiqkJO/OJrFb7zoPcZ0f2M5tLC1
bTZHLySZdCnk/WRyV63QokUPm4mKDCMf7W+ZjyL9yIsKTI2aFMdwOFQ+DbzORjmAIWby0TBcswx4
+ADfOYCX+W56mxB3luEVeyOOUtAz5sy18jzV9Wp7QTV+MzOUcTWiJLR34joWazojXWWFh+fSi1/I
CytkwUZjCuJ7ZCtZsE02ul/X7aT87VFtqDH0f9Ll3tGOrrdatCiSRgxbbUw6aKfmkyrpmJsGCFJ2
VpOmeMPA0LhpDPGxxW6ZrvycXfB7waeXIU3jiRB/5f+jD9itd6a3MtKE5dGO9MS1dQGBW6KAQCY+
mxHa0gcWoz1kL/YbHjJx9RIljs/jmMI/czdESD8pxWQj5Ygy5yXsIVWRMCB0a5gipgTKBxVbB8HC
7ky9PvJxzvjkxzznkxOS0gRhxhy24li93oxL+TtETnIK2u0cRO0orlCaoMBqaoLBDtAlOqCWWkXT
Ma2tRcWYkrt1knO7fWfa/D0EVq/3xhOHseXd7ZR960oHGVy2JE6mfnghs9yq6zpHGZt5r6Mm4P3C
+Q0sXrUB7eAptB5vXF7pHABcCpipw7fMGneRBCuIgQR+KShYiSYrIWW2uVIy/oP8H4AXywaxe+f1
KZvyhug2Ej6efVtnqJQNtUENJpiUb1bxvCkbL5altOT7GoMwGEOsfThuuyaTs7x3cxnUdE4szGwc
/L/kHsQMmemj6+B5OAJmgdiifRLBT7pomuVtUsoComcfDENb9tAYdYEkxcjmK+23XoFvZ52G7SEf
PZVTwpWUBxCmIVZ00xFuCfbdvPz0txILSNM5jVRcm4RmgFyPvQgXuQdnccYZjDOLFFWoXhsqajii
2cIas40wMBBJgISsNxH3RDrFuYA9nHi3mqtFczWv8dGjAXZ0dcU4T+k3ImNpWnYOVEQ9xkFvUpQB
XM9mbdnw59s9r696ZOPk9ChOPK1H6rwJXJ3Q+LmeIfXzVdEBHKSguvzjlTTtQPhBXrlqRt+YkxlZ
YZsFs3Hff0JpL42PQRG2RNO1cvklAKlMMVjStIjbVJU5/+IgaHwWvT9F6qNeRDrv96zURPpHSjKg
BdcNli2qjeCcehh6Bp+pJdc11ekgl9HaOFySH37kuz3W4RCJgsKrGYZyW8bDKette3rmWaB8j1Z4
pvRu+IM9b15Kpn7FcSNp/ufL+xnZAFJSUyrosE9473dNhGWoQNpSdcOK90bUeUt1forbP45axC94
R0V5m4iuyH+ah1lKqJgpiUMUVt+A71gjQlxLwjmnkWS2tjJUqsjfuVLvrdXdJEDf0YY4fbo8Q8Wp
TRBpy/C6OWw5KK48skkEzacXcKbx2ADTONfU7LCCNm9HlnlpkJURT1LvhDvS8VyVKa/qyhXCV/qt
S3AEpFdqt8H119BYq1KMO4QZx+UkliYbrlDHQwi21xE7mDlK931Wcyp2vKwdf2a7STSfMujWv0Kv
+IO1ap+nPZfY6q6FWxPF9FEPVGudyvjqQYYesxZWISRGp9ssF9hMgr9dAO9jkPF8pPh4GTXkPhP7
v402bESr79xXU+P2Rd6HhJnRHvt07XdwKgkbW1Y3/HP3oWFqJIF8SHcPzu9q+JeeOhDZWbUH/E0v
udw+g8hW5sBcYfTZYojA5IV03WxMPXqeDi5U60zwG9qSb1L3Q9AWzmzzmp/H+ixEXFh2XgEm7RcE
Y5jYKl4nwIocLYq9Todtcm/MMh3UMFMNyC6ezhGAUVPGCiZ89XRHVaQIAGjd+O2AXGLC+qMpLnem
hZVtZRP0HrGaSME0uw1uqWz96HEsN/jbKVMTumZRu17MmseA+jqlPrHic9s5umDG81l6VsSxWyRN
UrNi89GcY1Lg7LDqe9JxUAcM7QAOKU+uANFmKLTZ+6X2G+t1bFmksm7kkIlGAHRRPrdFyxk/39k7
KsPIzFCYWcItLE5QHChhDiCCstW5CmodG/tnrlzDtozOXI8ZxtdyFUGRtZBvRabAWJBQ8kMy2AKp
DVo5knCgFaDxHSHDx+vnWP7jfsEIiC1JZ0bZW4YJg0ltrU1uCYwORQOua2Yp2twsi5qBkhcA8fZj
2Hzk2cYg/ijaGiryoDBczAZSeSfaB0KfAFAD8PbCMJUkyRP9/12fC2CEAPeNaBB7YltKMQMWoicc
rFBjsKnF/g3voytF+ZRQJEeaMq40KxRzI+t3f4JVExbRGG67AJt88RSWFWTJ952/Io802G80sa/j
KXoXC58srnBK0Cc8cQReo7zyNYQA6IHC9IYnCljE8zro6esLaZlv+RUr4ieO6MRDrHIbSUBsHLYT
i2MdhifXr+QQ0busaF7wdSez5atb30KlPb5401uSghfwdh5To2oexMa18dvbIO/lSYmwjsjCXH1j
8mVK7L7EJwGYpwICQvAFuTvJ34JA3CW9rXiLg74UGelJJe1z/TdB2OP010fjkRgTR+AR+LsbcDY7
c+JHZ7mR0De47vq6A4T2iCuAetOwW+h3HHf4UZl7iwf6XdyEcg1zXWrTgHtfpQ9bqW//iiJnUd4m
B5w986u1zXZk6HCkq6ccDUDOjXRJ2VC9Oo8rGSzx1CIzo5wyiPvpqEch0j72f440e0WN4re+gUiS
SIW/mfdXSiGskMHoG6aoMGvUxvfxfMl9LSPZugDCKOw/eQIkPzGJ35bOpbzncOCXZC+TH/1xu4jq
EnJYmq33w+7akulVxV3PvizMbB+snG/yVzw0wgfBhizUgNvh0EyUo37b/k+GSFUgNtE9tUDkGbTl
R47odhgjeda9NokCJ7X7ljByKQkY0kVRPcVekmi2eY3t4hjWkAjo0udx73VwXwV0MippLhRpfCkX
x4Ryr6LuOr3iX8tYakHg9/rRmQEnKcJyBAsEIDD8acqQ18+BX6F+8itfLnnB4nQE3nIz2I1mTw3h
ZwCf14tbjW+A9u0v6sRt0BGG+DcwpD5TXTx4zIyE3XPEZjsFgEZo7rE9l2eMjH55eRz2UoTHRRLY
3DKxAaKNcGmgRxKmmAlhpga8AMmjxp/hR4rlLdOWzBIAKEWeCDDw7GtIvmb07u/WsONsiQcPu3h1
xcpEOfhsr6PPgsaoIo9012vDJEjNbY/qVbGBGhwJUe/St2Dqt0VQ/w4WEYoRuX9SqIc4PwdOOuXY
NOM2HpMV4F2muTRGEHplCAJ5aUEk7EJHqzQ4osMR5NzDN57CS5Wj7543So/N9toyOWA9FhseCZ+W
t1gN7VraWRTBn18whuw2X8i4TW1slz/1JmkFpFGypBPxZPqB+I335nHj8dMl+A7TOaSJpkj4ULuH
X+ATB9qmVdRyYnkN3nCHUTTtGdkYB8lUG0JWg1PStDylyY4/8QKk8yhVZPNsZTHqUKrgX+zI65G8
Oh6iuuZxQ1PozbtZwa/umHZfxRmNBeYyp2YiI8OYMHQWt3Gg6a3qMnZSumtAer5PsviV/ywoAmZG
LO5rCa7/NjMjvT+TNxdOobPBUQbm4vzEWlUhDherqFC+hiXjEiSCkIa8e5aGNa+Iv1G6SskE5cMp
3sy7H7xOH1W3BIsH51akvZbe0nwJfdJpqazmsTfExSimNnSZfAnk/AQT7mLd8SxJ7/1SCrDy5MCf
MmNAwt7QLI4NmVB2DSKCkybaqwyt0JJFciJZ9T3HVvsFr6NbHNFRbO26gvYrw3QWAR2eTJUEBo5R
wFXBQUrc8rswornsVxy2P2FdBVZ0cTd+71AIj598jRQ1CgAype7/R3wgxq6XfXfkzgjztBR8kA1u
lc0UQLiui0UkP4uTekiBKqaUyZACBdJmrlFTU4MRCV6TvyRjczq5ZGGlCe8nxRjrF8NE6C6B+fuZ
VQ+1RQ7AhKIZvDG6vWob+sACV3DIVru4Ev4y6MwXkaK+Xbd+uqeDSfdwv+YBtn/YiMwqFvUM0CxY
PJns89UR+nphyhkQuMI+uxtZazBiqqoWPzjxWaEjZKqWb2D5rB0r0PWm38Gpj/nj2L++WYWh5y7U
CTWwsfek5Eif3eBZpmRsXrYWgaGcAKzEG39hsCVa+/hOt3EN6os1Y65BkMeLnwrduLfe4zf0VOFH
9iwo0A9bK7Car9RBBKsskxSCskF5B/4p5T0Fw7UgLQxIb3V/5vt4woDUcad1Vb3a9tCZPriS1+Xw
POUPoH7BnQrZQHtrfA3VuWYuHKi2EF7cUg0HUqz1YtnLdARM8nRnbOLcRsKmMl0Lh+fotO0/Qp3y
g2NfW7S9V5FWmPbmmbXCFpt+cxfMamVfZQAHAxCMlbdvqPiP9rth6kDtnoLcgCJcH8RD2I2D7CZw
nS4dDOpmVpk3vOpxaetKf3vEsnxXbodQ03RXSjwsnjLPmsmUyEFkl/wrm1B+iRC33DBi/b4RG6LH
zbWHJKmTuH0bF3c9ndxnyvB7t87ASySmIZAPqhMr8RHUCMf84rOF/KDIQZAl1H5sd1WJ/lAmpzxS
DvBXT3TPx4i0HZtgg5yDCeYtDeL2G93nqY5s6TJp0nU7/6Quiqr10VxTTEq6MsjzRD6k+PZ4i7Uf
Mys++D/kap2HL1wxIeW2YY1WzufoW+mxyLbW59sb0wYWPA+8S0P/bH+9oohK/5ZxwboTTHdZgqIu
DNuTjOi6yFloBOUcGpC52u2q3gnd1KlALLWxWS1c4PhEff6vIerNGtg/eWIjnDzKrjC0Qv9GflxE
KfTGbkUZmlDN9Q33bgt9BbpdBBy8k6b/oVMOgpTKKyhvuY22XP0BQVw0YeCCxc9kZvXy37OddRG1
MQgLGoHq4kpWYnmmFKoLWHvJoC3kX56jSAkOl63hPCrwBXaHnj3s1rwEfiz74h49h9Thc/+X/1Qo
t+EvU2SUGSCbSSxa2o/EhLtrJo/MqVUU/QmQz4Bo7YdQdVGgqtap4pq4jatadl0Qift6bd8djrHI
0Yah/zDT6LuxbZ4zSezAu69LQuZu3lsQwIpVwI9J2pNCPU2P5n9IMUFaPemBAYi4jFm1m357Q/Ws
uvO0KwGNN2WZDgclV5pINq6ot9Z1+L05QvKTpGcCmujoeiaSbvgOU8iQW00EYd+8USq/mW2S/gXL
kLzeAYZwJ7soHCzm7BysRxS0uqfdh228p78lTt1YceeVY7GE38jT4YvQm3cFtfs3yC15aWpyEJ9r
L9EF5DuzWNZHA9WI5ptTYyiwQ6wFO5nqOV+IWGgO2CVxZAMN6YA0enRb9jFGw7JZRUV8cnyFcsmF
+IFdepRdpwwwi03GVU9/E0aHDbt5tEMwfndmFGpWmLOxZ8ZEifoG4o6Rj/3YAugVFwv2eQMpsZYL
c8AXt8u2PVBMDAtBOfLJUgZB0lsfKm7oHcKUtc6riQFWpn2iQbbZX12LYIY0wKup4bT3+Z/FTx4/
3trrDG3RX0d173ucxSAzCFYwKB5QSqD6WJzkR2eTPabKwW4L69LaoT3WnBBvTf9w8cnqjOV9Q2aP
24IL7+gVqTAkRezeOYT6Q0P6h09DVTaixLQuTdcXoGO/JcdjnUDn0BQHPlRFg+m75s9/D93ByfmN
EyHKT7kywScHN25Jdnx871B3zMJcun/vlDf7yDnCRtqgs8A+CaPOBRpGqTU3DHtYtMEjqXV7nOv3
KzjYgeNJJ3O0b9Tyw/4uDhka9xajaxMBmNIN20D7XGmH2S9PkJR8YJo0Rkq32ejol+Wce6dZcpPA
XcQxTFlf7wrPrzOhKPMOInbenMXYcnHPjIxkAp4E4Ga4/vwZ2s4RURM/LQHZaPyAr2iue0womGbI
FyGMdjasJ7SEMbsVDfO5+zY0mICk+6DSesiYdEI7fABETFbo7pdifQkKb+IfCmvp4ZhrlvkskFzF
jYDmsA6f3k8o7KnXz9HLO0dbyS0MHE1FVJ7vY8jVStOrru+aHeMkt+QEXzG+GjBWdkHdL1MMdwL3
91gFep3EuE9IQn/7ze0wZ3Yo3Esd1OGz7HaXe7m4pkduTv9Y8G0az1SxIl8K/4HS74kv67HIFv2/
Z+tG5MOvu1t3+0Lx1RQ61YbYYgd0OjrDegzFPq7F03krWYMQGwmBZVU6QjWziBCso2GSrYxzqeFX
TWWfsgJobH+XHAbv9mj9snk0KacyPhsfwWS52GhUIL2VJkCUK+vTGREyU6LUItezaSak7UN8yzpv
O7VvgZ6DpOJ6LxOlGtY+oAPkjLzo7WpwyY2LllFlTRo9yCfpOyQJqsNGpL3Bub+WvZ/M0u4GjyPy
jR+JRR2NyArvXMSSFZHuZPzUxMVmj2qPgT3UOzy3ypK/uQPumdvCKto9+VlyBjfL6GHJ3hs6QZ+h
m1tZXuyfyRl6B1nBctLCIcwKC6kpAVJ4fwMezVGZzOt698XweLPDKg7WS7iUcZ0D6lmreezizSwT
4tAjf0+EM+WULM/Ys3L0ObFRidATQ8MQBi0TC9h5RrCC4j0CiyXMhWXb/3DvttncQj370CPFBKWD
nCbC4k6jckvKZqDTLI1zJSH/8kODg6dCionULpmBXBe1/gR7B0Rt+e2SxUzK9j3SFhZ0Yrd7oQTp
qAqolqrmjVQrUqh6poTh8PBvL8JayDQ5K0jfLYzjFN8FCsS7FXwOMgMPBoEBSvKcvdn2OdLHU1Lj
fkW8DZX398i71m1mRpeOVkyijm7vFYK7iUIKVq+dzQQ4hvuxgVw4pd1mhgUwZtBVPG6h5jwtXHkl
RhpsRR0+MgFuagvzheVvDIIALp7innXlFusXfWMfxIVk84waEK5I+lkd51Y8521bviEwC7ez+ij7
YwVQ9zJ2gv+GcKZZURA2jSPMmoAfTaArrDCnIBlYDrNmCl9ZUz/zS0wAmKjG3BsMZIrbHNTTO/q8
+wWSV4c2nBPSVGatyVpLZbYyBltSPiEvSSlW7/IAqPAdDHZ8SCvbt93vndyZPtKmB3KSossRQx24
i4OI9tDpwm3cZOPHIhMX+jlNGk0ddwUe0E4gC/ury5uRDsPi6Uq8yruBEjrxEsVu/z5xzv+amFPc
0eLQwdHuy0HQTg8Pi2fLBRkG4Wmd7GypX8Y5bNy1PQqbp+S9H2ENNiMGjCX2LIit7or4fhm4ha8K
A51sUAnagqxCOoKP9xiMWXiHdMN2KX1QyyEGra2Rpo7XAypXkAXlN49vs2XsQTkyqKJBhU8rBzCy
X0pyw9bicKi8vZuxl4caIvTU4e4I50Qy5O0/rlUL8zZsl6b8rOi2bz5M9wSvfDLDfWJ6nFaiX8pS
Q6ntL2DwdDiTeoEs3g/bGeSI/vsGx2fIT7tKl8yQBmXI5sm9i7JuLps2D/I1XXya6GHXx6WyZQZY
noo1LRyKsRa/hCp7zO6XuBtZQBXIWM1/U9uS1pIUYx39uAH0FjYjJHML184/O9iXd9iatnBgOmaR
B2WmnJilmAvuyNSa6xso7lGwgjRjJuxCUTA2aU4CYiVYodlnPUxMos1rifEqSkF2QgYpxMJt9nEh
QVPoS4D4xds6/5ULH9LXsTHPNbzk7o63FYJfEY9hNVaaZyHhiuwPTj1Web2mDXTHQAwPex5mcc5w
qtPakmroOueReiboBdopFRGMFv+LKxOcVvOoRwSpp7AKlC5zJCTAvlAAwzNdqZVp6JusD9zbDD/Z
P/cpT5k+GfZnF5CKQK9Wr2nunBYan3WgJBOTmnVWlvu5MWKMq8+gAME2/fICmw9UnvUqJ6e1RRF7
DgfZImHQOLuXFezSbf8XrfIb6+7/ZIOHf5CYjpgjsqfoIC52qNXlcIkIJQnEAjMRCn2K1ubNhj3w
Ydq3prWFAO1UtDSBFQEeh/Pshn5AMdpPRs59gE3Inmk0L6XFcjzt/Q4lAsJgJgfVfZeKjHLLlYzj
lvspS2Hleb/ZCvQJpsSUGX7/DaxDeNnhcLJRDkdaGlkhzSRES/TV5YxUg024doc8aNVwpLZuoi5I
8N0lTOr9zUkMO6DRT/T3/XXgvmMc3olwlW041jYhh++QObURHLk5w5F2QbAuaYpYzGMy78gF2WRS
DWAuaXVdV5eqRxrOe8FH5+Qjunns8p4GYjD66U/nPYT5nHEqhIMuw6y2eFgFjbKYCtgDzClO/LCo
DkGOyVcTI8mAdYPSX3CwPcoi27g89Baj4GO5BcvWCU+DAbErV+j9txy2aEO3GCOYMV2mg22Xlnh/
xhKpIHRzHd2chO769Nf+ZQg6/nlS+OYPI3yDaK/dH7ChpEYuDrC+Auqq91r5y1K+JtulomIGpeJm
jUIGhF7jtlOMBsNMjBgtG0X3SYKzzjXZhJg/AWFqhg/BZwwDVDYEzmZpIe+p32Vr7L9l6jBUKhsL
alJwlutijk8TsGp1jl7bchhF3A9LPouO3tP1gu27OyRCoAH5My8GfcyAHpnWZtEyCqzhVByPqN/S
rfvbgqBOeSSTfE6SP2/0qgOPvDFC9rLJ/Hrk7wcr+eEwP26owDgOXuPA60HvcFV4YTh41MNFqzbI
mXGGakCZmXH+3cP5wOsq+OppgCXf4uZ/FjqI9ZHLel+Zir3I2fH1JrLi7Gqo3DSA1OrPYRmx9nRa
t+3jSVA34FrL4PQWXUtUO4VJDZpzZDUVvjSt5vTg3AgCdIuX7jXvaZKiM6E3DAd05aE1otNlv0MJ
5t6rYhBsQ0JmeQspDZEyCd7naTwlZbPYTeZ98yR4uY/uM3s7CfO/Kws0eg1OSQ/BLFmlove+Shw0
l7Q3f5ToSDA17Nt1imzWLrrS9hl5DYWtcVHH45r5qMZpxi77MEqWkypCnIdMhPgCjgG4bHRGGG4c
KXcz0Srdov6hCtqKjjbNM/7vj3fPVbYM6pR4hRvDifTayJJbGptyY0dczwwc+U9Ep7LtalBpHpqX
WRSVRw4ySkO4F6lklfYO3+xUk/NBo873PNzNmRntVRtHjQI2NDTG85lrTodoZUl1+RPob64dd7Uo
YIWlbGQIuMloXXrLee8o63rAS+LGBP9BQiRjm+gTxIxPIL6qOsIBFfXRo6BwesO1sn7mU39JGTS4
r2PMFUm2M/LkdDgbzNDHc5+ewIA2ct4bBiUiEe5WUVGvvd49IhAcCILns9djttIjLIZXCrHPQXTv
q5gOyUER1awsr8VHnhI8LXo2ZTeb4SFOA/f+ZY7O3g0DPX6MCfxYf1SfFCJvHIhftBup+q6EwK6e
VUKuoA7r//YGxVF1tgQ4Hy3n1nC9vHzG1xm02k5BeeWwd6fRLnGiCU/JxPD2s4OHS9nVRUo5Z/rv
xQtf6/ueE8nTpnhk8LJ8qARrnuKdXrvyhRQCLz4F7bJsp5I2oWlSqljOtflshXa74qljdv0sxSup
bGt29UAsXiot9zm9EYteaEsigfyTDP17lGPPNIXZWu9KKgQhq0y/aRvp/FbSaPLKPFRaUUdZnyl1
QiskWFHk4byyGwMmYchJTtijQ/C/jNXIHEXHfcrKJ/0ACeatk6bth8S9rZfH3M8qx9O2cGOmfr9h
eqxokAr/mM5PX/33wHje5t4fLblQ2ptWAIM+4+5ENwSEKq6Ez+fWHX929KUpP6NrkIvnCotiTGdv
OydeofQ+UmYzkZ0YeaDLBU3Inv3A3zbkFyqHA8nPK9xF5c1BVb1eomoDmVL3NXbVwb4mkCo86IkZ
W7qzDIhWtGvI42eTiV8tcZ9Q+DK1D3nxwpsegyyk90ZzSncaL2F2G5bgZSVLmGXGhJhAU94EIN7k
tuU6DPihBxNWkpG+N/QKqm3HVThPgu8LbicpbT3U3hRzjyWVdrx1VLi3ysRwTrPUW9mK3jaqdhbJ
LbVim60vMyDKYuUmo0dzYEp4uRoAPPmY6+yQT6SMjdRONrmQQe0SViv9fIm7sJZ9Cn8FR2JcwSwQ
iEF+yVFJmmoVz9A4TxN+VLXSmTCBeMpdBcYV8ecxPNZ6CKjVaVwUGS9HcG1Xs65P1VFrLLxOmZSu
Wfg05oCEXqNQ32cswaaPenbmFZExH4LdGe9qF6I0fKOJS634DEI/yUpox7JBU2L5x6xGyQmzgm8W
a8bkY4TD02ikKboctilA7/KRBxP4e0Aqc6GxDP7bXHamvK1pInkADm5EqIna8AArEY8LImXncJcD
UsfRM2pBCzu4bPqIyIplmq0M+wop90dGV4T+IhLoavN5qu/eFSqO22tge2obpcFYv6TH+I0fhk93
bhzKubHNbt/WsVsMDNzvRzrjQNs1ZHtzLi7yjUI5tjqI+WEMJVWBVt/sDTHAW1BZTr5uJYkJn7xp
etIYa9p5FqXLSnoeUvMkPW4ZVBQ8NULCxLoz3XKvzsfh6wLDZ3uoOzOT2BTTx3f9KDlo1+uD5u8h
NhVr1fH65/YdU0siJ5W+gmLRdb1i69kBdS6gAaCha5gOCvM2RyVIcbRJqq8nEV0UN3YXbNsFzwIx
aLHUt19ATTcsEPKeS72G5l8/L3jF7DbIYDu49qmUMhUyS7ibXSGSLnvJ731nlh1t9dYgtvcRlkEM
GK3KmgEWlvAle4q3BnK+tfeXgVRoUxkWwhj07slfSjKg37DeBFybODjy9wPVK8o/mAwHPUNyduO8
K0N8gpER6uc5LWIKK/TQJkmkpChycoIR3Wtsaj1RVkHP0mnSpxo4rg8oPgsPsFe2V2l4hYsJnr7a
wahui0bcnEbKjWfG3vT9cx650SwUJRTIb0Mc1GtM8kCs+WlwROZC0biyxJuOsAHVJzIGQb1ZQbFW
YdAzpyYXjBeW8ucF64C4AroQ20EachM78CQM1wiBlIqcBAZukN/6wFKVM1obDLxtfdd9xzKwMS7H
Vw37WaoQVTOQCvUYXt75rLHdWUV2KekAIJHvRSr5n2H+4mtS0xZV0z2jRUx10VFuzH8BMepfJVak
v23eWST8XHMJMsnPCUet19juLhHCNrv8YmrOWgyGhdLNoIVnpEN6K4zsb2D7shtbV0LWRSCavqdE
WFKGkcHrjejHI9LkpvA+xEQGYHv1UQb+lhjkG+0cGf96bkmeWYe7pEsyHhwExYpYcsVHZlBAsFIp
jY1igxkdvrANvrxJq+w1GfJ2Cao8yJDzEsIUzFZf7jpPdQ1U7Zq/nYBoeaDDGDROPFKNwy7ylr6v
ZgVRjtSEDkLIzvMNe+jO6clNgZzpq28NiUAisiZjt+fe0wRBt4/Mg/ux+d7vUDF/FekREVz5HctI
itjeNK2SkmVIjGdEce+89D332FoFXtRVIxfLpovTxQMFXD7ecNUcTTsd3B2mmLYUsI0nVogwa2al
kZ6ZDTuX2H/F9BIJayygCj5/gtJNkkk+N8ZSx0sHQMdr1x2uA6qsjviKJ5TE0ImlsBSmVoo6NSnD
K2C57vY8U9NGUtmeyMKvW/upW4mhbtqOAbKhsTpuFPsAaaojXOy2dPSxOpYKrgcfsjo3PDaMSqAC
i3621lmUUkbSH2+s2yVXZWEiw+WQO3MFdrK73/N9L9sgDgcW6269koIS6ovG2uoeRR4yvrLfFM2W
FdyYYaccuiTSh8qRjv7DKWzJ2siCKayPkP5fzxQhBc34LbuTJswq5CJtOG2NNWM+pQzXN9Wf9SVb
tDgIDfJgqz+GsLjKfuKZ+K2k12AQ276J8eQjiFS/E72jgft1ySwXU1vBf+/T9GzpFHofmcaaZ30j
f/BQibx5qkXi2T2Q7ekE4emdo9AcE86TnWee0M79emDnX+4uoOnd6kzK598Abq+LsRwo3Uxrg5hi
RwPgE+cepb692vvpCR96ATlA80DxIkgOfVO4ruJ8HcDt13jv0sFTLWo0DE8IS7+iC2yJTCY7Y8tX
Ly0Ndw5bcIqCwdSpy3sS50D6kWzzh4qksADxt9WjMoNROl73q1KPUseNbktW1O2eWNWZajwrYgpB
rWQcsqFq0ez1ahU/fbKWterjMKRDKfGM8cjKpF3ADXjBtBRGbCDQUwwoHTv4WwVexUYDjerSdKt+
6f3Tv6tphJy4O8fLX4qUZ8ySFSX+jh6030pTB3eXQw7DyeFiCMZ8ccfl1AZktohivT05SuH/dfk3
DIJsS87cT72sN0WMzBoamyOfGkJSgB+Ia7ESCkg2T+pJ9MbDlgkzlE5eBWJdkViGReumwkKDvulf
O8ji3X1sYXRARMxVL9WfxXF2WWbIvgr0KHuqQDb4QrOkLdh5OIYbzKoXUm2As0cq5/jb2c8+1ktR
7Q64w6yWzxZPwbg012Wgkt19rUCZd4VugbUbMib/exO5Erwmf1SR9oVm87+RPAyd/mp0PbIWZak7
mj9KULvaN/fxiKt2AiYypa2RH8LVnguWG03fyObXdQuvqx/xmZUYlKYLmUPxUw9sTD61AMzcjfSE
slkwR83b64wEYxIVkaCK1hN+4RDqggNf+XeQZt0q03cTZI0LrzZqUXoCYxd+X2S0eiyeYBPHpTRd
zPiYCpo5Q2qyWR5HKLqiIwo0vVOGS1C4pFuclbxxLANUICPXg6WRVelo4J85ZrVLjqmACs5FABrq
zRw1jzKYJ2Lqgbkk0ykk0N5Qt0qqP8BGFmhEuW1vq0ve2NLsQOSqaYIyJbeYP3aPT/tbvZSdQrUT
+hPwIzHi+DGL6piatUkXTjbLTS6iZz/xzFoqi3XI6SEVlHsEZS3IuTLAkfil9zXFUabaLEB+Pw9f
CbiPmojMQO4Knl821dOFZI7JoEvKHGZKGreMhHzEJra/gxlpDTJWfTEwKo95vsGdxpvgbUb9blax
K2GcDQAfw1k0RY4FK1O0qAeeg2n3cYIHk/ReSNqCGLn1uA35GU3hn+WfOc7+B3bn9QD+9hpa8sic
ODep24Kkfj/SS3JX2IkRiOsdXczfUHv80rC+fL/9F6q3nkWDuqkPhTE88dSSHN49yyLgfhxBbthi
xIbZZWxzETv22YeH9uyXS/EV4gKn1pVNIOnexWvNfVL12C6lUpb8GBtiWFsm8SyiKfF4VtdXnDX4
8OldP7+FekjEAeU0AqCJp+Mjc3PNW1B2fNetmrYTpXr3T+Grwy19Co3r1IR2vjl+9dyxpUZFRIUn
iz4gkad7TI8c2n4CqNPyRkGR+UbmOJ+zEmjJ43eqRtZBCJAQqoWYJ9MZ0N/ePkHIopdj0TXfZc3U
zyDnEebdYx0dRrYV1JJIB1t5Wnna6B8VAiRDgN2Ljd7wcErhcMGtD+rU4PzNK5pntBn/eOp1xPcj
DJqwgxW4g1cTjXZcSxDJU4DwkNTwabKMww0yAea8WaUTLSalMqmevh/kwU68Bagc1BvVDpgIoE6H
MJHRqmc8lkrtnlsiJVYeCKg/L92K26+U0d+wY5eKRjMNL/1dNWdJ8MEZjFV1WqD+J7HiKkNVQdP4
rTVX3CuN/9c7Wjnp8y7Mr9k3A+XRk0DquBvskS/C8Qwzori2vAdz26RouDoe/VCXMSdntn+iPet1
spoB3xOL2H/Tl7q+H2TXIw/Ky+bNEk3gOQ3u51sxLDuYctOcx8WBVYs5CDPITMXUpcxDHzgFnLrh
7W2mrNymi4Twzh+8BF6J0l+nKZKQRaF6Epqk9ctAjbVULvMI2ddUxT25H0kTzWVFlL9OC7pOpQJn
3HVejWCZ4/UBs3GG/Euj8mv7EqefNh8lrBYk6wfZWMh+QRDaz59wAn7UXqe5U+PaqnOas/UhVgVv
GcVWLuSpSd2sili0GhBzaRdNb4w0xSFsjud+1038E485WZAP0bct2RxjVMH4Mqyw6d0MTzdm/i9i
NaJnvaP+yGWZqsHYw5x9luD3UDY/6h34t4UJzwLps948/HVe29i1xrwEtIQlwiSWLiFw0iBAdikF
6mkjjiXbBvVd3QNxa480m1nF4wrlJytrox+ML3LJ7KFRRE3iWh/y+LREfkhFimjUrkQkslXo1PFW
MElNwxRbLeEiBGC+mvUOn1AmoGHlBCMIPmxERbeKiuc0Xmce92udh9mB2kKJkZymBQSKoAhS9O1j
OE0e3d1IpEYwD2UDwda+iBg61NkeDubuf4il+idHy236LQQ7J1219MaK34sXgMkZgtMq/cBTaD62
gDctJUIl8Wa763/Dx744lpLEv5YAcR9yN0p7m9djPBgLowE7tIiwXdmP6eMemub7BMtBFg0OEUY8
l9uDLMCSAi8uhC1WkZf7mjeItUNbdT5BTsdbQz4Cx5ROK0ZCupRY+0Bjtk36DVcRqeQWwl7n5pHl
6O8ACxfOiTe4NLX0x58PK5/2oTkeXgD8rCKamjXkJOVBto8REXrduWndtLEIu7sbBY+UU/3sIu4B
J5amHjtLc+Z7pHstpbodJXf3xgJt/rmHLNPPfGHidHT0m8PxHhioz81sWu+cIi1j2pg3PVwdBfQ3
mB+vfwtXqcqn8rQdMNzoAPkztqJq7nDT1LTH1R8GNALrSFj66QrumMU07GgOm1TwajkJnx8kXg9K
7r1nLQKWw674cj1ZnlQsFD2uJ9Osk1xRLWaClWwEKZzyKirRP5y1/auxLgRxPDeGGEguHA2Z1gxk
X5OKNAondwUGjqYIcpk1dTWVcVpPhMBrZJbfpoEe3zEwFkhzaDkfe9WcX0CHodbduXHB4r7yLeXd
XPjGhhgpIuVthLnWpJCbNjMee6mq2EZKE8SmGKfLxjDc/b69xmIMctmbFEN6jWR33NmSeBRvpFDp
+uYJCV7WIN5L5tgQQCyTOwutIwqXXbi3aQPpz5Ol1CrecCAJgum38+RvnbjRHjc+TuHvnG4MIQ+j
lBQOS1f98tBC4Sn+7qVI0ptClpyavkriINPbhc0k9RqTnJkuX5rhExz/WFwUryIpWBGSrGicW9hT
2dxRpH3SyQvn1m70sTdvokQt08bHlaO25mxoJQZD6sEDLMYOGeUOsgWkKlUmefIby7/HOK0fp9NP
i9t8b2Xrk8EvpB8oqQxaC5T9VJgTjHeCaQ1PtPviqANuF/Ht21RW+QdQvUATCaCspHzzc8JmbOZw
0Zl7bbSeRr/o2Pos3U+Jkuw7E9QB8M30BV1uwAxEKXQXRxv2A+SUDDemaBL4KtVWu2pwC7/vj/Ki
wbzDC0NldOVn7RsorAGa8d4N/voUNRxnh/lYezNf+i44rZcAHp0TRxJNdYyOWoyUmgIJ9pAXltjA
famgH49qiEyyz3UUB9Ts9vEBxxcQOCWE56xwisdl4UBYSgxGJsk7/k3j7IVSbywm/BBHm/+OqwtL
Ivw5/m6jWY6PVAdL3cxkQdVIvBNKVTm/QicY8vsPv737gFB2vwm0nVoBDwLS205xDBDZ6DmvagAY
APgyLLU54cW0y/WlQdgyekbDidmg4WxVo3A63P9DOZnBR5X/xDbAKAqmry4vhpyjMUJA0K3bfS3T
IZ/Wx7TSsjJxk93qKhY+cvVBOvH2PcC3pxsb9QibalSO0w3CX7+HRXz9wO1IStmECp1iI4cVXyta
8UZozbS9LBJwJjp4eXabqqWVZ1E7EJc2d/+fAAqi1lW2GbB4I8+ATiRKDs7Zi9/LDJgxqW5W9duo
DftBdX/fgNa2PLYKiHpL/pmTCk2jPY4+AvuPNxjUuDyjOnsr2EEbVYmlPAkcp68cJhrOp8ZOT7kx
uG/ScjVsthDByKv94t0DSpYXIGeiBdb7YaJ0b5rbJXeGjFtTqDYKH0ycMido9LlVOk8Z4C2UGpq/
CLmGN/6ln0V3Wki+CkAJOx1L+Gj6jKzhjfqKRadag8HO/0EDequ3Zj9Wvk52880yqiiECaZZeDcb
SY3j4k+k65P8Jz6wSrSmauQd8cML2ni+b9F0QR5rFDcnRZbBrwfZCaMO1/BQQ/Z4MapwatuTfYwW
bOK548toiFF2tKFl4ChHSivoWl3XcZIoKcz57epG9aBJHewr4vLTGURJe+MUeu51W2+A8gykFaxk
/Tr20JY68SHJkdUGJlZ2+ebTHc/pgZZhsqe3IPrFvtpm0Dys9zOtDKFfd0T91H8lc6DBE9RK4eej
C9FCys1K17PfOZYznlLY3y4FAI0pErT+ezk8lk0T0xNoEpuMuC1qNi1bUXBpCvX+93xR9ycwk6j4
ijJL+Zdst5oeGG+TTjogoIU0gJKTOMd4KfJ/HD718O/04dTVhZIVqoJv0qqYYeqX50kP5IrVdFmA
SzREP2DNGoyrxvEpFLC3M/IYvc0OiquMOxM6ByGkrxJ48tp+qMiIZPA0Rt7XM7K2Vope+fyQBcek
S/EOBMS7xW4KKJmylUvgVq1cxS557P4M7sSSxv0D/39nTPsHZXk9+ZTyq3HQfyaL84a3/onfec5L
ILvND+huPtxtQKF6UZ0+N7nhKKhUeYoRra3tSigXhkXoWbPZWkyyP6cAhDMwN+TjkeK1KkbKSbVs
z9Pva8/EUbPoTPfOotQkfu4G9L9SSLGNaYZcm1ZhjdzzmoZCH7XQwwcJAejDL+H4vljBELVC2/4S
DFBumAgYUd6GCElPc3V0FNSoyCUu0TDlW69yOT9a/jXGOm5uCQlga2jlQZjk2cms5Ykz17fM4tUi
PC1ya9FOHZjDYiGoOcsX3O9dpyf8uA4xcVzG5Yt2FE9pBfDqwlgPQqFQYsmAbvgNKHFx6HBouuhg
CEa5Xl71QQFVqfm8afvKJjPKcdzvKwT9f0IJK1KSfq6cUEN+1Z3ZRofdJ27mQz4DG6nmDdjyUNUk
FamR8oJ1uTF33ghKqJLl527SVYNbC9mh1Bnvjf5xRofxBqjRjNjJrt+chufSbmKuVsak+kVt9x3H
DgiwPZ+bm1q3bsgyt9ezc64EeBMJtGLI528W603/DYJGandiGhk2YjK7SH8JPkyd1gsYPN8ZUcvY
15W7xiC5GkfAUzmsieAA/kIA34eeZ0KFoG12Li4N+Tcig1bD7Qxjh36IdXzkGafVhMAzT97np5YB
Wi3J2DyYHpXAT83T6L7ruT/sUgU+En2fItv6b/wYTZ++gJZgkGw8jYKdlppeZdv21fMhsT0P/aln
7NF70xwe1HePbYeQhNAV/KgkspM7mmY4oyaXShrN61AHNWm2EetUSvzvkBzFRVIB8gs5LqToeDZ8
X8MfsjVz27znFxXQ5Q/HYS7LK1nZqdswMpV9VPs5XAZ9/+yIdGDRoWz5rCc88IXBLvhAlf2AbARg
QxgJ61jlEYph57vTGiQD+2U5kZWA6KQX76XZxdzkgpljZC2t0ZTOnAVeroSv5OtxJHR3//arrVpY
4s2D08hRLg9vqmf0R8wJ+I7XRi3g5BFfoff0K6YML+8hYK1wC4Q5vvFm5GaWxnZJqG9sLBO+HfnS
gT5Pf7ghgq+c1AHXt4gw2McnyaX0fg9Co6188V0LSs+1Ljxa/xy1i7zrVPWilogHsG/xD3OX7/np
lQwZ9OUBXuYK7q0MHvsFFIBQvfW/l31mldbDhkE+aH1atDsp67my4fsN/PJ5tNPWpBC4Ustscmlh
lgpF8MLNUy9ehbhBxY4GEOI1WOYpNiK6rjHBtrOZtFkGjQp6nMumdIiQ9pj6jpmFA2Xuz5LJluud
8BcCPzDH9uPG6yOE/CDDgjT6elPEttIeIuPVQqCjt3cAaWb0sR3dFisHlQeQtqivn/vCbxLODpR1
g+WSIyDLR/I9nsyQ7xxvLVtLFPOVV3vgMlfoHS4gbK1urVa6zTJy/ldhukWFcG0tyjP6yoCgVtVs
SMLmFsA83sUDkaHKMPOypNBs8JQnXXB7c06x8+Igamxav5MA4qqkmHe7jTiJ7Sf/rzi5lwERdowJ
0kqcjOMfCocLBkRGbPW0dKqvbMX240po1uYBWoAYDZkz7Hc8cq3yXJfvApC3EDQD94vMw7pZ2Lv9
eC6UJz9JGGVURDK+RP2BSC1SidisUp9nHZr2/SsLDXzp8J5HQkd6fOarl93OzROFjpg01v2zcJdA
gK4EI1wjUUvphUQ0DncL425S0pqOsnQEZxX8uKNC/VHT1xHcHrWhJsp88SGqOXqPmkB7QUdVdPJC
so9e3wigpsPsE6BVLhkDw6+3/O3h4j55iTY/zHTkSHoYtZ881LqObTx9qbNjGZSPg7+O1ImMKWzJ
o9oXpd3+lBuoHuOX/ZAvDwTOZBwjw0dM04/eeLcxRTq7xL/gH4aKUImBR+QrHHVhXDr2+rSCKcUL
88srfC0JQVVO/06fiyR5FoBFC8yk3pP/ZVjS+dNu805uJPE/9lCClYcExpOBoWitt5K0RPS+VwA2
hVzH5vKJPGBd+ZHhZK0dj5dfnbMCGnEhUeIUJVuLmqE50ipZZY4V+uC3qkdIxXtJKy2FeZwp9/uK
faehntuUBuDUVgsHC3SxXy0VZota6xr6KRpisqEoPKrdoLdq+mP3qOvW9k93Hn3+vXBF/Lhf6hHc
PyiXrwO8sSy5WfG3bSKpYVJ/in+dC8+0uRL/2O2OGQ0F2ZxHUACBpdoLc0GNkpqLo68BG5I1002x
lyDJtArozyblvhw02bCfTMlqA4GyktTXWmk0djuYYGp7KB2PdDN+eQEdS/eFASrTaD2gN2xUmwFy
W2zrOLRAkUXcSiUvu6OBTrPdO+Lbebdn9idNjUhDxSbU4FeBDeBF4T1FdNJMO5MwfdmjXYFxmQaS
t68s96kG/v5Bl8dmlYQFJlgBjizLBWuovpWTRcvvXBC3Ccg6nQik7oX1HwRUF6uKNiASAKrzYLmX
9Piqrpwa9npBe5VDAZ3xbp5MzyL5pLeeeIpiysJ2t5aYPF0+iV9tpvvk96WwVYERrBOAO0KHxPew
J4COCu3KgNw6cD6AcrOh9k8kscEoeCe5Mfho/zMIXPiCqcYaQBnl2uOsTgfzZgb1EO0+aFWFaOvp
whEAOCGI5MKtQ2vw/stGykyge/QBXxAiUYyGt2qnUHWAS6twseRvLhTctKdBusQPMwLDalAKNVSi
CfhKRZD/acFKgeo83ZmaEAWTp9vZbaIzTwuip1vDYmLv+9ycRqSs5DW3xPxLGDjGCpg76mJOhgsm
hB9AIVsFDU57510eZxuaCAz8njWbwsWf6RM61NpZdgQU5+/Dq1H13lebcLBVNQnZ4Bc9yRQnmbGV
sTuT+E2oHrTrtjy8LfwyvKcT600z+8Fa2hOByLnmD4NwV5DxI7/0zlbMnxxkm8snGE0KrPoWqYhB
0A1zajXRm6rQ7WB9kz4SFWjthLvUaweZLOaZaLuQvZaNQhzFINWoZ0FFnP5ulQPZSlmb7cubtgsi
JGc4Ezj9FQjxDEHn1RC/WHzyi28vYRgCfr88XnM5LFZU6oD8LsYpqSfHFa3QIWfT2H7ToWP4eFff
K+zRq+fY1bywC1oMZeSAJ8GI/edu8K/nedUUXbHEQBAo3i1f0vxgXNdG0vkbVPTKAzcUHwjdFhfa
JhREBl4tPxdAexvIQbeahu0rSUmswaie3fPhpGy98X/FaD2gccSnVpM/qH6CQmvv6xFGVsLWTBr6
6dospXY3q1KF0RzhdqFaIrjXmHGoDRltMqPXXBGg5qJKNsM2ViiyDrIRRiIMb68NakI4SCNv182P
wouBVdVaUazKuERzpJnhNU41OB00lBnRMmaqpC57+zYx3QL/EPWxD874M5zbjJMf/l0OI7p3xn5Q
xwHLF3MA3huxSG500Y9+LxRO2gKpn2qvzqzdKESbtLwSaZ2xxZJW1YK+LKsakt2f94KiijCBgsLO
Wd8g0hBtsnz5BzGsZH48jcx7WsyA8SUfJ13dOON/XbfAxTMMsJCsWXfAMnl8obnhH8Di6RCyRVJC
5p02tu281Po8cqGbTfmk8EuzbJbrFg5mH9Op6q2Ln5odfElit0ZePbJJNApwrCeP91eVUfiwnUuv
RKjMeWZ/DM5hNBd17iFv5YXNsltufNkISbNka/wRqXC3AjkwAC+aLiwv2K/jMGvv65k5VTJe6yKL
FH1Jf5wyV/BD1lsOh7XuU95K5H6deB4sQsOv6BKTQ8m9RAI7BZJEGaNA+czLxtuy921IfNAIlYYL
bMuMbVCZDNQb05xH7Wz85BUEiky9npjw3lOD4yTNk/wiciJFo8pOPocvbkSwO/IN0j5YJX4GoHgh
nxJ79kF+V9hO1hLw9Q5eSAIe6U0luRSLsLwo11IVoIyjTmKroRM4NNPo+V/AkoSNc8/paFnJODPu
BffI2mM176LzM0rl3VlutDONMOo/0rkvPyVB45aOXyVA76M1S+oZhs2fyCGcfA/+g9afoJKXRNvI
0OrKFtjckLin3YYoljaOEwlHsoiiONys0FJgOhPw21/NezM8wIsOVjIDgGCjXE8XQHWwd7IqVJD5
1BIdfGhghBKExM49CB6mQVUJ/2kFqPvIFA8xz8lTiWMy8lYNZKMMI2cwRQG0WT8nQFu/EKCDTOgf
IHsJ+eq2Ca85cq5rdv1piuxAbmeLFf7i2AK5Zfnk4bovQbybZ/7HFjlBolEUUAQ5K+yxbwUI8pxP
Rhtqt3gxyegogIpXlfBQUbuyGN3h0bi5vfVDHdnrIHfkogK0OE4gKRStMvd2VprMiRRDzjs560Sx
QE0dFEsGVzniIhPfBpHKz150N/lpljOBMUYsMv5IteJsaHxbS5j7Go5Ttfc0DeG3bXlg6AH6Pcjv
cc1FNDJdNQDH0kHBynjcFh3Ok0PkTuLpG/tCRl8vQAkSstHiX3dopp3dc658SvAZ5Xf+nCmuqJQB
3JQ7DoLNvTsf16PdyjCwmLpKnm0oAmspxE4IH0mh7zStBLj+6eOqdv1Ox2dMq1z/+LjJbpoJJPn3
31VTpaCu3MrjVM9dLH62J/smY1L+J3QvWIZ+Ac+7MhgT13Sw06FIeI38WkWWRQqApB0ku9jnMfUQ
gH6m8f44XYnceAl4kPOOzbBjThrKvC9uCGghnGulLBEZWAFfjcfU/7W16mtKNXA6Ldn8zNNrUC8V
Pua3Bmpv70wT5a8c3j714Z5OXeFA/s9WIC33SJEzvDmulTY5AOwx5tT1JW6Dxtei1Xdt5QmZ3v4S
HNT2ow1TuM2S2QbeOY/Wm+JTw63ScDiLlWEmq7wWZ+LyG6IHb9Glijg45VJ5ppSnG8i0dsseu7Dk
r5sp3If955OJ09p+oBKo6sIesKnMNYsfFeEpVinQabZmnmOMUTXk+/cZogxTkONj2bE++IP0hh5d
Xg7h0ns+cIKEe+9SHRjGcTX2OC5VHjY97qm85Ckf1air0ImCW5pmU2s3vDfgz+v0OLuqZH/yOaqW
RnA07ysYDpl8S1/zhnzK9bIMkTiLJjzi32ypsPu9r//88dEsRByeD8grSOTW/9Vcl3gu+S30hYG+
w1UCa2VDkU65/druHEH3tLrwxnDzljMpGp+mKPywy8oQqcRMlEmxV1v68eet3yqxvpPSsH0CBjZN
XCyD9EbglsIfEnxqCiA1OEw6O5Ykx6KjxdSyk3HwvDremr5Rchyopzg+lygY5oY6TPDdSHS6UQRc
H63HJHPFy57EdlT/T6AaUknKFd/q1HxgJiW1+45BomA54qUk2V2l4cBS2uH8yES8j2m8Y4RHtzi0
qW0089ZU9Y1ZLZ/HJjW+K80kptBvEdjH9c7y4CtSNUNDdlDOxeBcBGLHvBE4by3Iu+82u0CRKvpp
KHpxWpBCY4waaMvqrwoFGvPC6oMd1GjwCRrl6MB6e+gSUpMAqDxQi2rzgHeViYWkgCaAOqU+YZX0
UG6ECdyD6BrPJGSbkjszoxaxpj86efVjjztOjUpxaCIrqhcLJsAAa0jeaWcwMiy/IFnyKgWDoB9K
cJKzLEmNhspW3hYHk40BGkA/x2HZsLXhLTb1fjtcLvN3++KQiznfcAzhtSkEjEjKM88AL/hVN58+
AVCP2uBp7+4DOfyAMpNLtIIR7vOMTZS1xJ8QuHMDrewQs78UB3vOSCV3oce4JJOXRnNml52DJdDb
3Jdnwkuo5/kogcx9HclBhKRSK9zGeCtDEI9tpWsR1pombAaRp98jmHuSjWC8KkdmOwJFDfCTppNK
m0Wd6qJXdhYhcJJnCQfk9OXnMu2qh3hVbpUrPqtLrcAXCY1oGFVk7OI1Kp08BTZwuoYRu6vU3UzQ
mCaU8IM41cmgFUQL8A+MrjbyPbYzb/evQebvASAW98iWrZMbGlXmT/1ttrQ57v9Nl1fv6+0MkqB8
GLQreMBbrNYkG6RI/F+aCaWrdwzktWAKcFjymB+m1BZnGw1O+avP6vXUxbIbJIJ+z/ij+8Rbi4Zl
DtIl5HcGmVT12DCJ7wGF6hODu5hfXe5n3HJO1TKcF/zM20jLZaXBxM2ANGHiiDNV6IAJK/YWiThR
Farx4umi0vWAM6Ew7vOZ2s+jfDKzpXwkBkuAuHEB/Aj3XkajibzjcTXVPEkxmRCaJkx4p0iUSdeH
lPzFcCiBkgVACdqhFUAUXWcf6JyZedwki7rJ+rrW/YmI+yZJ3v1ZMeskeoLt1LzI8J5gGCsermLi
cZjmzS/PZRO5XxHBR3RanH6Amjo3Pw/NxDQgLH+SGdHTd62euHRuOgnsmVyKox9+HbiLwEDWqZbg
b2a2OyOhISiikSxn14ywREsE/OZzLJJY/5LYupRl1v+3stg3KvqLVodDMEl47LsmOtMrB25vZNyJ
/ylKqSSozcqpyyyeUR1xLa01FL7O8/BLt09yllfW2ePn3Jvohx7bBxd8m74cjHw+Oa/UJcglogEt
YyDNQPnbdzwuMqkIqrWRxqw062nMyzttoQmH8qExigsKNhjv/bFG/i1IxJlsUnQ16eW3f0quzeuD
7jyq1WCLSh5mSIm9vr+tp/h9fI6fSWmaHC2S5R6Iwt7xR1GfSp2t5c+H0Yeuo//dnVPVK5n+pXUe
PygFmAigx+uvINL4jlJewfcdPUJEa+6gSLzX0nvJDy/vkMZjbSUhEv+7fYs+Q9+u3dENsUSi1/LH
Rdbn5ILWoblfTZt5NawisKtQoqvgk6X/4Lu4V6qLzVM3dhR/syeyNiaKAivsv+TslsolWzqDoIYm
O+JRiRdhbLmmepRVQYPBZ95+fGyfFaCdrTczTaFqO843khmDyg+e36/TK1ocv1jSkPBzfQ9W7fWE
W9nz//9B/kalGggSO35Sw3Q5kmgbFB+sbxZuutS697LxQsNYtM0TEaPVvkTV/QN4QBTYfBFufKwZ
c5nOvSiovKuQSTS6Ct1TQNpttMq0lWn8fsHGQ6T1Q2F/7MesQWmR3gm+iSG7VDzdw/PMx2gR1BJL
3XRcNCSWlFmYot+LKRC2uM0ihs9tiAPoWwXp6ixy6RyLoaMlszp3L7WWv9p9K4cUWwhURYKfWlpw
xrQ4RCz1U3Za3IgSJHieblLxxCeQ/xadalznkkO3jeYIAKEq5uFHsme+n62kGZ/6SUufBXxQiF99
7eBmbMT6PDc65Ix7QRcEPzJ+oLEL5+nrIluKcq6zRAyUX2DE2RXndVnoFQ7oOcyLW68Ms7Fc2ytN
dUxsUGFwvVJzshqgfB23eYEvnnoFaEIi8DRhgl09nc4r+PcNv9EUlMqCRUC33uYBvcKsOhjn1oF3
R9HUaJ25644bQB43GThKcfyZoI/vydQcs5mQD4Wm13wO7hVHX41vOcPl2ukJ2qRSaH5tOkPP1a75
gD+YAojJOZtma6LDyc17w1eWIlxyFhI+TUD4eVzjcMO7Q/zVX7jjnNa165RC+TvQNSL0cgctzpTg
K8sl69fyoAEwXVq41M/ioEebMrJaMQ2WrUPyjGeIPiqaDs06lShokNjyOVWZxt68ynIqPsqLmgMA
XmPfy/ng6OOxAkpd/yFw0V3H60go54qqrnogfuapjxQD3ojgBboTWzh32tCqER9Dd/8dckEoGA71
Ts1CH3QlLdBI7Z0xWa/4Hg9PEAo3ybAalU8d7A2IjyjgOzwOlcoOJF4thipT8oe7cLQqDrIPqIwQ
iWjP/QnjlgPqp9yIRQtfQ9oCvdiAeLJ8wCX0OBTURkyXSr7d9VP8QvCsPfn+7TLsLgE2Us99fPHQ
Z2/sEK0Qf9TOaYXvqUdRR+ML9+9pbMO8eZUrr/wG3tIvTQIEmu/aJYtvEoCrJlh9oxVFK4oE9AkX
E0yQImI91kaNCtR0WICOnLNEC2tz68x2F+8SqcqL0HeUrv0ZfoqGJvZSZZBe0rL28bwzNTV9E2mI
qhNnFsoaVPqXdQhVHDQVJGrpGwRa/HEW2wSCrvJhsoqQ3l3HwydxRoH+7Qm5fazjLPbwYwsMo8S+
wFDUVCI8llUy3Q8bcshkY7saqXnFntfmRHrtVENrIe5KlbhWXb6imyVHZCtAz9XEibt0Fdk2dWT4
/BgP2Qc/IplYsiOQ+OEtdfDuNTrweoSUOq26MhkpLsjWGpL3kW4aDHtvPqtwEWE1CC+q5ZX4YysI
Gl38xYmf21kPApPCMk/DN/dMTXM23/s+6IYaWNcgInagg9IyocFgcbUmZpK6y9VKRcccYDEGMlmj
9wYVSFrpllsP6FLPBGNZNH7YGy+s9XhXK4x8r0pHgKv9Q2OwBHlXODdWUIwfWwIQioBv2dd7XMJH
/Qx1IPyqa2mZPBecA30raVAQ059SpDkG7/dp1Gpc8tIHI8pc52u31pgMFzawIXmUNYSFghDq12Ja
+jpgYfq8UhsONx1jTVytja1T8TEZJLkaHpxuvroKqS8UM7pf2J2dyzK701t2PTVeg5imsn6GLfWd
R5I5/j6mlhMxUawNRyrryHE4X4FIXdyMqzUP7LbyRgTfHTMJMt86dTyeWvnFcfYlGIcjAS04nhqz
aB2gcVR7SaUrA8EOylKMpxUHxUNbL199CrbK3pEqLAKwpO3NKgeHqHUxTiqI/7t+z+ZhOXcLVr4n
NugIshFoR/NTnlwsMWixLAScQ95GpKWwNIrtlTkWlfnubAN6JyK/EMqQPvAU/HI4dtw6YWpn9QD4
4Fi0I9TMmOfZefxUBFWENeeYW3a4K1ihcEpxy/IeQxbv+6aMzSxvRvXNAtl1jlJ/Dpuh6DRNPjeZ
YtwyjVjixBWakdap+YuOzfopz9XXVRVomGBV5ECYUJfg16IKfXVRMvGDAhW3ydiCUNvY8cog+pGZ
kHI+rE5WgfcvNFD3qsuqukpGESJBcYOw5oYaXM/gR/zs0AYncq2etEGwMG7jA+CU9rPcosxTYT79
HUYCarZeYIZkUdflOJ0kcSFq+33FF6lvE/cQU1TDjMRyKDnhZVagc85IL699p1RmTz2Aa2ElaNEu
gelzCmHTliPN61T1Nwu0kxZ1tCzoNFsBnweJkGYdKLqeBnZO48tEUYVeDfI1R38DWUalqOp7gx58
5x29LZaW1+AgxRbQQV1WoFJc0jw6+eLe4XQIyGjjItOoSc6kikjVu0Dgrm72kTH+Mj4ydQyZGJY2
IY4ptxNHsg5VTRRhktzIV2CoG7gCfFwI+EE3oIJed7RknkIvx14jRpykk/j1T32CnleK8mft40ln
m6u6dMZQ/ROIcTKGpSqK+qoLKhUz/Ae3VYywTbIg7AvxVNMhBA7uQYtcc5bJy7I5D8HOiemQ3Rg5
kyNyZKFy2/xRMiXWNKy3rxJs9rFKStbGTaiPRqQ8td56lIaFjrR6rUtcXh5hLzJvgpZlvzdKxEU5
12S5o5Ge8fSDfBlmzCzgCAY/unR4UWPdK+e/CVlnSRR6cUDfmgTKanQF6kcs7ObNMNUVP8vxOE+y
cnZ8vgjOblCzy4gkQ2DCdJUfNiEhY87oNwqHcv24dtAo+K082CWZ2xTLj/JihwXSJge4l1pBbqP2
tas72FPzyXLm8l+sB8Mrr+cAgq0lsyA/0DXJZo2/PfyEE+/mEinXexnQ/7QnA0sbPJcuu6E5Q+H1
5TbFuJ9Zn482fKV26fw/I7QMbtjdrmM4UVvYKkzRJgTybi+M2xXDBur51l7njPzxrNxlsGaYXEuS
3f4Og+uBno/8RjgruXOgSl3tvjtmv/x3+sKtjZwTYkGB/eLacdvZyWryvs9KACxH3MQ1gZFZ1YIY
3tUGgxPp5J4yqBzAEoKd5yvAJQmQZkbxQoTyGSqe4pEHh7XqOJUzBdtfzqyl8usE4eIs5qYuEVzV
1VV3xXIX0+qkNVynvTUGSYxoSlvqVR9196C3S+Elc57F/OETqbfgZThVZWYfio36VEB6eoPdkSw/
QEkEJNh5pn4sSY86C4yACIjArhjDaXFm5bWZ2rsId094Qa2CPuDSePuAVJPyHXDp9D2Qj6vnna4q
XKnjImXAfClDWx6rvRczRvKxbuJry1hBK5KljHXjcw9pN3L4sS47cB/VMFGoA2LMSpIETorCZYps
DmKEfSv2u7yvqgOnLKt4TlczISW8iKQqfmbE6N61PDYSzPbKE6uVuTFxHevx/p6x05UwnS+Z857I
oaHa38ns0BufOF0JxZcppufhrmHnQ3Ucu4PAx8H9mSu9szbiClkd+7T/QQazFjDu1UcTdF3M3eWN
bz8WQ4laIEmf4tY5TR4yHt5sJiOXuk7vR8DyMY36rJxozHunzaefOKfQQcyaBIzbj3Rif8sCTcic
XV9LjM2uv1iJAA8ZwbG7wkmZyf2BOYgx21F2UIpLEn3jcTI3FmJXIuvg1LfEPUAZGDNt8koV6pX1
sTI1GBQzWGuAAEwfylwgYb62i3+EOs+XUXdrlJe41gTaR75usu4fzcN5yL+ccaoRa9FbU0LLolWu
4GBYYDPpAOtFrKRYkCwR3oY0grOJa8Yrr/JwoIPK3hZnTN6R9CghGuuqlSIPRvgzSMhed1kMu37Q
9GVnik4MUbu+W6lJsQgjzxQFiPmqSMX2aN8pMP0BjRyBwdydSNmHzh+3MaqdQa42aL5o3xNK4tFy
eETYOkgR3UuNZ8rTXTV6k9k/qxInQV+KGeTiuf6Mgab2Bqc7t+SSY+3xxzHrnxZ5dEz+sIAsU9Pq
sjQq/Ownb1858EqbDGWtPELnMucDGQl2rSXYxAFR8XYx4UUZ0IP6HsCF2JN1YjRwKwYNAoQmHiW5
v4U8FmEnEBx9Vb5BrPNgySUlBKTIL639LksskwaKEZdjRrCFFKVS7wyxPpmTiIamY+RdfAyQKUm2
WOIet1V+KLzcq8p+D4Bls8g06cVe/e1ohCBFVPXR4zeUfkyGx35mheZ7CuuyxCsRjMQHIHnQULiu
GBP2ec2BKlCujMrTukCHsg2FiLbkUg8YdaPlp2pgsiV2YmG67zBsdSXnE9mRys0kM6bw9dB58JyF
w0bgu/nztE36ybFtSKvD2SpYleMwrrb9zaedpk/+VdOQgleNj06862X8MAhbG0KnKS5+puaSphdM
XZ+DsUVZzU4msAjzUJlO4hrVldUTCwdDGo+G4Di0EqrX3152P6C+uBKfoEt2qKy65wGrmPCAS7XM
WBxk9Dv7rs/uPWTrkMWTt8wOzX87l7RXUnaTyfxB+7qlH8fJ/kJIulONj+w2KEe0w9q74BroHtxT
nM6gct2nldwT/YOGPimUj/eJsOt4xbEu0ftzuUaGA6908DHFnRxJAane2+6QEWE7O7PfcqXwTXwB
1quRZ1vfw7AE5hWYerDIaQOG35FnTeP/xTUe1oUPhD3nTN8y9d75MKU4ixXEJBLPeecndF6WQNbK
nAUY3JF6ILRJOfskWytJG6ig4c4a+acRK0dh6fj/nvCFxjMErogkEN9kci9s6+Zo4G/I8zBESwTU
bTKtC2qSEfm0FlY/BSCXldbyHwyAiH7525OkbefDaNK3fOh6MnYqlGLAHnU8jtefugHBx11Gz9pl
YP6QDnEnCm3mWg4Eum9MmMLSSFwqpSw9WibZVvA55SVRHWpehg2T+RvwrldfcPjQdXnDMuvJBmWL
7wyGo16+rJTciJ3Aifggff3a/7/mXFfh8ZCtwroo0SSUiC6fgA3iFp6ptMb7VW6FN+zuEBMO0GFY
xAFPNVaK1g2RBeab0EXdAxoQGv5PcU0Lt0fa+rJcDhn5TFUz/LlbjlsFsaoBe09RbpZGyFnYooA8
s+g+XlPnoLtbTNQWm1dlHsd/68iaLrvNzQwUvinvxdqdQulPQf4dFgYABpAKGdJs9FRUT3IACiRr
AKAhHkdUm1mC8zB+oUCu6NS6tx2e5r+67wPTptyJK+aMR0S9l+Du8jowr+ykdFw0lEcLuii5WeRn
BeEz5hqvfdC/b2w7Ag7CB6QiVGcvib5XNGbwiIPUhHkdZIuLsL3UAnm/yXrCgxJ1DprKOeF2Bkxf
ZZbX6tWtdlpSvBMGWZRVZzQt6kgKBLhmMU6AzLBs51gnZfu81daU4aENzSWIoj0HoOws22AYZEqm
RR61YineUjiInSohya3//tTVQpnSzy4KCSOPAKtqdOYzmYcq6jWWpCy8cAyT20/vjCEmfaPdPjku
JZSHzke93JhEoFRkS7BuzWc9R+L+1GJhmjPt2MoNJYlacNOjGp7gTSuRbLSV9/GAs8Ab1/9+b6n5
M2IU8g4b+0Tk+PEkLllcr0NF2THuAAZHgWxx6aiCp540sJMH6RyW/4gzXX1gdwUcVvlurO71l41T
8DY7X2feRDPSm27pjUQMeeWT4R30cZQi8LB7ZhQGW78I/XK0PbBrImevpnFRivUI9wjXVDZR+K1Q
E6GylcU8bD6SRh1H7sXdzkYM4aEN95PCgH6tEhGUfFFQvuAElLYRdgNwW4EjoToD+QKwr8uNYva8
cBlASCe8epUzenFEhkSAJ93+2qwIQFISCc8Gzpq1V7gv8pOGETQ2yJBBr4/BLiipZBoWgPY1idDz
ZWFdJM55cIQ2kgdFObW4vc+ZYonovTSwU406+2rcH/8EzQe5j2Y/XoKQMW8KmibS5kRtLbuAWA0H
vTPdiIIfMvnD4/X5o0XVEAqxzRV5lJ4YPjGDFiISSjMnHmoKUsd2SBHtQbzfoS3fqfgH+wUBMffa
wy2li4/hZE9rTuE6ZQs5Wpv9z0FXvuyDGQi5ODKvOkKIhqcX4KO+WgbpTh+s2XlfMfHOhGmv0awG
0XdAp2SGA+2pbEPN/I/qcD2D9qmBzDp8+qDme+kHETGiocuIgPXTqTjKTXrxaXmilx/WzAUmkqsU
fi1eigDtLCayyCtBocTIc5mhuXW4YvP+Ho6hZyRr9V9JaAIf9TL6EfvXG+Ys3S+qoeBpqtjvAJ+E
74htfbn7nfjkxbkCRoFaqDF2Hbchi1ift/JXwXcymsQ7qwKw79kqOkH40Ofl9NwA7LFZxa0E+rmX
yp8x9oz9t2x8X+M0bMPFF6xzpvBlJUP9cd+vOxTwP2Tw7MSbKeld9p2W1a+ephbkJvrSFGdf2pDt
V9X63+O1uTixYDSK8YzMs5FUWaoMbhEt/TLar6SBRW2AIlL8O/lkzeJQoqmhW0t1TPT4o3IvJVrT
jz8gd/v8TMqbgPjTrwnneiOmFCaNh+8ipOaAJN6iIeQaasKMPVLca8CAomRF8aWPRH0154Psxnza
CZyx9eADlubhlb418qy9NdyMrXhLHVcyS+ozexkPFmUQ+ERqqvwHgDskUiPzxGjzApAVLCUFUTnC
/fPs09sv4JqFFtlHakTWPxJfQhcejXWTANCoTci8KxR1lgayFOCvBDgab3Gq4Waw6edHL5zg3Jzf
SUHsKm5/ruUc9B4sXFL/C2ucMi3XTBdlslWyOlE3okYN6PzPIjUJFZrChnEFrVOPV7C3ccvrqJtc
e4NTHuZfhOJDep3KnSQb62/3DcwAU1phG+GtBZE+z7gduFE1mLSN4q0y9GX4+9QKykVHEeG6UrvZ
xXgrDPFyWZw3v4LfXwztUC/0/J4kP1sbyeAkhfWd1i/C6AFbVVjZdRVOPtUTNPDsFFjEXgc7PzH4
pTOB9Tkm/8N3VK6Yh3B8q/yuvOsSUPHit/IuyC21nm6lYxuyOe0ltdM6nsC4r0trFCsDz7Bf9QNh
jYWJvLJt8IeaALNr3NZUuVosR54kwBwxI3/dUTsM/PD06OcF5At0/guCprwidEObyI31CqeqFagx
dMfnVQ7fEHCRlU9HEB5ZF+gIdR511Ay/K24DOyw9RSTjPKcyFPQkHlQ9xV28VZt0O0f1jbn7jtnk
nmCfozBGFQtUF+cIaf1x/lQgi14JkGxnd6t/fWlqrS4u2XbodK4AleKsi8x/1X8rMgDkxDKCYgfj
PUiw32G/+NLLpaRwyXq0n/NvCIL/To11CAOIrRH+C92npoOIG0jvbpV53/fAAdZuNIJqTmdLcIYq
+Y7Hd+A1FiiuYCw1yPS31lxoFsA7h4TN4dno9vfD6tFGp/WCdOz7wFJd3HGqp9FvvVeCxBppVHVg
mNGvqTwDNzUTUZdFdZMpYeZUd9zfyIAVc3zUAU9ni1RVTxxdd1vy4VcJFuN2ybR4NchULK5O+6w1
hAPbBoROLGSbjHgL72Bq7kWTbd/W0WuNHVDm6XbSpK+I4Tfsbn0oks/zY/SXnGepogHmsryJLpCh
Yo5Vvfy3JNa15DofB+si4rxz0t77hB8ijq1MWVNFrtONFRu71+vssv+mtPyR2h9bA59igPiRx/rL
CylSQQhkhAH63+a+/wZ4wJ5XSk6N6itBAtOOJVYNTGQ7ku8E83+5r8bhWqe4cxU8NW9doGc6I+y0
J2T8qs3wFm2l8oCg3quaB8V/r0CnqvSSEaWcmZaihSs1DFwUat86/PGoAfy5QIQgfQXg2mwjG+/F
O1WVB4KPcGOyI5oFxzjS+P66TK9+jy4btU2MXGruwJO5i3yzF8ABfOOJN6wUqbfxnthchj4Z8z6b
gUEQwSsaNo/Ly3FFPvclZ9qpOmxCILPK5QchnJicGDdUl92V9Gumd37tPrinW4NUZI1rR3l0je6w
Celk1u4T8Y9GxYFqZSm3zi3Yha6LtnII3UVNR7lAFGy/jMiZ+7EU+4lIaNGRcgaVx6ETpXj505GT
aO7HrB9hSUW+9gb9K+PykvobMVA/bL+l8BlNZNqUctmKAKe2T6qkX3K/nGUygJh22tDe3minZFZm
ywwWI6XxqQhTXg/LqnlTgXJB2QCTntrjh0927mgViP7Sy91PJlj2phT4uKUK34zYkMsc34/s0LAw
RBP2JpLyffqg68oLuV5No2p9o9EtoTA6NDtYnEMKEcmZ3bRnLIWIBTABXwyOTXWLqZBj1yXESe/w
a23ymwfwJDRqaH7vqMQTkcvhlNsOiGMR0VYUtwVEhY16WPSTxveP5G+aBqKfrZ13L5B4ft0H3IvB
RhULLqwzFV7e/Ap08U5TyJceadFqsABCZxMjO4A7TDF2AgN9GVfiIsp7uEfrTiZZCd2A1XS/slZM
KeWnEnkwOtn3y8Go9vkzPT42PeZala7AGMWb/0wnFrPn0CN0MgdweUjUEe2VuHrMUB9Ls0IlWOeR
gF5ODyb0V1t4uonmLzTbwFhLOt8IyVqt5i2mpUjxzMVCA4S3+lYPZeQU0n8VUh01IDhFqe/bv4t1
svO1TplC59YbYNXZJW5q/WYg2HysJM7PXO0c9woi/9xd7X5bGlvG8xhtYSUw1HGCdSEE0GfMNWXl
QotgJJRix0K/8/kx7VpAwN5PJpQ/NNynKNLOlgcBPLUevCGdCcR31cI8gSZh7H8UwM4L8Ehxmkii
ZcghCrmOlHP2vP+rWB/SaDNEdv8Blu1hlufrwugz6EvEpz30L0L58yLkaZiWk4xAyomUDJJStu8u
ky2HSsh+QRJmu1CtklXhadQWzNY/D0TVcotBYnbl2UaLC5WKkrFsV5k86avzC3Vme+GVNGVZ/49l
TGZCMsfNT+576R32hGUK+iKFaHawAKSbWhyiOdQ3W/3O5O4TDTh5IQbmS7PDQUhDJB1NNVl1VQfw
yEY4dmlIJ/t7q9ED+XD0SJJA6pKJPN2utdqHRpOa6XUv6iSb+XYiGTGSoshraKKEqwkwOQlufWVd
aciSoCvikBFc1zydVNgKpriLw6ik4fODMzb5F9AitJrn584Q6hHBTH9Cjf+9y0BFyrOJqXDPSfTO
4AM4uFMApytYdMZdED7HVG2E/sipTma8OTA4bBc5QAs94pxIPFg8r4fPna4NFE6avud71tXvKKeL
pT1XNHA6AQw6SNVvyDzdmeTz6SxuA2yJBcOFuRfZ3lT+ZFUEvVuOc0XReew5NP46OLAp4pazk3vR
4Y0GNAh20hoQPj4XS5pTua+GyKMNwuk6dBRSv69ozD526PNTmuw/rnmWw57SH13rCGYFOFQ0zM/y
ubtUxHCkQ6yvpeZHaqE1dvVWQSyGmJ1OBXJb7HppkBBeX4pAoo1fG2Hf7wPr3/3dDGU5sf67Xboi
aPcent5HdymhzfUXjR+gv5+3Gk8Z83J+NAPwasAA3kGwc6XKH2mEi1UA7pUmUOSA7amP83rdbwHz
a0OToO0aLrPscoRxHYpARmE2kUizhtAL5weWtVwdsk+lNPzTTlqdg5Zj80gMHWSbH8s8q01IqeXN
7fjYzYpwLA09Ha+8u6OpssjqFkb+tT+Ru0kn2fRgXr9ZGlPJj51Bk/nZEboFDR20/BcyFqRzEW4o
HjBoxakgO9/DVVyv4gSxBaPTZwpSXVmEyx6HGcaqdY5aYiQJhWpeQ4/AhXf6JBo01K+anBhKorGd
jH5h4dE8axu7mGEku16ca4OJjXcUEWuW5cWBsw77qQ7sIfAwxOtiwNjPUm7mYtGb6F7X+nFYl3w3
d0KaHNLECdzZOKGxlgxc7MzrHzcJ7LmddsKl6o39xAn4aqDRaOPBHOLZasOU2m5t8X4wAH6h4LsG
+j14zwNE5ZxC/UuQPQDJ1grjTgZualeIvsc3U+IEhR16ArIrRbGCofODDZitnrtqHHKpBb1YtY7Q
dgMK3sOuUUOEzRN53Wy59rTEVNyEmwzp9tP4wC2tk7npZOIL4AX/YQFHcOnbqpchAS+cczULyjaM
t+SvrojQyw1+R0XAinsJFmJ+hEp0vdJHlnOkfHZ0qVLwI+tbvd0nKmnBbcgMAyGXcGHXSzFv6get
KU/Nwp8qHQNV3vQ38tIu2P/YpctebYq5hvCaJWG5jKgsEh7vxBubSe2+QpbLw3GyLCEV6l7b+Mew
poWI4ZNZKMPUncobVA+gFxhBjpsWx08t+AHidCYqw7qrvZeSO5zR8uIgYDvuSTiOexDK+1n3sE54
K9P2xoAcY2RKgTCUDaTCh3f0idwU7Tm8NzwwPFnJnqAqQveKTEIN9JNaMir1A1YRzBG+Vfcfhtb9
8zBBx/AWQSK8ADPWuYKLn2rqnsUOJXO12izBLbYIBvCl3aNZsNbEVxKayYwIoPTm0mEE1pKiigCo
qBlJLWcBRhVpiG0bH9XIm7u6xgSwmEvsYkt3ZPdudXOgt0ER7fXIwtAjRZl5xR48AQYV/G9NACwd
IBu0d4fzCUH6Sgldegjw5+nRAyELMF1vj32+uoAKm1xoqvIAzovvTrQwEjYzlIYoxVfokCEAHXRH
DastK2GIaxoZHQFtZPnBgdA9TusqHiKKGV0ZpGOmJEsRY3QPcJ7/oBr0o1SncSA+pVc/vHm7RLAs
YOu4/8RaqcN629ET3MNUXxEPhFVKfbrUCFjJIp2b6fTcGkZTf/ZdHer9q6bQ67wks49vfHGNJEbN
Ni45Ui+BGJGP+qQpRKDSiXDEYhjY4RaOXA1YRW0lhytEC/+1FpEhh7kvdiBnyrJK3e1GBI93Z4I7
F0v0AE/wVG6QnpYjqsL2lTDH2eo5+OTn3wEfNar/qoLRDyQskUuxCog7XGbDOTQ5VXu3J/bgR0qI
ZFzxyY1QGxOBrR4F2PiX3EtK0gR4nU/i9cnKdFX8msNv6tmVeiV/kvWPFoIIJ0pkJjA4YqUbdXpE
YY28npcR/Dn76TERYGpW6J9oOtYPO7aTWIS1dBNE7V9DksjJcbSv+eUa8hGxE/U7RrI3W9LTRRvz
bTovNIC1tkjoLv0oO3WADGnVD/NEHFb1iBII4YtqeTJRw5NxT2t2eKSbMRiZvGcxb+5mxDdmqOXE
AwIxBOKK/47vev7uvPm4gsufLZa7eRCsGIuitzJGrh8Fz2v6uTzmdE1mFHvOxYucKvzV/28bqcwi
MEUWrgt4ShmGbX4aO25Q5UmwnnR30q6TIjsI8S6W/F4zk/XaYYJcyEALZ+33b8XkHGz6jDtn2HON
YyGaLc98kCEvhVPfSLChxkXFT8+gsPyUkm4Zh4c5+eEwnpNhjasygE+IQ4QMkK45hQu9WSLqL95K
OVeCjihGuG759I8Fv+4uKTfA/xJevSieKyjyOT064EV1DAiPA0a5uIoa2+5DYKbeuKYKXOYpXNon
MdpV3fzGmWB09YrEd2Nn+sX9TgcuFQyF0/PPcTaVBer1hroHe4vqAMdmzPl0N9hzpJXqPQljMAxs
gnA6xwXWX8oJ2vzBhvn9YXVzV5y+MOp/pgt5JuARs6QA8vjqO5IEBtrmEt8zfjUf1kh/qV91P+qJ
ECfULv/d1voHEkseTZdYVOhtnHgesB68/M3JcsmW+XjroSKiwTcg3kVZ3ksXOZNBcNBnBUtRsaWw
X1LhLtYw9A50YjbJhInKJwGF9UD/vApwe4UjA6mN/R47qXsUg3ZfRv0tjRNnlmjTnSOcFsWNeqHr
QxmcE9dKntr5YhYqK3AzptKPSMovPM0ulnPXBs0eSaE12+SNcggZtPGaLvVAeYgLblAdGCl8F/Ti
Y5AEpS3d18gWRiT8vktpSNjk9N6ITamWzETEA5gS3EaYu47p0ItEnt55l2mg3UuwEPIDmS1vxd1Y
u4/ZU3DQSKkZjqEmkLwj1ulL/g7JOJHN/aS8T5OmZ5/Sj++8IO8AdBZO7pDJyJ3f7txUoQv+Qi6S
E4UG+WSF3g4wN95zauSDNGFGBkF25VH6N0Nn7nFJfpzFjVCQZ8H4qo9qAzNiGX7aGJGraQLsChhR
8d6aD3qfdS6MpNA1KaIFRaQNzinCNE1p2DfgcxZM0xawWku9kQWuNuQvgMkfmdcnpseyybs66fNW
wlrVcVgRCJ5RF20NIEr/tpkupTfVNt+Y/zE7qafyIpUdXP3YlGlTiz8Jbpq9JUScDfaS7iK2CXp3
2HRh58i2iljiq3ys4eRa+HDxqfz0eM0JQaaHrauF0lJVWk2S9dEt8F42uABzGY2dyhXHHyetOmkd
LupL3Akfo/UyogXs712g+a1UFInMCU4iJSUUMHXK+2jQ5GPQ3Vk2IHFc+f4NsZJ/9BocpF5t77pJ
L/3eNWYlRyt3FzQ60BSh6EUqJ8A6F/dSyzb36aP4njXUM86f5J7M6EXJbbdKAKIB/sr2PHtJyXyZ
iaFPVizQ4iM/aJ2UfmKOO3lPSSQ59EqgZGfT3NI0niaUdJc43V7D9KL7WsPXCg50clUqJbjHPFmr
jrt8vfX1ojoJTOUfAUywMHwEMTkk2joV/inyB3Ou/QCkD+gA4DVaOpNu05qNfPDa2VATL9QzDikb
9OBpxle6Hle9a3JsfNRijlh7dyPR9znjbuMSg2nf50YHxkfX89MkNnbkOOWh44/Xo4shDAiJtGRI
hSMpN3puo2P4lxwLvpxa3ADaLDbSvS3bfFkulOsZ3FJ1sUVxtUQg4RRqro20Llggc1swMgo/fOCC
6PdDCEza5YAjmrEvIqSXTEpWGktzsz3EgJF02sEaZ6+hceVloI2tYuC4jGDhEGi2tDjnGe9bdgOf
lnot9qXy/iHDqvP1ndNDL8oLMKFtUUM2eYw34Zyk3DXjNvJr23vZloZKfELe5eizBGJ4oK17CEnL
PhS3//fNrjG+1Qesfj/N3Y9yfUD41CL92m5QCWDIb87PnSY2SZHohjov9REW9jUV0ZW5nGsFQxDj
wfgJP8NqsFRHWxkB1za0Vr5HZ8TzCSHmbfBSgfIOOsGYNDrtgipzvr+IeTth08TrK6dLx1xKoATv
FDkejiQmlXyvSHmiDSL66pn6LLjgGY8F+6DeCPE5vqbPB2IuIDUMPIZSlAzmh8l/CfUUEEfjrliC
rhDV0VSQ0gVq6X03GXIo1v0NSUIPDsrnub6fWUZpy6304e1x8tOJOhAnfOTuTrTN229Ylv9KW2Vc
+rg/xODYiwfP3fy6mb43aT0oOlBLMfapLirntU+n8SjvoOrBy5XWi7KS3h7YaqFHFJ32Z+55drE0
/MLgM/ZpF9lTFHmzx6WIqj0fKPicFImNaeA7sqagVvta2Ar+dbonVpv2EKA+crSoLgRS3uLJr6ut
vjQmLlmy+PWe7BlXhd3G814bXjeAkSylXII0MqUoKKR2FVsLXg4PNFyUjNoa+Q6pZyxWMCvz8FBp
ZEtVEPTtrsfAzWD79Iatzcwqkf9c/VmIDyjv/ZmvXRWkKNbl3LUIS+kV7Csw1KhzWrXNyp3PixSZ
XQfJpg+nb9sPeUWRIhgXiYiPXal8eb92hSdWahyep+vEsq9ghAbbIyug8UITdM8Y2EUZ6V++fG7u
jYNNvECXte2c0v0MJfdfTHPzalanYpOB/lujDja6kZUNv3DxOqL+9Qd6RFXAUJCIgeexPD2wzAJV
Fe7Rf7YHA03gZlyCRPjyFyP+AqEiA16l69F2Z2WahfYPgLL+wmNZuk8I2dtNraHaIYCb7ECCr7JD
GNYhbW8wQMRJsBa4s7Xzz/G8+/TPnry7FmJoSvgKlNHvHWT4sUPb9MN/vyY7WzeZ/NCC5gQid03A
B1cEHWU5RXMrUbXN4R+vp28KS9PAizGmVate0ATx07KpTIhul+k+7i4tcYS19+jubHg9bG2lDhQy
sE1qW9oVtJjhNY4qOpP0jVSQcrCtM5gZVZ24ZRtxLDriuhknG1cRYiTKRUmPRVjkbPP0kBJJzjxn
eKdGuNMIXUv0Q50e9iJTRRucqXTWDTLLlcwm1+kg3DVEw364bq4VnuOwzlZJVsIkl4DAmdxBivYQ
hYFsAIQhKUkgWMbAkNCRxkp1qeELoDibOGFm9/K/Esn/Ib2WWRblKooBHJtIStIrKorKjMVKNNWr
s43PvYoCj0bWEMCZKJcoQnGpbjomy9GYDsZCjHuySn9j41GJ87cdQCrRMapjIAMaeztIcwV5tt/m
xTV+TrXG3gpFL2NX0DdI3zfYOlpuAvPaPT9slbF9e2HT6tQodQ0B8CGgP7+uoOjeFMOTmvj2/acP
34G3hSx274TgCKgydPybDjy8e/3Gf+ewEPw5ODqDeuuZ6MVZAH5itioRrBM2LfM3YDjsUaXf+yMQ
X1hyUY/2qv73SNIe0p4LCN7GVYDC3iUVoaEIWY7WrbJLzLKB5mwGOM6NkhqC1OctSl4vwNkVezUK
1CIzvkDTf2m3dwaKrji99/2L1Hnr+T5TZDV4Q07MVAZZMbxcoq8zFWeBFvDsk+KMEYOpk57GeGCA
3HrA45HlylA0/UB4yKy27VVWNBYO1a/CzquVfv6uAqPkwDpzSZ3ikGh8T4+BGJWGXTX+ZUsY3PqN
VT97EjjbDtcFSUYSNMMJ46BJnKc7MxagAZBSe4dIDA/Wrp3+y9Y7cSTjoPf09P9rb40MQz3sv4bk
NBruoS+JCKeL5wbDrNcwsU8XnTV3Cx/vkbybNv3TCdZPyEJry7gAGErRLF0+VSRF0Q9aRl+IEFqR
h+jKgmbA1cw1Yf085YvONqdYD2SNVLffgc2cwfzZ0jnRuELjcoR5pV3Ujl6omxnDLTVfaNrcqw56
t0YT0Jkb6YSiP4o3m0qj+A3g3K5VsE0etb0dbd/6zCGveUk5UmqzZREqQgOSCKzzY5cIisuNsMhl
RpgIW0j3VhRCQpatEuyyB2x5+m8NvRo47HOZ68fdMAPhz+2CFh6ZpgNRbv67tGzHL09ac1GR8Iyc
UzXx6ef8+AJuQivnCm6Uu7gpzmc6rvJLNHLnm+uj7TTj03M12DTtWsKOq+nXjlirGM7UQ4zTJQB4
Z+89VgEHrn6F8zf/rv1FKMRuKe6Ia4X3M0c4KEyGCR9H/6XD0ei/wS/2cUvZQLiYXv6MKwBxhjsE
GOHg4CDSGcpoGrPvDBIA1Pbgoo29FPxja8iPY/2s+S526QjLiOxMSP3qLpcp2hpT3R2hlXU9DGUs
bTBrkoNsj/1NNodD6NXYAUgq+72JwySerUp9Bk0T+g4mcIQXx8kb0h1fO0PX+mS9IkBDbJcsJtpu
ChNQZi52fV1BOg3lvKYD5pLaP0P8nbuDogqY/XoJk/JPQtcBqV10xQM952yiXkb1g65BWgfCQv9W
6I+B+2LktMwaxxxEYdVreQzZA+Qw7dEqckJM4x4jDPfBTHc/ckL2GBAzv26z8OKnfD+HV+YBX5Hf
4rlLxj/L9Bev3DSwaQuKrc5kxlsh5+Om0MuLYnG+Vz6vV8g21Zb0wF0TW5Jg9TfOsSPWcnCOthFy
gyXidbGho3bH1crC/RZ+MkD+WuOy90AJQRykfnK297lLu2FNVKoOqdbZie9I7p7H/Sd0nhE4+su4
OrKLXuTUWvXPOpfoIJdeqhx73XNEpnmPlK9X0TMkj0/Q3m8y9MhzKoS2zC5x7aJuG79aKED51Q3W
VqYYHGHfZeKkzouwjJ2ATtA3Y89CL14/CgciSobVa+rEFFdoki1NhM6WpWJRwJpIKhn0qDd4I6Ov
SrRdpmxsp14qudHFdW84ChuL9+0bze8jd+frHa+vyjd8d871Md0e2PazooPOkamkAD2cbU0zJSYs
JMhBuQTNwughokhchaGt37zGAAZAN5C+DAqdSepp1RCsdxpYJIt3HVCHFJ0/cOB9L+qLxFQbkmJx
jEYjGGrzzhLa2RaxOKPASu5yZRoiOas9X03LaCKsWLp4lPTvNVWNOE9jqf4M6qfdZVpZl65Lr3me
5b8XU2boEXh1KJJ0Wv3gmA34pfgUvxetUy2/my1yrgD3QzuYigsAO5MP4Gl+ira442pkLyWXb5pQ
e6ksGo/O4aklWsHM42BPPTOZJIFCkYOprNyt/+kY3ND9prqYWHrQtp+VLjZJask+2H+gwSjOT2Ky
POcde8bNWdEbz0XcwBxTFy20QVX/7FSLMHRG2/qq7kl772k34/wVQe/v+iTHyymjMIHox/L7DRy5
fCKs6U7K3Jy7JjgCHaLG18XM0GwlM8Tcm0FjND5dBs+WoUuXR9tLWsA3AVu4kIQo4SMXcD6D+NWQ
4pYQP4GHIYzuNZtOLC0KI+0XwOPVni3Nynd56whgXnvoaksKXld9lDrp0ciQqIezlPuzfQeGrgYf
CpuPQqtjU6p2Ca8mnGaJntcOvOKovC4td2m3rz4VvvaRdvWH9zMee0gjaRInFKIT7CruS74EMQSH
UwaI79ULRzYd5GKXG+BMi2CYl6bDGeOJzrHJMAGjNEWJmmlaE3jOaH74ppIQqurGLCxfzCKd+mWk
YJNteSIuIrRcxUY1z0pXro4UU3MNAOesPJdB9oV5hl1FQAlPsShorbgNjnFpdpGyRWJp7vamca4A
yaDf7VDImY82/EX+23k4EmkfQHHtp51G0HbroixrIYmlsPy+Zj2Pw9GzVLjoKH0rY37loGUF/ZtR
aEl5CLIJXa36oFfhV68BQVfpDKqp4aMRSRf+75K5IFfdXG9OPXyUznaL+M3H6kTht+hfxIQdmN+F
UlMLeho7dO8jo0v1Eh+U2TRhR/G7yUXJSwi4HVlvthN9d0losNJAWjuEDmIj+JxEPER3SrjAPV+n
8+3Z7iEYWGaeF8zLZNby+LdMTCMay0/rP4+TC0B/TJ7/ldK8UUcaQw+BBZmWKk/1BMhZjtPHdK1g
ENVOKiHz083P/3DN0innh1h2x6D0G3NXhMpKNL/RgP1ozraqZFI+Q9I4FV24xVbR8nIdvubUWAdM
g4tcGodZjrRjNmssSoJx+h/Pc1JlfUZrYRPfzDejoaTl5YYXYEl4hoz1QaPM8PGTu3LxQZScKMlH
xIyYKMzNR28xaSX3CXk5u1DT8kaReRlaFsXaA5qT4gr9gn6nGnjovV5V7IVn8oyXglHAnMnGoA/9
7/vFtcL6y/bCPKOzPr8Gy9EpH5rLv4j+sVJWwlTmuNs1S+d1LwU2lwOb/0xOzR231FkcCwr7f61g
tTkbd6pXTLeOTGkdcruMsywEtse9I31olAmtcXzLoUcMlcDyj9nw+P7ZtoEfce/o5NDZttGsiode
pYX3xNSCc0/UF69wUCjtShazg2fFHUx3b1KKwei9//RNrV5ManARvOyx6z9KRG5CFeJ04GY1et0c
GU5XJCRr941xhIW1hp4NFfBbvUGV3kUXpLQRk4CKL/iprOWArTdBt2CuieQS+pDQg31dU9I3vVIf
MoedzjErlhSi8DJl9WCnDq35wETQ87ETGtqo/tnH62TYYnxSMLNqBSOirAg+rZzxpp2hBuc4bxyL
UiABOi+VTN+Q40zdGtJB1avQ+lwd82HEdWjnyX0r51amUos4lpxrd/UzJoWow5YSiysX4Qy4aBlL
X5IkENh3FbwbZ06bJdoyRbqvW42i+mP7mYBvqpV6K1/jGIpy3VtE88JLafeRxAPa9dJN8rN2TdEc
hjUwOSLippCGrQPbRfWQcgUE5tNvVd93l5Sxf5nks02c1gk9w/pk3IsNBNoFyPbYtKJgnKifuqfT
EPO6V4Ql6GEQCr+mcBKKNDxW2li3YxTfmnaMEgHo0YfTRmKPsrXHCE5hqmWtrUB7PShYzs1Y1SDU
HAvmKSGHupSSyf44PRmJg399LP6u4uXHCfHxdJz6DHPSHbDsIXwApA4DFJLFLl8WKoTze8AIR6qG
2uoxn8ARDrhBH3Ul23pIyy5ICMmyo/cjAgHtxzN5mbmPSfgN9AwXMV7vd6/hkniIcmL0YALVQJ97
KHvQ0lz2Wmz/06O0127I00Q3s795Utlk5FAIq78/zkgD2zwkC77Z46ebS7j2QAy/dv9nnfyU165r
1oTOHe+XfvPnCIfBWBaugEVZKBN1g2DjHwSTx+Tll0mISbBbJMDKQ9KCZGtF8apztsVKgRO3KobY
3g3kKmyLHMAtNrE2WsJv5rhiQv9rF7i/R/QFUEUddW9S1qOILrRi8y+74CW/WUqFO4GeXIfnqJgN
MZ81fzU4FNjaTgT9fdEMR1H5nRPTv/jQNXsfVK9ZQjeT+jFpanZasiXLODNKqK1QIpJvsuABjjag
QKD/5qgMB+zmwTm+75ik1efmcnyEx2HFQL7RyDowj0nfa25mqZB6WJmxngtE+eeTU5e+Evl7Am4I
h4ShkG1bW0yvHn3Ct8HwKk6bCrvQnkWl0ifo4u4dbswk75qF6pgwR90rHRQFyp5yAWs7eZ1nIi2D
cxzUVQHGbQYesMOe/8tk8H897IL6mv8FVOuh8lJT7xKjt89iNokvRdYoArkDEYU0VXIx0rsl7gr5
xe7Q+U9VPOC0UOOA22WIY9Tc2nvAYqfWTK9vCYAdGEF51C5UmK5jq4KHw1Vdeo/VG23S6tcwCG87
+uCg4kiYDuD9DyyWFz1USEDtRhzyxuJ9zdZBSdQx9o8AwveS56yhF/KpgwHuTgsuQCogwFE5l2tC
vGJtEbDHFKJWf1M7xj1fdaSsfw9eSxCNF+rD17HijmjIuGvkRTxH8x5kZ6ew6Gea9AVtRuoJLsrR
WJq3Uw8dKgRS1plMp8itz9xlaWx7LzQv2qZjESJBE/aHrU/Cs0UeByrsmrBwZBnrUUv5CTO5CcX3
f6MhGqwhKFLaVyFlLrNpMMws5oyvSW9Kkh1B8nB4TNrQtwspq/iy1kFxuhu1kPHv6AO8dQYVLpep
2LZYt5pGe1UxxCDo36fQTf878Ijkw8HpmovHCUNP2xzwubtAY+Ets1xwgnLNayaMQw1XS+cUnuWi
G5fDV2nsIgkaqqJmVFZ6U9NTFCqvps9vjD+cYdha7Xcnx1OZr4WwPx1xNIO8gBIQkbI8fVy4sLs/
GfVM0AI36zhudj3RegR2LhYdTIlkuaW9ICXItMfXxwygNF7P65fVClWEM75QnhabKe4cc5IB0p6I
Y8Bmf22WnlJFPO16eeDPzWU9VX9KJCWDsdX6wIUkyyw4C7N1H7m0yfZC3mEcppygkY/YDkqBM5sT
N4LU61ZXprzZ5khHFs2QZtmF3AFbD2F94d1KhdEJAAOgV6haqHn9ybJ/g6VtbD4wfUGQyIdeFI6y
EHBDhG7rmUAQSa4Ja4AzBuuru8A5JibI+Nfov6ny1xPAFf7Lqn47/K2NkR4SqjlzbuaR0fNN+4o5
uWBVLpm3e73/73bV54j1R91mCAn75kYyCzhOwytTD0+ESzHhS/XjY9+skJG7vlaZsj6k4qEXWt3X
T/iW8HGfRneAhNNF3WEZTAfzFg8s5j99xjLuZ6t0cKdG7xs5mHXig7YxE1srGivt3Zxk/g1DpuaV
djr+8UejmwfV1Jpn9ZAaTCeqB7lBFjV27SZeOCf7YZPfN8TN5eExAWpVl+72CRJTPjO/EpoZv5so
EiqUBnkPeOVrhTtiaWSUNOYvr8qIY+oMSVpgfY/HzVeZ7Q5jNiYW9j2qqtyKWWJ6ePfn5Lrowgy3
bYqTFzU45cVIhWExYjUla4JNOz9DziPhDWaAabkJw7dS28p+l9fNgU7kq/W16XjmuiW3bDLHnFWJ
knhjui5CnPXr7fNizo4lEJtxcgiztzuhFLvaSD84ZJMED4F5ghAhA/OySD4THn7GQtUJFL8VYn0C
7dakX712LSKUt/9jJdPAyi+JaEFffTi5GrKMz58igywGZJNLnbZXeazphOWbyeEmxXtwCitNRIGS
zhmlEm0hfJPR5lOKbHHc/8UmhRljSTh/TE63XeQmCIkmT5ic3Bs74lneJhcviM/8C2bbLOcHwaRX
2QQwyeNisvvWqhefKzkpKGsVwBEu6gm7pC23223IbW0DHYnbc7T9fgsUsUun/51AqQMmhO3gEbsB
qgtJzfU0INQUb5gmVD9w/iZ4uwGuCYE+wSEzZ1loAySGWJ4bXxgkr7Xb/5T6clJOpqkSgzpzqe7O
dgrucetEvMcusxds6R8LXx1NQxuxb8XFxlqhAfMFclL8ibTAVHjnivuii9mhfdbNslob5utN/t4o
zvNTLBLzd5yhTkK7BXy3b1PDfVLM+kg6e3o4zVzxcxVUw5ZBtVgoyNY2CCouxvnVsQ9KNQYiytUO
h7WM78za8HeNjkL8SPWnz2697jCT9EJyEMUiibQAmoHgRdCcn4o6U4KCijWKamwI3VGYIx1nD9fl
KoTCMZsUyJEDlUf43HVli8m2+/oGzQxtLXfXOSPhEXhOvF5plxfmfWU3EuNEXr8em5QUlO1ZUyPT
9quHZpZyfAHMSbDBotAmXMm2uNr9B+rEIj/S45EJqy5IaszaLS7fsufe8SBel+/sbhxZLwCwda1R
02i26uC28M3nVfHvGvo3MFX4RtPZsEvMJAYtCVWAKAlHFQcVnWtWxRXReo/uYesEG2Xb4yKkjd3Q
cJPldL4OcpK18/UNUE7ZT59zIAMIj3xm9zVHSqAwvsWpNtt7JIvzFSOBX/tfQOacLv1ZiTwy7a/W
VIMSHnFadJFypqWckYJsgTZWrPFnSBunOVdX9aPm53kEOWjiu0Jw1K09qp22CXGTGX86g9qvvYtr
OYHcLVyWrdisU5ARHg2VDRcRUMMowOPmiiON3yUbffI9giJR3ygT4z1cv7bmr7rYOkPU4ZBtnabS
w1c18lu9USJMuKP3WJYTvfYmlEcRQlhg9l2q6NPfGOre9fS3fSj8YPcBRKk6/4DaK2U/YjIQdgJI
L9MPMIXAVbHnyIWECMfEh/2qS2HBHG5v3fqt2sF272PtMYN2MuQymGUppsf8cIlSLtzyzRUFXODL
VPlKGt8Ed1Tq7E1/fnmUHeNWIkwPToOgrzKOoE0H9Y8pq06gTFTIRnZSCTLBXH03h5LNSENrzNyi
f4vEcKFStAxuvHlZP+FEHBewI8+es2H2sgAHSS6GeF/dOchoDIZ3m2oQ2KuNupoewdP44ZXY+wfW
EuLDZXvF2OQIK4KVTD/hMur68IG8izfO1JonTggSmDuXClAAXABCclRZ1hxC6DssN+zCol9sb6oI
fQ5rjdCI8spY4DGFSE9pGrnch4EmAlYbAxkpRRudJ6ozzZ67NmcVBO6P3FicUQcWlj0DLMdR/8EH
cxBQAbv6GTStKfiYpIFgCtqL6ERi3dATKpeHF6BHLfKm4CksN4JGKmtb+oAzxLSirhJFtXI/S429
n9mCxN9HEsBwlgJf8DaGLuYfx7MEgozin61L0xVPe8J6zGW7oLkNE/uUOSo6hnOIMLDQjZ4g9XfS
vxkzVD6qmtJzZ2CKKbzfXNVohCleF7vNEJmu5YF/KvPxwLE8LGd43IF2pLufs1PIIrTqxKpXsUcM
xkA/XgUI4v8RQvfg0tE5+klOFxx7QDMTT8v4PTUN3J0EGSt4CFklgJMLJmnq7xH2rS//OhQVlxmK
hHBuXDrylLktGT5rrsAVLpc5Qg2L9QqIWu8lXZNbVQUgpdIbONabXCn5biGnGFGZUtDSxKDLnHua
tJjZKc+BMlflzFHa+krgI5Fn1UwcufyNXtzjIzjI5/rvhMY1byL8hvRa2Wg0Kv2fVrwcVpF95WfT
52qQ6NWyAVN679iQzksBeUmyWGNxJnqSvgmaHYZn6mqonfs1Ikx/5i/o4TLJa/2I3JJpJLRHOtpz
UanMyhnEeryOoZvN8q85oRPL5w2WbWOoqlbaRcmPUQoxg7mBuKPU7gRI0ZTz7c5xndjgGCfdG1f7
O2AuwhpgiGniTyoKHOG9Hh/ysGkl6X5cT6slSajyqWyAeNvXjlauJpZx/4wUtdaiC9lxWYRYfMp1
BLByPfd7Lsm5RR5/903vtsV+VgtDRrzMgfUeyLVAABWb3Ql+LCTqWmmHUaVHczhY2p03rq9FZKPI
ItxOW6A4/NJUNUw0juDfc6fv+dND5nGuqhcn1QbJ+Fjfh9/a7wqc4dKDvrJZVHnxqN4eJAFauy6K
BzHMoWXZwDqhSFLKBnyQX6iahGK/omdMWd8+IdPVbnXQVK31HbGLpoO08N+Blv1d17PPDdWL+Ihz
rLFCO4AM/lKqXGZ7p2jMPw4j3bPWyxSO1VMu/YmmB0CalUkfgSeNlcvuQZfrI0ZfLayKpVGtDUas
SAzTGl6QDULlh+CCgSbaU0rsjzHEECU4S9DBrhSDAUJr6r+ezJB5Kw1JfKOrXUGE1IImfx2pxWCQ
djBuyVcvdx1yAzKAXIsE0NnIuY7CouEJkd1BtGLhDNv3EcAAYh16shO+TSt2shHHaAQ589gq2O3X
T8GY7egfe7pZjExiWzOfBNcOaoUy8nbjAha6tKgBwgNxlT9rDMfGfeiuT78OYU5bamT202mM1O4Y
tUH7Tft532Zy2uPTlqws7GTp+PU3I1rumrZPSuOlE4HY3xgszKrS1fSZloX0Iv3yQrD1OBw1mbTX
ZFdYpa5Bq1rrFpXvBQJ7mlvgnLVXSJXR+mwYwvat5KtLHVhe19n7v24G1lAGDAkYcNuruHbnWrIG
kNQSG1MNRtNsvvOcppH8Qlcvgb0bemmnB2TpnuJ+ej+EAwH/NyIbWKf9txws8v0LSYugf1RnT50C
6jM2Dkd/M3IFu+C7VVfT7i0kXLY+NOLTgHQZftmIsPSVP4W0vmghmFr9wL/1m/9RvmPZxA3hVfgA
DoMcOx5LK6FBrvarg3oLRRyz5B1lfb7V8RDD6LPWOO/uCUYYgO48T9kgJfNixE2Zw98jaOuVQ0qQ
EhxKmNSs45Up0CE/4wvjjoxXwqUkN4gubQk+bJgbYJwRe9+5pZq8dFvL6TmG6x6bpZBd4a3IvVd/
HCYiNkE0QFhNjlKCdrGMcJnBtLGkG637xS65niHssSWH50N+onr/6Ld/w8YZwmWxVtBYJ+fBFbUf
Rl+qiI2H1IYu7X3FzxTvW4BgtIBXwG/Nv8QU/ItufcVv2vyyWFiX4YhvdC3eq3EDVW8fy23uRE/g
c+xykvNk2qg2Qpok80in2xYTgvhkg97Tg8rFyhZ4c3IjSGIIpCJXemqeCIymg4BcHumB/IQYaR47
92gK+ERHbNA9AEJlvBPdqJRDZ9EuZ2ITC5+pPzI5OuoFmGkwxHPv30rfWN7hENc59Ixmw39FYMvz
m+/3OOQong8haiiL0hrg+RbXvrAs/auCt4AR++wYZRVC2dnGyaB9AathcXdmULlqJ8ebEi3ueJN+
BbChUViI8l5H5js9OGAfTzW+3T3Wspt6HX90/aH3Js5hOcEs7z0aL0WVL94HuIH1VUwS21csot5B
9cjJmqC/NZveOIrLLC2Mrp8VnAOvNOBhjniKHiT5XUgeJUWIy6ZEDE3SmntfIXkDoFHbTRcAmknD
s2P6XpXZXqDSKEV3SHn56f9m6t2dAl9KF0732ZXNw0twD50pKxvO+uAirBwrF9+EIqRQ1tL56diW
ukh+de5TDdTMvMSFiw2wszQdRByjEgCtJ5DJfV5qQG+0A1eBPGO9Ktk1b3PGxYCUU7UVbSmjOhBG
K9mzKGm9d7Hwpv1ty1xwKSOjFKgZ/W4fAOf54NNUdTt+tvBcXxwvs69hTgIfMk14jbXRd91XQO/i
/trasGkJgVJrOqBhI5ssFUcaY/c0pCmW9YKUpXJUDYoKfskoP0AhdLFrQL0yM40lAoZhNjq0DFSL
zOSiKixROWNKSwQhxR8eJf0JbHWwXjHCnwJ11Z7IkQ9YGaxrcFxl5pcyiMg3QuOOb1HkM6RBez3p
fXrrQBmmzrHRSKFJnTMYn1WpO+3PRKO5V9CUqYe+FsHY+KAMNqXZNKfelF1acAVp9Ws3/C8cRltl
pfbl9408Ll7FIs985w+e92eTGlzBdOZAF+lc9bfefNIW9o7LvG9Rp+mNqOJ5meyL9who29lsvJtd
ZoUFp0k4BrP6ZE2lsfhJVwz+x0d8nf+ge9P3XTuJMfyttFdLy1XRvoOMYcCcBjpigSiibZttb/oZ
xOOzuzMDCVpS9UlrXiD42e8rSWRW4oi6PAGtuDvdl7IIM4HI5aipFZy70NgWNV0vad5vWJozN7kw
qTtMnulYsVqGdJ4zlwxUdCieIy4P28kxN5QTe14hxqaVyMENHMIKq4LG6wTPvinaky+nnG9UwWM/
rYgljSxZbndizye6rozMzuKAGXUmPQo62TQSY8kq1AgBw2tVATXOCmt8iG/wEDR3aFKGYyjvev59
juVhPITYIe8AyY99Qv2eU+a9vJ5GLRLYqFNz5CwF9xCZ3p0S41Q0vWnmHjAM/BBB9LpYMy9GcExh
hCsfJlIen8+BDXQFa38kpVKQxwxMBUmuQx1mnMP0KIo+zH569irqb/pGoJGLAU6jMZqmrXgZy+sE
47R0Za5mGQbnLWcOdF00A+m7H4lKIbK6kLmR0Vyf/6F9/ePdnAe2IsKNFvzXFAohOQd6Qc3BqbTf
HMnz72cYnyBxWhRNaDWcrFlkDaUsWRFC7gkQ1g7L2fyWxRYFRl1O1Aa4vXlyTIdSBKBqZINiXiOi
jIAIrlEaKkei1aNfNy92Zw52L0kJ+IKr/aKPeMc4+poz9Vj/U85xzwNKzndR/TYKv1LS+5zaMnCz
g0z9ovm2bavYjhpnR+MezR6wgjlJx59zFLKWAtyE2drPVto0BNYxbNLsrMTTw+S2Hu1HJoSEfuN0
gYDQnz9mlsB/zRoKBQYWvuf1OegYpQegDC86MHcYu4dTOv2rvBJY8vx1uiLMwzOKFaeCcWIULfoD
JT/E/wRQ/QS1D8qOzInPT6Gv6mcfms0v9t353/sPhf5m6+WC6vJamVmZHRIy76UYRpleo4SudR2B
X54fYiNr/8FUBsCUJIjTzRCCMn84dXfo9wkrbpGMFq7S349FTuO9+0eeTv6Nr/K2SvhtDhEuUJq3
lqueRYKwDy7UGxx0i1/EH6yUW2BqdVOJQrEQcUjJQbEnL+epvcc6KnYILEFAXEsSxQxuy6pmWE0A
wTxHYdiWtaPAT5UKcUNmKYbk6dBDA59LraHeQEHGb6wJMdNK3bSlVussAqkRGqHflK2wZIR11rBv
JZTRcUuNvp+fnM32Pzc2GEf053yYirGdgJQNagix/geuqg0igHGvCAnlc+NkLUOqEbUCpq5J+2TM
cskzTmW48pR3JabtqqbQc8gUOgx2iyBiczRcNlRaOXl12u6JpxwdczFleDFC4mDXJu8VNoHYsfPt
4CBaKqgSpCUc0Yf6nJYIFZHzkA5uRGuxwN5aGyYd6WT743AHK07UgKl8rzwrPkfsZLJIFz5iWoH7
e6A8fTNt9EhRr5OsWAe3lZYjRRDPdT1S+46Ww/9jEHPKPSVQwuWl6vF9PZCLyRKtqdNNou66LBbP
AcLGLMBSBFby3QBRPfS3WThI97p9syhOzZ6/K/OZyOXxLMhNfrIS/AiRoqUVReN18oOji4abtKvl
8Qcfg3gKLmb0Ne/fAlz8kA965xusiAesq0BBNVlRl3U2tC7ACQ8b5ovd34TopG9tILKjmZk1LVnr
qrv9hRQ66DPnylU/gTXvdkfkUqE9lbUkLqHjE6wn5ktoxA/oQ4fuazLzdPD0GcIBqHmGudROlSvx
ZLJ+T49d+v+g37pLrqK/0I7d4uvetmw3+I0QnQDLeThfDBmI0dbhZ1cG1ZoCPZsBhffLsggzrqop
RoCBW1Ozp+OIRBRi9sjiAiEpxcC90AHbxH3ASvP81ekTLEir6898higXlm04URIRm+lGwjgPdGbt
ZWoaaBnbpk55tcCMiuF4LGU4Q+UB86Aibi0R/Hbq9/4idY0KXCd6WhgPVNMa/UUrZ+ekD/nmftTi
zZBwxh4DKfpF5qwq0rZiALxm0v9TT8L6wxEZGMQdbjwP2CcUOVmPjRvZnPbN8iIRvP8HupHWzKxC
1pKKhXMGFV+ingvzxgNWB8YziRaNAMmU0Q+cweXl2vRUAyXYJNAVf4GzHlobZJWW/5iRyj4cuG8w
mI2U5zM1AWsL2onXl6XGarMtiWESqTO2jTYKjtC4OdgyJv87lcxnD1yXPbRtql8ZWrOAsS/Ysjxa
AFFiQ2PB2eN20CiBWwFw5qZuniqn4hrDkyyZtfz2+jL9rodM+89Q14JOEKv2WP2fb3SRl5+ls7zY
S0rqQhIo793diZrUB/7zaGC4PGbIyLNd2oxsJYxDYUiHqN3Zf7xVhmJW3Uma9+8D8P5brgFvsfgt
p5ZvFutofzmfj0o8digpJqIp/R+ttOYBGTzXI1URDlNUcw3d851SPXQLWggvz96C/VeAGvEMwqNC
zVFe3RZPIYDU6ZWshkYQOicJiVibhd9rg09gMwnauXrU4F7Ymg/tEFB9SlI7+IMdIMRbHiGPAkPM
DsOkcQAdmp/MQxxFI1HTakYdjtULF1drCFN3SLWcQwANt7D0ZrlwZBxhxOldYZzXdM54S63Q/vUR
/DV4yFwjq3wCBDUAFmajmDT0iyFhio3qFa67DEJeLWpqvnMbHRz6lZ0oT84XDoJjI5Udp3f5zoP4
mayXsLBgxnp28pdRFKoeaBbFANRfn/+7aR9xLSpklrAIgeFjPWI9OjPybZCORO3tZQK4fBKk6U3p
aZfVHPVKWalxFmgAW0VwqvWaEn6ItOMq1y+W3fCDp5aHY1M3GwWZot37oYkE+lA9xKoo66eDOY+S
8xtFp/m7R11GS+xt/NMtWJuPFDUhw4C4MMKU2JNIaTtoFVByRXyOLcKA0KN+8Eo/D9RFxj3Dwn9j
cVHv9q0G5/QVG2YsYUhqU6uvVBN22O5O9kEudI+WgLQVxhHyIFal+akNSNQl+rRuqVe9qT318Dh7
glFlOYjNU95Vfu+1o8COUt0ojBtv2JdnREMRLopg8/KDYcMH3VvJSLNlS8WFSaFZxd8YwUo58StH
nXEao9+aWqakjhqnKfmefApZAl1YTAPjylfMt+3IPgT8lKYaIZcmpfz3jgtOUCK+SykFZfo7Z3Ac
jnXPCfkxVQ4RCTMlYAEuuxJhScUHw5ZKr91PZJQAFg4+r0oemZ5pcrJjnGasyW0CkDbyKSP/M02B
0gxnFut+lTKby01GRl4zXfCIabj36hU/VWHvGfAEgmY5hhrcrUOY2HkUN/4yhL99qqLGxFvPYLc+
Rw2/e5koUL/pOfk8Qd/nsfztpFbdlfcEo3IP6dDQdSA2DQEVwsGsV8b/WJqKAk5+vrQjDf2OK8o0
g2hpTLGuAfvTAeG72NPi4PXCeKi6MeU3SIHvXJRNfca1ug8SjrYV7AOOC2PmVrMyAeCTsGuPYMIb
WW/qMHyWy800p1F7VDh2xyRFdfAy5FNu9RsSFJgE3jESnClDqorqaYti50BzUfXEJ0ZpVL6tfzbZ
564pNaYv2Q4UEdgcwgffdsOgdLIViLZ00vBsMu/yxc5o4pVjIHDEPTDEyychFRm+rOt40UT8xnyy
RcN7dRkkxC+Ls2UN4JIDGZqAD4YiCv5dbDmytK17RKkOlBkv54dLKzJB5oJebmlZhHfQGnR3iypO
sSu4Nqqt8YN4wueMa67r9qULenUFNBQOyeeC/mUE8pW+m85l4KtHGJsGt4yYUmorasDLSmK1SPnF
/liJFIItLk917ut9aPK8EZ89xQLQTUav18x6GSyQ5rh2gojIy76MQLBpvMoUAHFE6Iwuva900PxH
cGn12WnRuq/tjrXpqGoLriArtDi7l+EJxzkuajnGBdppd6sJ12V81aVctL+RUdYXQ+Mbt/hSDiEO
y2C482fy5z8x3ShsUybG6RYty9CLFxxpix8X9r6nxxrrCt/A8ZiDrQw0oS5k87By/UefMv4aVneD
54svprtesoGSm17J/ch4hJYuX87tkbn66R31yTnF6lBFyuoHRVM1eRAHpE/2BCVxNIr80PyELsNI
zVhzGnJdAsMoLRctTKqbXY2F1SxLfdmgWQ1663qNS4mlC2qlKK6de8Rz5pm2UNHcsbppKmDcuKt9
sLZ+TieioUohr0jptVOs/gJDqbXliJs6TCIAy2ltgpZnRItljpl8a9CYx+aKJZAaA1uJBvyAwlaV
HI0/2NI85ckhUbK2auT4cmv3UclJa4zHPdWtEAxAwffmANyn1sg8rLF1ybEk6INwtivoKPgu8UX8
DszyW4vU4cT9t/WiUR8AJzbsiT1Jsi2TJ4JCFsM4Gsd0uwwsArF7taLnw98V94f+PWrA0PGNeGjU
H0NCC5dkfwXwEVP8FCw2Emv3URWr0MWMdutvI55DgsKwgIrl4KP69JkwrPiw1van7m3DWKJfqGG1
9iUpJKGBhTbZqtNmJBNB8CnbmKj9XcNjATbFpnlAfIjs2t7fLGV1XVvJWjwAR6YPZ0tFLbkaFxUV
7k1+HMIDvdnrFoKTAav5JLtjSrHfM6bnzNvEljtmXspvxAiDJUj1aumozPXAVphZvQYf/P1jkTzW
7Z6e9UGxi3iQKJE4F+AoukyTofUG4EfG05Axqp3M7M43+Akjz7yT9j7WMTFWExwR2DD6HoGwxO28
7mnbcdubOHoYTvJm/mlqbIelrJ9+LwuJcO6X0NWxJndqTTs4d3vucylTliURJtqEDroMkwm+OTK9
Tme8PXN9Owc/4Yaxlb4MXhx1bDMujT3hfYr+uZNu5AQGHovdA7BkzN4FavOW+RpfjyKaqxQz3a+7
TX7mhUVINY6LmR7ZcQt1Mhh7Zl5Nk6gAnAORBGjMrgQjJURT3f2zMPQSzBvNXd929+7ggC1Knjp0
cZaxDEOWOGxw4BGJSV7wAYosm5TsXBVRH3oDo6IcKUPOQsmV7+OpCQvL8uUhrBzDcC38F/h4/wY5
KvA6plIrvRKvsLcLIsVBcGwpbqfoIAfBnTGxkULMLRaP7QJ78Mk275skmBzy/AR7c7GvIu1Ge4jd
OCqDkG7d5gYLO2+ntwa+UMBXn9ZI00TDzrgReUZz2LrLUYaYfw0uhiVeVrpeoa0tyLxsnQWnXFH1
oUJjT7SMS0sQVhO2c0X72uD1bkHCTVHfJfAr/x4NM9LDtCrTKSa4f61y6/aS37I81WwmIB2xJUMo
PcTjdkFmrdFXVLEVxpxXGkc0Ti5A+JBLfzp1sjvRaD7+GnFr9Tz1kSDW8rKsTxP9P6sBm8Xv4o8G
zXoqYmFlOE1HO9l79uK7GW0wE1kBUm2P2DwmYfgM76KrLsJ1xAy5RqrCRn0dq3BvA+1FN/GuIPOA
k2fpN6ejk78rjv9ty5mXx6V21KoMMA72J/0tfCZy+LdO3/k5nD+eDt9GBlcX9qQf+XvVXtYm3dMS
4g7jTus1tqKelD1CcGro2/IKFkpl/ANCqCawCSThE6ZFO0AzsnH1UNUo3VeiEi7SgLCIPimjBMJS
i+Me68Qp3GFljwlwswUxLLdOMudqAZE9pYpHx+atlNngG3VhR03Dq0k6bgQ7Yw6X/sGJ5rcE0f8T
bOZh5qqtruNK9pkqFNLaR4I6IzVvqqiLAKnLnoan+TcvFnYhzagpL0Oadc/OcD815kiyfgLPOYPl
7bAkI6nWvgNF3Yyh5aD74FWBdcvVrPtKFs2vnfDdvablgr2BtwR8pcWnNJ+a0PisPhMoXmUCeSNZ
170EgfBwNcYYKdR8jwWX12caZvz+Omf2dAIdRZ7vOrwMehzNIKEypRecGJRhFg98LC2eHTc7lfo0
tYJPNX6NZSplwNQdnd6gAjbnA+Y0rNSnTDxaryY7acrdwl1RyqSa0uuTQK/k4bkkFVuNIP/GArkX
ymyp8ecjaYu92Bg7wf52U0N/RxgQ0FITjasJjM4OzT3O9VwK/f4yLdJvoWJQmZjdvD0h8F6k5xDp
BCd3sq2Afn8VoFCsuyNaMgYGvUAWxJKr4yz+anCv+GKjJQeZW4suSksPX+I5hegP71Gp4XC5pG4u
2+O0hnc+JH6TVQiBPcnuPt8w0/BtD0Om4nFkkDzD1rOmgIB4ojpX85ziZls46he3qli2y/oUKbFc
jCwQcdOisAoF5R8VAdd9IOpbqa8PkPI4NKtF22erVo53d8Cwde9CHtv362EBBbjTFEbnElQrSWl4
W4JNRthYgQLf5oq4bND1AJy74gYFoC2Z8l9nHOtGaxLyBDq1j/CY+OH+Jt9Tx0donmJnW98WK2bk
Wgz/wMP5pCaOa+0JogzWIIftDoVMSkEv8/jbOYH7rTOX32KDSH/h8rURy44WZmm2+qAXwnoZD1nj
65241HTfRTNTkbwPUCTQayH+OuQMCjOAPW/BEC4OFuE9i26PorAklLV2JZIp4pKLRXQgftEMwpLL
0MjqbgMb9Vy7c4i7lUZDN2W9WdHevkHw7v6vsvBDbYYEwu3fcSQNeD+wbrwhCSKlbCPIjUBzt2Ec
xu3B9eIbASEMR5VXbL/x7VpGsmm8hahxEvzlodlNRVD+cG31BiYLfeAob0cvm90tMmFdsQhj587E
jCYu8gCQDsjYnlVFhZ9UA1+9y2c2ubUHQc3V7Igb9yxvfkZVU5a1erNBoVcErRzrAFcCXmJulQZ/
Odi7RQoB4pjixLo+e8nQTadOAk3qfaFsk1Hr3V8CF50A7Hu8Oh7tzhxvadHMt9LyergGNwT22B5T
iVuuRf9Ec9522y8ozXVaA34fYDHh/zANsIcEf066jC++LjgNsDIWGHZxPmQVk1BuUmP8XRahQ6LX
72ZSvpMhG6SSIYAMQ5zZvFEreX6loVnHywIoruqGhjLZD8yG0VhWBvhk7BIdk4NcBC17/l7V71F2
T8432fmfZceT8jyg3l0SkSVahbMFpANzHFH6Ccjwc3/ZDH3AJi+6o+3QUE70pExxColfRy1uMiap
zs2UtjLFBBKbtnsoXtPBygIkduzubd8xdhJlULezMI19FwI/dCANM2oq1Z+l8ck8QYN4idPCPoiF
PGE75W/WjKvdt7VOutdEKcY7ttftwzXE7iIdMj6CtgIkUUPdSM2qJSkpMmfLx44A/zFHQ0NVdFHU
CMVlI2zrnNlA1CxKoBWgPxZNoT0SvfOEL5hGtoJfT4qG/3/va9CEH4HWUe4gbKZqpg1BZlrMlFJS
sGy4u11C/ixQEq592UTKGwWs9pMc15A/krUsWEpuRH1AWJyiB5DAPvEbP9mYI0tk1gffAlCoawVS
4046OhBlrt38mA81dzNlGcntZFNRZKj7lgJ9Z0WgA+LPzCdvP4ZPyY2CFE7KkJUL+tej5sFWAHNH
pm+fEQvh9whluS6vQVS+d5QCfJIvhUDKbzRAyj/Xx2rTTavhU4dok3pP6+p90EbQv05Y9JMDopYb
hz4aIdl4UZyeorKha3buTBfQZR82xIZJWVTjpw+zDVEEbiUz3m/FXhlizkOxl04fbAFRvoxP1NOt
N8sUWgM1WSSe6B0pqUB6V8q+6luZ35KnrY83gQZQ/fQCp84/RcGjcfEeL0dT8Cw+Paf6FwKVyUDY
xSajt5/TU9tnd8jEBUPGYy1xzUrS9PjkBYC8YSZFMyI6H/xK3WO5eQeJVfqWup4NZGDFzepf/k5Q
4MKaFZqXCJvIrrhJofZYDtKXuOzvWervlHoytvqV0+1dOpTE627HeaX1bQRKOumA9cywvaoB7E5f
e9cmtDHt0HAFj0Y/MM0vqYdFOiy3jp6h1R9uNrmDDMYWvLG/xNrPAMI149YLsXs74qTDlW+AfKgT
m62zVSRmqssZSKjM96wSfrSCrqP/HALEjPx+OfdkQHtrD6OHZHgw43kktRDqXWQ6h2T7JQgP3t0Y
C3bcUzhpJHsDS7l9Dw1i5W/Fg/podAGE23uvvoFGIAAv2OHokWiUiuZc80VcD2+AXosWKZRQfuDd
LVg461CTXSTiP01l06aV+jTVnJtQ/n09VS7Udil3Moa9tBctCycu5N+/5dyZoi/pzkTmWGQGV7kw
TDGewR/TpuYFvcELYqh2q9t5WNCWPLSTB6n9alN74eplrCRA/Av8Fj7+Tfpqmu4QLSlPH9N/AJl+
0Vl9Pi6mp6TsF+fEVpngdP8x9p6LJr91veIuW9CgiQYol7IowmXwmPc17qZWHSGeO7E3k4Oxsq9H
XaI3z6CK4LbPnzAhx+Vup/yhGOGKa7/NkclpNX5VtFtMNVe4N6YLw3glRTZIhTjC4+T81N8fOa6h
47XBpHEkxdo8MaAvJcu16SvHn5ToFWyWUbcqeX88FW4FdAWW1vbZeiuFVUC2rQMQhBqgfR4llxFg
k5vfqGGndHuXoFs8Z+QGykyGVQjNvjldvyXVbHVDrw89hODve6jP8H02HVK27uzM9d+OuR3fH6Zr
2BODkbexmobgSzJjcpIezNvzDZoS1fbAfHk1j0YEJmf0vsMOXoXn6sen49+GtxcYW3+pMfKM4xWn
WHCHfGhUP8NEUT0E3XU7ovutCNYvgb7S9yftUyNnCmSaf3P9FbUmD19MfM7cZWh4q6pDAUGQvirN
aKO5H+nQpC8WfWVLr1dSO0nEYNLftDj6oN+3ARnbm7NszH9bDeIBtLqmMV/4BH1+ZVdb2ZMZHXuQ
lnx2PtSb0GfazU1J+yE7T02Nz/+HAetfQmzAOt3UECjmwa/hiHICKZbe6c/km9LNX2wdoGlRqcx7
yMsqxFeAy/QoHFizfwJw6vOvMdmfuWBcDmdPi7YA+nhSKu/VkRbYs0QTpB67QChC9M0llTDkEaK7
jN43vdf4SnDUNhL2K89SNNFUGacaHXWVTUKs8pj4IEaq/TkxENXHqK6RXIGBrqcM6MlqbNPSBxqM
5c9OQ1Z7HyLcHCOXwV4k4Xo8vt5NfdUstqMw1pW+uzU1XyyUboDgw3Kgm/aysidqMNCJ7yw5Cu3T
gbxJ36fNJe2fUHeptv2pOe/Fh4K4/1+wP1CZi2H2nadZ7zeRFwpYDRDxF52XdNvFfWs+/qnXZg6f
2ff/tzGGUP2l/NEm/N2e6g/8LW2PX3JtXZYGf0Yk0xvFctk4eeB+P6SXek5Bc5lHTEtQMfvf1WIN
HrxP9vcXOgPBnajgTBumhkh3FYGcmHmRZp0QXOXce+ZGUQoYKQ17JA5bnnxWeXu8etgM2gB/AStq
++g6SHjHp3AjCUA3dJJI8xOThtSu3M0vVk9yW8IKw+/Ru5QM+cSddwO6FKkziA199JkA/sCGuOrc
SPow051/yXu8fiGZz6TmPsF8L1hYlc7CLuihfUpBPKpdO2tTnilrVJOmVVRoqMPDHr0S7sbZPEpo
Iab+HVB35w+Mv4gFXQFX6yVOBnOdx4k7S4UG6e34kpGyjXdKTjwWKBjwc93WNqmwdtyAd3xEIqNH
dzmYyGRsJDbO+PoyhaM399jI6GVd8+YOe+T5NlNHux7073PhQjebC45GOoyocQo9V0W9/ASaQAA0
E1OI+BOOR35YJxzHpi0AqFxhVR1ZVSCO73Ao7SgRPyoFDdMjVhihXqYC/tB6xQc/CvjGzqEssbU9
dXoeV43Ex5acrRAtryH8ekG+c8gxf8KE/gQcUM0yDjIJ7UVLDUALx91ErQ8EnJ5WU7dCzK9e3Iwk
J3vFGUxj4hcV9876IxOt1YKNwNvfWjbzylM1NtkHsv7ReGlSICTWPdvr02M4rxqq9ytpGpam0wHZ
mVaozIbZUonJ1g22VEofqqhabBEMMeW2ChMwgoFZt8XCXlomBkOJWuA7WbKmVpZereTptD2Ds2CH
ZvboXv7Dmn3aWFwUcwBxY/gQn0X5NPpCKp4kGklmfxEh50fd3BNfyqRtGvulrNBuCQTSaDcb7k3L
k1jNeDxTmCtFDojjurMKdB+xoHcFHqAQ7uJqbd1chYnNQdJUc986B7MDx4QJXaT9Toz7YwIWWjt/
2O4taNbNkM0tsVXoa0/Cq/75mAwQHXhtaYGW2Pzfif8i7kg6x+hqHPCsjQACuSACj+OYYehojcV1
rFPDFeYIJ5kkf8XIRRMpCtotbqSwS1/y4+5AiCtmgQz6xalM2PSv6e48zMseXDNXfuNNQTDKGoHa
8JSpVgzy7/5/LB6gP8MJU9P+BeOdMiooOXddteibgX+fePqBYzf1rhDV/pylv5vhRnJAYP8s5rJs
jdlstCoZmd27JalnKUXvdp7URyTlkc1E3PvgRrCfWHFXvnNBWUKZh8af5VaaB+nxjY0SmgcsH9ke
7lYWZNCR708X08CDJX++gUwLv4Adv72OLtItuFpoHJ0x5suwcQLv2I1uDXwLlxeok+izqviiDUUJ
MqL2MQzEYcyha4aOFBW9DCpjlNH6pDJXohCDOU7AGRh6oDH+Fd+bl9eAm0ElK1PXlDzKaFKePpSw
FzVZfXjk9PF0jLNO9WSYJyViASfpFghC+Soi8XDKSE5X++fmh5GZOPrEWokqneU31PNZXIi/P8VL
j0IwfgzPl2T16V5CVpB47s4uMdFCVCXvh1omNNtC2K0jjuKIMOlvZdPBLhlAXKwPwVGzb9l0u78Q
+66pEby+TKCKvh8dtDuwU6I04GU0eUI4mU5VD/k9d/xedciHJWSAvZoVildMHIiwdLPXvFxOpajF
YklhFtR/UIPvfpgf8OjQR4wEglsCbFw217vo9qEoS9Cr+Z1mrdqAY673d6p/jG1N2DtIUnaGWtLc
YjIQZ0ruN7SJnXsWHXwC64Ql4Kj8oT79yXswZTkceY6mtZFYCGP4Uy1cLxMuUe/ufj8FaXCp/r+Z
Wa6EidcnWT7woRxKtRr/B4+Yoik91BkCf9TzAC3tQz9PB9KaMGaJGhnCPb5nSFkO62idijfRJK+K
1eFnGfN8hWXshtBuOKzoa49J+WjQ7P2rlfzTOXZ9EeAPBNqgJ0McSrBakEVB6LuCZmh6eQT3Asm4
y9YsL0pjdzpbBct5kZdCI/5DD7MSqGcu8RkUqYEvWXy0gPktJQM8JAf4ynQJ86vfm4PLZzMSJADC
oMtSJqgb1vHArczrSUAPWj3cjiGwIAnd2I6kpVUgpiRb0Jip/I8JM2uVRpyvd3wS7Kbf4J18hY/v
QXGI3fz+ndQzuNXccc06wnCNqQiyuM7r0YTRg2d3Fo4vsTItnu6FBb5q/H8GbfI1yMHjn3yXy96z
dJMw04P34UAkeGQ82sEQP/GgfGMONpsesjaPugJY2v2b3b5aBvChqkHtcmkR77xiTBH3b8bbVtdF
DBZaj+oOFn0oOGzwHxkWCjLBH/R2ybfu0vFsVQxrt5bR8+UCg/FRV17I9n1tFW/nTl9zyovRwCiP
AmzsvM3jGV6ljWP4HzplFkKEJY101JhtkuyhSW6wpYxOSL1xv2e3X5YUKtwco0VN67J7Z9ex1Pd0
Q9p8n1KQ9Ds7cSl2OxVd/x7H1MztpfkRVRAt0RNQ8LyH0VSrraurq7gR8F9BCWDTMFzSbZHqXET4
dWekCeFMVyZ+hTdqEjM0RGqc6Y5ubhcvvIODeBaIaXbFtEbgRNgMaOBgbdbRHVTxie133QDs5THz
PutJUGiVxumQXOSvBC2gnnOCM6+RgxloV7DgqgCG0h4CTZhTESpmY6oFSWoZ41cXXTxQfIK44DFu
U7zAlGQGnddz86UlxYOGElSlHkBAV7rT0iwEzfeXhMMUsBdAu1EZ7/IEAASCX54iKGT2XTbKSjkz
jYnGIGrNs6MAzyz9A4GAb9RmOrAm45WvQGI4P7DkBei/JOuuEEN1ZxPJahaAvPaJxPZv6jbeMiPM
cfd7XiClhLaZIafkCIWchJTz2TqEhabzx8fMJlVyvOPj9ainDBK8gC8wvz1rlyAOsZwgCAOZBY8a
o6Jgj7W+LQ1bTvEfP6aK9lNMMPiMAYHD2QmlHRyev2YnKwFN/VuCDALFq02Tz+D4VjYKFy1IDPMH
8H3Ft85FW/jGUwleW/jvUKv3pzhbl3AEyRIdNZxv2K6fUcNnUz0ryWI+/L9AAa4JPgk1GBA5yuxO
OYgFZ49jMi4MwbH+jiWkYgCgbIUdwpDVg9dwunZeXv19F82vymjNHsTbJfqhGqxbbCij91m2B6rC
kfjsDBF+sWgzJMnIZO8m2x96l51c7Tesy4IgzREEfp6NjY9jKFXyVBDLmSFUqkaCMPFXbSB8X3kf
16B94xdZSyy3DvM+slb5hSHsbSt6beW7duCtz7WCIZazD7jqdq30H5oSsc89SSoSdk5z+XIFfCWB
Sqn0gWeMtF7dyOFFQC+hghmizzNuQvJ/KsBfoY/WKT0p6TlSA2EeUJT/yDZ/mzht4Ti3NHZOGJn4
7Ds6QFou/tZdk9+CWd7tcrldveeiyH8Lo7MckcJBpDchjaLBLusPlAHx5H6THCjL5selxyLYT/CK
3q3LnJ/VSt19gmtT+cxLr98hdaClh9fRd47FJOiKrQ2fyeVpZ/a+LxzOz3eTrvh1Hb7i31t3rRFA
O8PgWCx2sVt5e78Z9KCfdlg26+EdSyZTEm7volhqOE6TU7iGAeSgjmFy7SOzYdVsG/cJcWesd/dI
1Pi69W4o/Zz0PFUJ5+YDPRpsYXIuXtJgv6vKm7JQcmHPmvkLNQwe4I27xtDJ82hqtP3+SYNYCzqb
1kgLJP4YVo0OydAQpQK0eWiRJ0pHlCa1asEYrq5hK994cun6zBwhcxSuI1OzlI/j5oyxnd7uVM6s
MW1N9q0BhD0gDxcn/UU8dXX2mUA0FqrQ9nVRa4eD4aFPtI36oMfeSglNDslVqCgVo2juzVmfGT7O
Cej9hJaCbNMRu3AYqfoHJr0A0KnaNjPFdYblc55MH0Atitf6+ZHL/BdOyj0pB4zmnYZ1J9OjuhlO
n1ZU4eYfr7wkvDYtbZR7cIE60ZdXK5XQBdcoPu+M3kVLU4optIsfFnBTgjJ4lm/7SCnbChgpmqEQ
fHsaPzU11ceffmkNDVyYwvl2mlpmjsLlwghXz7IIQjePGxDaf1OdgOUGgn0HylacEIsI4b/90iof
BUftbBoucsCrxmvnP6MKIh4tWCcRJGKKVriRPkEQMgO5dX2FMods3A9yX7oYzDYw25nOyO7YP1mW
Ov/0o62grxNeUG8/3vM6NP5b6VkxA/ORuAY6fCa1aAzkbqQR4Oj09VP3f4vbCigC+SyE2TdlQdaA
mlN26ZZ9kwT3JHGAKKQcn4/LImlVCTmFRzaPbpn0vfKl7tqyk6NSCIk8fJzxJL4dNGuG2RExmyK8
eO3/CscbgHPPJXRaUJVmu2VPPKzCBnD26nye7fEmlf2Lcy7bA76UZHAJ7Bc6n5MyUf/dB4p1KArr
TEFdE68q9DCHnDgxa2WQdbKKe0rJ3ONQ+dLyeRch0FDKV7dOtCv0uDq2IVaQwb+zGeV60BjIz+RZ
dBKtP9hIo7DM//8g7dltApr3597xPGPbvahFw1yQkn+Uv8pmtmD2Gt/osLPhK0SXp/qyo3N2PA6u
IlYtpYsmh3PWRpIIMlOeq8vxneIfgB7EYrJCsoABXIzOxdZa4Jxp+ZzCp17qB5wvdg9MbxW5Drqr
4Bmig2pXmfMTb64oWU/URKT6Lgcg2jsyEr26cJ6WQI5CX3ZqQYIojTLOQcoS5wavNyna7LIofdLG
B2xh6iw73MewEave5WiPMB/2/K3fFSGIS9krOBQpW6douMApY30yNCcs5nlKtgHlxTPbp70+v2xE
JUsDtkTRTStf6Eiu/69KPj0a1JBmo/7kct/HGtvBNNdvLsq7dUfYrkEij4dq30tsE5HQ/GANM1i2
rzcp2G8QVwRerFbpPjb0pLEuQQptUe1BZIx2jvOrMoVw4lRyx+kcchG7sihO6YP5i8+sWqN8UJwF
kp0BvN+w02ydbKh6EZCjkol+qKJgMVxIIQJx7gt4jZgU3c3hGeKe7RMK12LOPvEuy3GIp+M6GCKn
KSdoM+FW2W0pbPzwZF1EcKZMnU5DN0wALV6nq4CQRQ0E2FQ8hIyopXGoQ8cCTd1GfBpXTXwdwj2C
QYe5FN9O9FAQXtbLhptFORkujfY1yIz86ckjt3CKPqAaJu6Ig8Jb831s0ycyDWKk4rV7B4r/XueU
P/Leecc4oNuTiBZqVJ1x4/967x+ogztFp9xI8hXHSzKSO+sTPYDzHpzk6NK7Oh7cGPsz+4YtV2BU
QeJ1NwU0LGGEffsxPXdbr7Ztjh2cLupTwC7GAU6G5phVETOGPJrCUKxk2etTDTj+G0PcUwF7Y7fC
uaHMMqOadsTqhIa6sabaik4mlchhlftN9QfxdZ6NNpoguplP94m8Ef6ydw9vxc6Lpg8aWcv8WDDq
9/Ce/ScAdfne6yboTJDr5k5ugUxENOwOmsNMBH7pm5EFEP96pV9HLLs2DjmtzP4gwF4KpZ8l4Y+u
0VtfJjhg48/5b8DxEdd4aznUk/xFed9XeSFfuSVzFCyGp1nqb3clzRBlIKF8DDf491nN+WdfACaS
q0qswFg9IwoyBPK6uorMs0XxiZL27GQNIum+bdl4Xu15Wp+Tna/QT2Ng0baojz8b0d5DLVoxiI6Q
qtM0vAaNUbSN6Cu6UlITawmgrBbdySXEaRKQzz+jHCXNv4AObwoH6rh7ihlk7xUSDihETuLN2XMb
hwUu3NxkhWbPLhhwdBZ5TFE7VYOiqY//BBgJVkXzkYEp6YuvJ8y18P8XVM3YU0WmvxLtvpRNYBLo
Gyz4JyVgyQ5QWxDvOfbvQytcQNCP7jSUZW/wx3ueNg0TdYhjPhPiHJZmN8Y5GRqg0joR7o9wiNc2
s4DrdddBBiQbROoSLRs8WaWZU4RVONNGgqhhIhCyjiXCPCYMjane9ki7eYbp9Mj8VQs7Ve3LgtAC
d79owcn82hYSo9Eq45dKEb5gA70hdGZ6Yv1lAn5iHcfmFlkZQWKzFvnlVuwAGk/7kv9UMvX72wnp
rymjcgawFazrIFp0l49KxBANsl3xyLkZKWmhDX4pqP/Ec0xDoTeMMLin3jXj8EPrP4gP6nxAznZ/
/EgCiG3R4X3gnk8sOCiBGBahiYTZvvuwmFEDuEZLRmhZhlJA/Qp/RFGKW5Oqh9Pm/14Xw+mjq2As
Fr3vjMkm4z/lX5i1rPFm6Qc9Ep1r5AnDWCBdtaPn+Vk7lEwcw4jHH9eyMvLQsUlaiXtrRFt14gZW
yK35SXXuFYELTAn2Y/5X7SsbHWmhRLGffp9+ikbhbMp4V2swvtmoJAoPzY+JVhZAOa8VFhDYdyhe
qvbyTawCyY+WqnTHIHKylClzky/0SSByjBQyl6dHpOZCv3/sc/wuJVBs3Lc5h+oO5KWlVSeToMBB
HSO56h/1Ubarioh/KkcF8xq6Zu3a+NZCbGOkaqBZMVCV1Z6rcEsMegQ+fvVIV/HRx5hIoIzlCyQk
J/n3RII0Bod0ZL3ox+XHOT+21rEwvkP2L0BEst07Taqk8aiQTwllFxxm5PHkaZ+MS3Eu9h6pJw0P
7Y4mV3izvMNgOsz97voRlEN+xLiRVe7AI3f0/g2tIx+KPyhQ6pEHEeHrQAgNL5xfuFX7kK0zBXVn
CAKlDIYf/E/8vaIs3WAxUVHP7DghMJrbVRcDD99QcKlVntFCFXlTP6LFb7m+QuJIM54BlN113tlI
Xl2BULrKAV7lwPkDzPcZ49yWA/RcxZO9zXq45jf2qkUNPJ2OHDMJkSof2GJMoSAeTS/d+GPXb6QW
IaJtie+5u6DicleYIhrnzt98svcELucLhDOBq7mMw08/0BUaO6wyKHwYRTdqVZJauoKZ3UHbyTYP
v3iYIOXyrxxqOETSvajYYSsiFbHoKWrhQK2zlKho0Johq2DxKdTTril7qTrCcnvcGknv7rdLROi4
z9F2M08UbOUcEyVLhhBCvU7ra5+J/2e7hxBpwYNrVtirIisEb2Bw/LkLQ09IyRHV5A0JpX5zf440
Y2+YteScciPvvJFh7Y6BsizqNk6VHN06rrOx2Hp1sY44iDsZL9GoArNtbvtYNJnZYKZeNMWSUqiU
MAjiqUWpaXEvKWwOjNmRR8ZuFp5N4TGe+jrUYnEMN9kcv1R/zAB2FvAk6n03rfxK890dT4xy1lGp
Tg+qdzNo9K1kPJWOPGD8d5K5H8JZIx3AQdoiKw2a6nSauIQQWHTi677WKoCBDuHMiCXWxIP9EWKy
+ePcMzVSrhu5Echi6k1WCx8sssBfEMzL+UQET1g54EaBo7+ROqGByn78UVQENqkFI2i8fmHpsCz8
rc8y7/oFIqP/putG+AaYwR+iFtSqi/kDXJrpTJlnPHTG6hqXJu2Mx6Wki99yuo9d3DUx23FNR3d+
aHKV+6FAspepuEjPVN9dX6TXujix45ib1TI6WI6FTljDLvTTdCk8O6qZc5Om/w7RMPktITaNa5uc
DJLuMna/462xxgwtbrPUms/j1QKBBJ+VcNVUkG7NOUHg0wf9BQVZ/7R9QNagye3fE3c3p18OIicR
PyhWOMNgOEw7LlqaQtBCcUpAoXdz1wTF9xGdGByN3m7kEiDss5moYUhaF7Ksn8g0PfVp45BUkeKF
sHFvFa4NmJfWHXWGmAtasezt/Alm/Iwt+v2tL6TZwphocNtshRY7c1k3dpzIeroe3zphwvsr8raP
05qNTQsq8T4sQcsR2z9blwqUeXkatbFUtBfr5MN64DTiuOmGhBcQpnmhs+O63uZQufOUcvLAPeN8
M4FA7d9kihVoWdWJKjVQ9kJk5IdfIue7aEZVhsAu/+0JWFC/gJt+h1aaQhGgpXIWMFo1yn5oFqsV
K33aEzXAvMlKQYgOlkbO4lDTVfYNdYq1gc0VfaTUKRjDXHWz6iWO+LEF17j54wsy9FFUbQWjF4l3
8rLyFIC2qMc8y+sIxZhw+ze17c46A8qjz5C2I/u4lFmGfe0u+chv/DOPOytYcfi7ZVl8gYonC3Mb
4V+aTbqKQmipHODpOxs0fSQ7NZiQ4xyL1q75P8MbveGy8fbNGRjRJJU/33KupRd9Ru/jp3zRBuvU
RppHcDpvKNlnKZJ7e1iel/J5pGyTGpYvui0niva7AUu4IdGebpZ+ph84+K3wKBlG2ODRnZS9YpfC
9f5xAuHb9ZwkZ1KgAGsym2WpdwqR/XAJep6lRJiv61cDHT08A5F0gmbZefnUGaglIF31lXpitwqM
/6mhnbXQgzr+PSAC+9F7PjdKV+Cjr9zxYxPIEH6PIar3bGpcWlvIx9f2R59q61B6/3XYHbHOl0GE
nDnPNoGWQdFnDcy/LaSfGwzYWBWyJ8WiXgymVkp0ZpD+9Np2bHVfx8UQh78VUf7tGDmyA2nV+ah1
c1n3FW3ZrOw13abnodCWDpXflBG52j0r6tqP38fbzUU5Vrx93/MUawEFZg8RenQqTn0ULyX8rX+4
X06gd/wnj0cJksjMk4eSj/rMwNhYDKR8EIHVnJfS34fuetLWh3YCztulhddo2otVKL8D6dV4Ck9t
agMC7DeOPCbXVh2ZHwUsD98PTLqYSIzf78TxcaZ3cIDGIDYXLVyBGPU++I61RzCuNWP7HTnglW+2
U+k9/nzp0N7oFjo0O4SnHOWYlXxJYhxQW8jNEznL7BJLd4HzqRUyZPJBRWpPdR+n7y//fr61bFy6
xVWBvY1JYwwFQtzjTBgRY8xcrJg1CttD0rxrwUf7ov2viCwbqFeOLJ+W+km/eZh0pkcR/VT99whX
07rvuJ+CpFsUBDLgw18S6HPRlNbAosgHg/+oKvWTu0++hQxuF89Vnb6td48VT8yL2bTWLTFBVEgy
WYeyRZBXuTMqkap2QarsZRuPeAENXpUObEJVoUHFhVN2pasd8pVZjXNFj6y1n/ogB1TFv4toxo+N
5ToSSZ5n3039/+wAFuvpXL826stShRofWyBkpVpjgVZzPRc5GzO6ZWu7Q3vrsdYTk8IZRrzLD1EL
PA1xpaATy8Od1MkdYmzfsdUTY6PLAx0dWrUQEGQaZBEh13IxpNhSmdIm+M9K46O1UoGLYUIroqH8
uPDrNVKGUwFcNpG2qs8YOrH3gTDZcXZJpRk2Ua9+6Lk0a89FHhS9HhHj442/k6jiHnj8PrABTWy/
v/JpimsMS5MVN7PvTNmrBXHMslmgivQdYOjx5LsMqodc/LyH289xIBxTpCqMnd0H8wYlDHVGE5zE
cMjUv1D3jflSxfqcVPdn91zJJJFbCHvKOFPxuzhfI3WKVeH9zwW7Ey+cMuqGziupENdcpY7mUb12
yfeWBYBtL92n7Gqez9EeFjUvNI0/pa12PT0uq1BkqAwIZR623Bqho/RXqPQVWmvdkC3kwCEG3W75
4uEE40NgDSwLDXuuUQBvWYmQw9C3dJ2G2o7JTpi25dNUz0JjGqymg5q/lHfqVSwnLHkfFAlL4AVY
abcCkoahK8256SbxssG95/dnIqirQI51p6INtUhx05oq/C4JQHvjDF5Zw1I7JqIXtsWolgt2KR7u
GFCkkEjzeMXoupn9c2vKqXVQk0AHpxA0RIE67rFIMXcYhv/50bvi+NMJ/btRfPIQBO7iQPnuA0Jz
a9HC9QsdOhBxpKCmbAySPcoJuLwsbpoQoJTjX0y+jrEXw9luxlE1py/DYIBGxJIlirwiU/nvAtMN
nHtjpbglFq0Rr8Q3/zpOYluqYHKp60N6Yo2HkGw6cot6EFe76ovtwVEmS8fZT9fcpunwmvV9kP6x
fP2UsyaR49Vlf25wmA4ug/z515t98tYMGbi1p3FH+egJ5DT/BwKBU1FHnq0Gq6lIbJBnzhzwjVZK
gIdoUVEC88g1NuZvodq8wUAhT7pSIrqanxgwFQWK3uT43AfCkcKGjMc5arP+H5baNrKStS3CYlzP
GaUpZ0rW4B5xY76nRUfA+z9Fq2HJ2NoztZkCKH0fsBoIeDIprLJyB9gTtm2RmpZAqcGHg65bRae1
+2o5X8HcAxFs8vrAZ7rHzinIi1CfGq6RUkv3K/CGl9VEgWUbRlOlenJHSYZz1UdUeyK71jJJuldO
dS8jwvTmSrwxxXc+AhRSm8rpouR4piCEHdXC65XZEW58Z+X/Vq74vd135MV8qa4BTfmC9ULdB5VP
6ZtBh4zn/UMbEQEwwNOuX9oexPBryRfdT+VVlFo6Lsx0BNUSiXWjO0dUF5knOOk+H2kO5r+zIdRt
b+3JUdwQAnowAF33JxozaYlmWZN83xmQCpACSFqDKe8xlcEXowRc1oZFaje/eYJBgdHz6oOGdWKF
P+HHBgFbxadUCMrRT2FKbgHXrsNh62x072aCIfUweQKGF+nlF1P1x2IpJhL69i+SdkxATIw/eR2j
EW7fVSegCd7UbKEMP5I54JXh+HEn7RKzz4kgc58vqZOpFqvXJTmzMnahdtXPE30QNgvQi/sPTcnC
GgTaY0z7I53CGOLLxP7gdWUmwP8AYWN9qBEukXN38lRIgcThPtDO92uuhLmm6/UxzA/5hqLrdDXL
QE0QxaS36pw+ZZWHQ7AOEEB20AYQ2NyLWzCi076gIJtLZI86ddphDKrkdpeH4nwClbJ4Jcc2O1lM
gbyjIDFAVqdwe7n9cm3vJvT/96j4szxQ2thr7ig0widJrCufHgX9PQ2kYJny/WY8I8vamzabzwo9
duu6zbkszSPZmCO3ATqfBsoTf9hx8QzGAQnyA2roV1SPAcahdh2yhjuub58hh7/qGvabM7wF9UFe
MAAw9YesBE/ljyWJLs6mF2w/qerpsC/HPTxsfDYTu16t7jVmlQlge/BEdoR+G0+x+lM42ZktnVjv
oS3hhzpk+60fARUPY1DPJU9y0HydtfXPziZmYsnnTEyFR4YhN9O2zhNTcMPp8FKDOiAEnwX+6lHj
GuFMgBsIFRPPNljrCUQ72VTgkrODvr1XiZa+yTmL62I02n9KMpWh/lAhS0ox9RVEMV+cf5M8Rz3X
24Dso8BBiV9QKICPyAmwBloWjomJ6qU4RqpoAaGqRu9xTSWv+cRseMG+lyMK2yF8Ps/GFq5Sxn5K
6qPQGCHiYBS61bszppqExQ2htgKoEkchxTgSSU0MV9ogYQM0RLXREmKJ0uVkCJ9F570Mumy694PS
5G9dgviCHlFMMOLlv8ETxUx1SN8XPaXo4C5YWeH1f3zjfhnlr+cpUMDOenobGbgTcMs98zcEZN60
+jScUXR2BHsBN75JRa2N0n6pBOuZa/7awAyK9vX/SC/cKOM24DEf9gqFUCPt09+/qqFhKY4ZOh9m
6Qd7DPwozkcDYDILEmTB0LyoKjGyWxx6UJ67mDdqnTEOkQ8D8gdaT/v0idamEg85baFtMHbfvclM
7dtExeTF0u5/uMjacCTDBye3fN80ZTcGDKANmUYo0Hq54ZI+cUidI+HdboWjnMsVmGUPTICt/N02
LFr1890MlzgGrzqyuPcVmXLmB00vO0CdCPaOYRtzpGhzo4BAMMCCorM7kUNJJQg/bslZWPuMx1xD
yLsZ/AYrvZR3P/W77uBIgscexruhCEx5qjfsl2Y/UinuxS3nW1P0SSp9ptyNPvxOuYfLIwSxlezH
3k6PEQBIwwvx2KEngNXjJIOWIuBS1pzAyCDgVfc1Uq8NYsF2+GLrUEkLnBdk8tiO7a3OqI0BYNhg
adDVuN09z+4Lek0NSt5Mj73AgsdII3Toi4kiabi/F99Dgghi/uLQBlJbqr87k2g4LmC1VuztJFoc
iTKHVwUhiF1xNHTN8AfyesC8c/ygoK1ozMAcH/mWmniExV6kpz9WJKah4Hu1FwdlPScJ53k9WKib
3Cfh97kl8nbju9po9zySria6Let6ScAQ0XpjovaiAUCp8n/cOS4dNI2IUJCgRMsWnabbqrRWw+yi
Csijx6JAn0ZQsZgHBa6NGZbp2si4iCu9rC+nTVCtM65TmkxMB7HJn2ctcB00qGSxJPoG0aWj0Yuc
UZ7rflvBYaLgGM/seJQctQTnin6cRBD7tKwHgyWlDu7B0eyIRgLiFrNFf4KUD0WMKwtVp7MqnQVo
On3il93giEMGlBp7LskVrvKmetFwI8yNe/mMeP+qUbP9D1730y63v12fkuRFHYPiQA5yF0t7wTUp
ZVRZMRoPfCqnw0Tzs6MoKNpvqe1Js3Sm8FTn3p0YMh5YpUZvXA55Vs+6Pfg6kZyox1QxnsufHvBv
p4MA1TUJfHNjE+ix5GazW1aBazCuMyJTVquYksiCbNzIKPahxnGUtiODOFIPs22wph1HVVy0VeNW
f1oz5YJsmZny70Z1PE5/F87C7sMJmAqSgljXqpcyMEMmcgIOYDDLJuCVVL/b9Pme+j6l1ypg8/fQ
rWSemo8iynUa0hqvn+YLAnowCG9uw1fq5uB0jccW01ONKmcNDBhaOFH0d6ydSnqKJde0CLh9K5Bz
lPcwBz0Oa9mQTn8fVqHbByVgYRcIvLMGmZGOx2+fsVSiM0I0FhQm01xcLSTPhx2XD9vyV0dQFRzI
aFx6E9OfFOl5/NoiJ2lBmpNF6fm2224Sx9CfvBQHhwGuz536rzOt+6a/IVUIdDbnokjaPybOvneo
Mb2IAGsdOWgxvt+Tmru0hCgimH7nos8t6kJrF8Y87R3sl7mYYn0pkVGVbBHs7LQ5eBz/TgCQRGEo
hQg0fUWED8yjCwqIR8ifNEUHgEFYCES/Q/6txtF1c71IRC+gHsfXMTQEockOKkasK2AwRShEQV/Y
RpXPut5YS9NhSryBrO6THgs6DhnkercBLJJ5gy91ebxv35c9Xfd9HK+5+ElVFOqjItVUgS80xrGS
e9xEtTN2dfsLXRpEJhG9wt0cCTyyTN0Wcr6hQ7VLn0oCCyk2o7lUZrIKX9hHBwU2wXmcdibltNjO
ZZzE5/7bBUi4IMDgw5Wo6Xa/2vCFtLzgL/TiV0/sQ+nxuVTzzTj4sVF/UDD1DxzhoyHNzbIJgMQ9
VRGLBqv3z9iVbmhmv5U0bgawTI4brqLRXlsxP6rOXtbwViSpmxC3j0uVksRqvlxXXjxgJaSt//Se
NV+yi//oLJGVpvPLkyuTZ9KQfUOjBzJ5fc7yH1Fl1bmZTyziLFCxlQMARtzqwzAPNjq41AOnLrPO
4O1u5Hp0ul7H1Itw6I0502fgKSzDREnfUxztyMDSh8xqhEzzQj2pq38ySbEiIrFOu8/nQbDTboj8
mBSf4Mp6VxZpmsuz3jnLl4pLOcKryM0WIzOdzGfPo6W8HM7KihTVc+AJNmtHNxMVqC9ZOf8PCeHf
VtySiEew99/wHCZB7qA77ix5sXR8UF9/R3/prbxpktyVhrLu79PGYGso6wlHx1C0T8LG+oyP3RVi
AMACjx/ENrE1JH1rtJusdu02w9BHA5c3UErYddh72tzRh+qZmHK0WdHsZ0Noy6XpTL3qr5XVYEpR
OZJsCoJPWH9lgLK3+jY8VmehzmkNi8wILdDgNGVD7/PSKGHGearg4mW/FuUbAi891/DK4o2U0B+b
NpPucjtTtZrIS/qzSvoUzEVOEHyv5nvYeZ9Uh4af8pzOVZog4DRem2nV9g4VMg6h32LqpRgEvEEs
gvbZag9jP1kgMuzpPn1H70Z9jc917B29kzcABkzOvHwgs66iQyJNSY2/WxAb6roHLCAJgKeWfjH+
6A1L4zt8Yx0cs279n1RTeE0teWdMLYrsLEI4jI3Vjg0GoKqg3yoWboMz42QUeI9KvMg8fJDiDiFt
6GORcKy/gc6wUJAnx4OJ2SMImL/nShKZ2eWKBS0hkSu2SSbYS0tfSGlqGuSHcGUn+7cjlw9bvywh
1XZ0u/z+VFRDYNeIcCgH0cBxcK+TCBHGu2OsAucOhvqgfTbZZ42W2O/pYRzR/hAbCKxRT8XNFSub
gLGbkYOKv9+qr8oLB0UGr/gAbRgErpOV7vHItVxuTKwrhzTES/iFBcWnwBwjj69LB7V2YUOGi/ml
g8xtOf+QphuwCjSj2DACZR5Pmerv0O0RDFe6z6MqrrVvUEaO11ylNi0Q0n13/mmCe/s/mhQ25fJD
E3dzZ1lPdtbxgNG6OGNXlMMaalmhujg4FGrl6BcrVOucSWSdQmFrmxq3tPX6IqxH0/iZ41KdW9HJ
mmtL7h1L3TJ9CQKRv1PefOTIMvTS+Y5fNeuQL+v3Gk7zUSnll5bROhJVDhZNt5/Xoe+UySD8zOrx
4qdcmPcIkFSV/mm6s/dxhh2sCuT1G6+/eyHyhEIr41yqe6ovrAritc91vENOxhQaGMMwji0mgUkz
h0a78QqkHtypyKYoL8qvbN6S8kvC+Mx6+eeoGNK9ObzBuupEmLX0djwKhemT/ezN48tAa3dEIHK6
V1GmW6tJGNTT6sNuTf7l3YKpKkPlKM6AYEhnEaDuYvF7BxB9YXfNwRnACURn4zZvYZZ6Fytc2tE8
OPS1Oqpf9Y4P8BDb2AwFYWcT2d3kDEl8DY4iKWsMvvUE45I/JuxE3mPll4UhTcwf5Zylmf71aq4u
b0McbPGuNUPYTwmofoPlRI/Oxrk0YXze5hvQ/EXGe+NSmKQ9Z/oBFAyeAvVnSjXmFf75DmfjjVNV
oz+IvqRBVim/NZy1JDRpZYo0z2/Vo0KPXj6Orq9nlwjYRPVymYVGc/8MDB0bmVLe0RgZwq3Bz0V3
q4prHitiqqVFjc8i5LECPZyGDSc7Rf0QHhBul9VYdCqWd3TERE75cBQxq9KxjqY7Yj0Zl6za9Kec
yVniXWzSJnMELkyu9LEQKfbJjDfgrWZQat+gLFq4ji7+6X7B6FqvG62a9KXuX6fy6SKLlQRmVEfM
GxDJCJ/K9bKCt4wh2EpUrngmQVqjYoMtLJSn+nFRJoP9jFKLKrmIEEXfjn7QiSmwG4freKVcR1pM
yGkWiQFNMsKXfe53y2dHkn1LLxuvtvtHlxhQI3+OvngubfNjFEUs/n0T2WbiIHeLK5qzfYicF7jI
bux5rcOmXPnG1XjhObyAHQ+WNEGCEpFiNi+JI8+2raSIn3msdO/k1QAMJZ9zdxkPUzxV2X7JzSoz
XyKvTXeygG4U/7SYaqjAVxOnGlgq6pPR3DuvlD3Gk+oTB9tZ3H19jHlTg4lmS0QVGelN2RRTOrTV
K3zBSFakBwgfATl3MUbHKz++/T1K4Tq0elXmLbZlco0lMT5WhQ9vs74tjB2fl+glejZ4OFVn/tk3
fR8HggbVubXCleh/Wn8qLlM39g3lz2vj0j2cJfi5c8L5lw1rif9IUDfnix4aQ78r+P5qoFX8BIbm
xAp7Maa89poHJLHA+3kwYEIFVLxzW+uxdROW3l7S2OatdMYOR6n6IDL5RNs9Ou8pgacKh9XL2O4a
N9jbkx8zQq7eGvCNt96cmKkpzOaocndFlAA07TYf+tJ22wFlSqJt+TGMSORgK/nPh4eaC/QtKsHe
i6SMGx4kRuLTje6UruXgc5rkwlZOFXNaixJkGBjsGeMNZi5+dMF4E1t6wNIgXAnU2CDaBZU5K/ga
twzYUXCj++ZytcD0r4emDmbAdKL3Mq0FqLyjx00xpGXMxpUAQt2ZXPsYLIZNPjQqNQMsQfszh0+0
Xofv28YaFlZS07rVYoQl9UhNbZbuldIBHMbj2qxNZw4kGTotrT6RYgYQCI+4augLjkY0PicGEhCj
zLIdbnnpIRx59ptGKEeESoucaAOluBnYftu8wCeLYg26/x6AFf+jpH5pV1SnHzlzFJnjVeXyfWm6
t0SMFno764WbAsdvDs/qVaQ5LFcHX9ntFXM//dUvZTImZ2WBiTwOdj0rRmzQTsKq2kYtgxxh4r9P
xSWfp+9rhOcyUiWUUivgDVHVbcy1RhntZ9TqDJVBcHJHEn+f+t0hxkdOlVsg59/F27iGRAtjTl2I
Szd4tA26ipDVLisIg/YefRKnsYp83VHxQOaSxtwHsD5o4ciGvzWYJSS54yjfyBDEmSu/HVF6xath
7F7w/Mp2ApCeUMjb5h/3TYleT5uPNZoQMrbVFj1jsO0bqp5ZnvcdSvSJrpaOR1+p1/6u8LKKIHu7
aQNplJFwxn6ZjcOCcmb/xyeHmOVPU0ImXU+3gnz7b2vu3j5wjH8yjjkhH7KAEO+9EF8oNIDok99b
Y6JCqVwUgp2+OXGiJu+cCzmcSIzOfCiCnQvG5iAvCIpJ/qfuro/EVnOxjh/vUkIRio+mjX+WbVg0
AJ8PlFe/lFS2rKDpDFH8guEAFzoX+6UqYMhCxY3MI4tgR7yAoHzXC2OyyWhDh335jV2EKp9RccDx
DQ6EM5RgY6UfMTZ0SQma8aLHC8r7dapyGDsw6ZW7Cazfuw//fytPzYY7vDrfBM9NgC5OKi74/GY6
G8f7H5Ii9oyfqTlodGUbqo0QymnLJKda07UBaNOp84BEMXEZ9lPBDoo5Mtz7I6LKL5Ethnj9Y+j8
Dr3StTOGdblG4tFr+at/4ETrnfTGxH8nQcUCgXVvCiGf70GcF3zDEv3v6JiMP8j7Fx9vtdCAP9gN
fxTUFgBD+VTgC+O+Xm/4SJCawTaBafrlEZNq+PNCa/849He/27h2gG24HX7OO+9w5rbZYSt5JUOO
Vwrt9AYCLNVDESptWKmUTBF5Z+KPflVO65mZrIvzTe3eSIwBpf0BXQ8GnQ9o0MYJRuitBpAgtpG6
YXvKGKpV2piO5BVkIFbPy/Xw96J42wjvoRH9L1hLjrma+YP6WehVM7yGTZjIHMAd60yZqKOrtKX1
pr6bmzwRvM7Rm7sFzFL3MIYVpwTi8a8qFMvNR8R3ok8zCey5S/kTyiODMmSMuiP14I1dbfCQydcl
Q3clEylXvGZ4LxJDBQ7CKrOUuum314TuwTliVV9z8Jv6mPjNvbyGzs5IvA3h3XEr/V62EIu38cl6
6iT9hIxH/+fjOqnu4r2rJNv6pWHjMnc47qDRpQ9daTvUNmK06j6Nq1qdhP+i0bkm+4rHOQTLY94D
uZfYMrPXhLGjJVcvfosV8N6EfQauJ8tY2I7AyAUHAo9tyC3Z6ccIS6kcxDCQVEc8DkieOkfnsRyb
jdU+BN9HxFBrgQ5fT9jCVAn+EtM7MaHvP01cOpkBzaoWqyQEchwug8VQ8bpiSdnk81T3P5qKinsf
VbtuFh2Bzzin8OLJvE/uHTtnOdI09oH5xcqXJIZht26Bir8cLse2eWHOhtZJ8uOwe6ozfqPrFTZA
XKzpLgYdsYRInfV0VrgfaDfUzKRnlRZJ7bCCfuoUqAz/dxL9m7rTMBWcV3ptoWYt1YDbGhpH4Hj/
jfAEwK0RtnvcntGOJLr8xWJAnrmz5kEmb2d0nVew8+DL4EaW5ZzZTmltH0B5dFVKH39aMgdXblbE
CI9dcWY6HulEYxCcwRP8seWEzklbwjwJD8xLHWRE7b1V4sr8b7U+gH/PuGCYVuyaTK1tZjttaY0F
7+YG469bXibZiO9ZlV7tkVv7UWQm4hX2lvybjUJsRmHzow3pqoWdeH4H3G0lNSVv+6fQgZ0nYMKa
SQfDu9QqUQHyjjFUh0dnxcR6qe1lV9QXrbIOqy9KC2hYaFyGcEJLoGS7swuYHj2bQc5wr95ozwfU
/elDDtUHxM1RKvo372Ozd7g1qMti9avVyBi9/aaFuN4Ei/TT6sl98Di8MbdD4dlQ0OKkf2GDQFik
6j9aWc+ivPXktws8WyBipp5upWu1Jkkk155+db28sVam8y4t0pwA07BoZAgwiC6xd6FMKgNM+lIC
XQiSzgXuqIRuXlPjJJJRV5YWKu8JrARm/wI+RCnLnaLkYSytQOTwM5P7CHu2AdKnuKtl255QlMpU
N1TZph00GDCIotj3zPmGzA6Cm9G4G335Qi/imIk3XDrASLQqFL0OeJ6Eh9dnwY+k2z6JXYGI48mU
fUP6EXuKwZJqy0tUjWhik6Prn4XljVWm6Hd4LGKoiQOguap+GfQS58o0Ay73Hc/OW7RcojHKT/sf
t0xqtO9UzS3j8EqE/EJcHaqnDmUIpHMWuOEs3b2dNTQJHXk99I5N1HIdiSaB/2aYNV00TgZ8oi/0
WszUD2kIEq2aEh81LEcRrmDS6TTnj7KoWXCg2t8EUWV8t/Vnwuwtchr+UOAFo3a9CXauFJt8BtfJ
ZkQLXvDse/tVXNrBEY59rF59E5EbU6n4Xhyq2hwNcmpCn1reYxRWETdoR1MW3KkOHXkj+Tbhb9ZW
gxR06kTZ/oN2pU2jzJWSE1vw8frAmBjeuwduzLfapTsUWfleCYg8xjAGCAYQTC/ROeWRhpwggrKd
3LaZv54zHkXl4r2Vj1Xu2+FFbr4RJrVOPbcEuCuvKJ6xSz7N821bBnuPgb1h/Ph+rx8SdxMbLJ3A
uwXhP/WMvGmU6kjaajPQOVoEA50HlRieWUQ/9xOJkJhFHRVDFNRQCg1HOPEnAI0gJQwHPbzRGtTX
yqF5De8OJbzOKroE8/r/vt2HF27UAkjb/G8ZNDuXJuQPscGafGvVhEglmZskBZ+2SbcZ1SNNjy0a
gFp3CKFc7iz2WlxNTfl2PqnEwgwDvnaILmYjjbggzPNj0aj0X4lgaUzamoOlhHi8AZcpqAMUVdwb
95j2x+AcalxpLAYeFGHi2EjNvfmUmDNZDwhMqkyJFMgqNsBqlfOp+wH2bVQs2CWJy9FaHd0dL4Ll
l5wGkdKzx5qcbzHfD6V01tP9VF1x+lE+zDQjU/27awhWDaYgjMxsm7XSMXzcEQ5XXwjuiNa6eWrx
I83boGgUoigBv1jJKK3uCz9cw6XAlwgoSVCthytTWczXH3rvDVe/o8o7bpukjKdCfVaHveW3ljU4
oqPFCx7bmvYJ+oZ730d1VcCCqCu3bqav/mocOkDPQlPjIgNLNRfx23ANtZLncjUovb7oDb23ZBzl
Y/aSED4cvNGRcm+z52hf5c+uuPTf8BEhEXhD4cSxF6JLtOKWhG1v63ihpiyW2CP91ofN/MzeudsY
qrk7tU+arvn/aE8p867aVaxhgMPZqDo2UzGrncxm7LB7hNtvlw08h+7ptP7CGq0TkjXUDaeN4PV8
Pi7ND+4ooLb9OKCT88ljJ7uwfkuJa6LI7NmKUCCowFYn6LJZpwJuEVFN5C9kqK7YKk4bx98EGPVh
7mpua2e6zKqlQh/VlXN9FXZKP2LN4PjsdSwRFdnuAlWse+ioQCzChxqzWLxaUlaohLKCWxZm1ekU
VNSNUXA1l6ON6+qQ3FMayN3TCLYUjLsaTYb96kb3IR5u1GAchS0aKpPD08euVPmrmNFRXuzHVng7
9Dj48rBiNrjE6AMS04AH+v3iJe12/duHqI/3XBIHNEeSwujJviN62xSM6k4MpidOrvQZKQ8TODwl
9Gjda3q5D9vGGkX6tGB543xCTU6zW0tbpEwMsgboE26b43JA8qY6v3YyeEUqGhG+Uw2vvHYhfRO5
dtjmulvzTH4SLF0cpx8n2e6TpNyXi2RlmmlBz4AL3AiJtzQuXrHc0lCZY7H3I4I50heUfGrWvGJI
zwV+DLUFypyR71kMg8FKQNFZbQLcPykIv1tKHPPQZBHkcUYibHWfaBb805w1Zi3e/MRKb5oI4RHq
NUFr4WgA9kSswdM3uqBVg5L6upundnuMpNIifK3TPFoIK0Uuf6C3x06BKzD8Je+RS3ajhUZnIW94
+JZGDGazavZvyEGy6uxihTIe0j5JtNKCq3SFv9UkxCoffeNJc2HvaaKOOzOkc0iyfvEBQoSen5Vr
AzbAg6JB1Lt3GXBsJYwiLyLVgmmdwzNrhYajmB572CX2E+pOJ9YCoJ/H2Adks5K8CGFE6P/eAPW5
Fx4cYJJA4PsBrc/MgQvBh/dCQoess4UXLrEBuWKdm7OSE1pDXjazVuyHTo4FCxZ92Pkjl6A0MCKQ
JgICzijAShT+aJ6oyLC1XgstLq0c6pNrKd5AvKNHRTYr8Rc3wlS8JaztbRyauA8uzIfPT0zLpNL/
hr1mHBWD6PRSQbIyaegjFwRwR/yeEnPQyrojT5Ac2aT79NyET/2vACqJItjylXv2FlVFk7iDbM8n
A0t2ogM+mLlCZ6l2r5qTeS7U4Fza46jOKtzNVZSzX9n7H7qbRqZ/cO2c+0YU9Xw7lmXNRPQc3Bkj
lO2eShMdSty+cJ/lEXGf6Orm2iwtIpAFR572ttrr/WN8p0KC9Ip0NjWhKbTnAgb/EGU7OvQus2tq
EcfN7nXPtfBqcEhwKFHErInH3XkLfiaAmFBCXBske+ZV43mWWDDm1vinmi3Jq+m+juy8JvGiYewA
A5Xy0VcE4v1aCF1LpPqmZmzgXysfSTM695iIhG1kzIDgKi5RMtOcvjYCfGmb3BONYOgGNDIAC+fx
kspjNND12/BcosuIgPYlRJU9iXKNHffWjQ5AMfnOcVlczfUS5EjpM72r2/u24aSrE+TlfpiI151q
VZonZAW7yrVwRmrZNLJVc3oINDLT0wUr08fYSD6TblBLKnddldCS4xlpgMNV0dbE2DTWlb3jALEo
UNkmTZ9zptaoZ44UTeAolvZgXXnc1EpXt+ob5w3bcKxFgFjUoWMpQpRbG93W8j5Y6Nny15RlSVpg
tpUuoccnsyhfioet1NdoUpij3DIpxffh1uGQtP4RN/QuGgCXbO6FxL044MOz9f8Zkn4EhMPtOsJ5
IMpahpH6HYjCGYxTJX2q4VcnzlpB0xIiDAmN0nMIPtpzN6EO9/DAFpK/oKgHTfieyvEZlqrReGqR
w2bPpqWz81rK7eCHTNmziUf3M84yKaHNd0V045UkC7AEuGfqqay+pKa6AzaQrIhnVnn0oFGnIjPy
Co50NE/8ZsfXD1LdD3x8SeVIN/E4q3eK9HN0fhWSYzxQa/emmKoln8vQxpPzYMcyEpCFTVbFvCfI
qJaCXX+KgV/jk0rsvHq9rRYmQLDsBjrCJpatR2pKuelX9UfFjF6A5QXpCzKIQnQUnhhaqcSnBbTN
yz+4o8ijGDGlvvgA+eQJIXOAqKoqKEscB1l28L15zBIv73zUxB4s8CEE3Y0QvHTp4E4fYvYycwaR
ZCX8gPY8QKDAwv2Zz/oXb32RmDOY/RMe2gXe1wsEEOHzlB3PDpR0EvIQNkX0un83h/sOj3eptjSW
Kw5d8tEJK9KfkX+yajO7CRz1dudqZEdXT/kXN9Uvt7/+nbQi92nc4LNjf6+u38Kb7Le7kk5vrLnj
J2PlBceWqtzWjsLXQOGpykBcX1EBlN/DfmREUi5Re8IIH18vtfPav8hnYfowcdh9ccGP6yKrPqr/
mStGDjwuW1xdoTjwYeNAekrOixJfL2G88UTNPqIpVW2+dNuHbRp4t7CpAQJSSh6vX2N7/0v55b8r
hmVBd+Prpyi7k38hlezlBnwO4JzDlZHdoMOqib83b9YUfhyfeeSU06ELRGWRXAKCIqB4M5xkOeHJ
+KpR+OxQ5WouiX3H1hDZG2rsjZFFrz/CcvHX59PjCb+uxYi+iQsejgiQxvGhKKKAVNJ8WQTPBHhd
TzFpuPsN2DqJnSPfn3bykG/2j/RxqxxifMm95ChyPB04dB1ixJ1XKmOIpzIIFnAq1nqRlWRAaBmo
AcqikngGbuWYtxKwNJGZbzMx9eVxlPjzTPB0ZEnVklZzfxxSMZFRz5GVWKjblP2ncGSyGpy+A4h6
THkglZ4mQ45CTYV420v+EfOQnbBPnPsqtY6gQce7D9QOLgPp9iBi11zdTTe77WTSylzMY7GIo295
luxzvLbh2Zl1kWmk60yd0g+FYZDOUJLW+kh8le4gn2OnzkHO5114mlVD/DFa8Va7mrWlVRailNtw
O2tXlEJxfBGXIDjPVpp7suLQDlt35q0+WUdPQ/qenh3KGXvSexE96FXNV30a2IemvUMB35qaN4mf
byAA9wvusbE/BwvTy5dowOtWcLv9qhXqqUPGDf99lyCVRo309oCvLnggJlMmeCZ0ZhhQveljW+bM
A+gBAzWOqJr7IY2/eYWXwTptyjFmpWL7AwvdwYQbkBjgmB3k+/355TOZA6ZCWkQXICLgD2uStVlG
CL9UIkNML4MENb+cGXKVMfEV5Cpqxay5dJy3foyuJNXj5PEYccGIZb6e47iB3IAImC52vz7ViQdJ
ENVOzjdezM82P4YdGLkENpPeYIA7p3QBsEXkPV3JJIaPAGItKtiYLVCWudS/9HNwIZ9Squ8JnHzp
ExPqp0myK7OLDO2NIG4GaqnBaY32RKrt9CxScbfQwt/uoM9tF6C0aK2DPh6IYLnvuss3YWx69AL2
vwzgzyrQ/GN/z8mJyVdRhEnEALZFajngb86THVgXw2XWkcBwFw8lQUjlRwlHRTPB7itccAdZI5ML
VMBcep9kjpemBkv831vnW3pgSN9HrQgJh30nevbo98Ww5T+AP5UcvUBqUH+JhPtAT+eOv0Zpe49x
CGmki/aYxF2SgADwkG79d7gkXwGIfMUDmlUb+sTd08AF61+95Q+MHrDKGhIvScZIp9wfinoAoTw6
Sc3XJ17yQrpBfIfKKSSXTOzt/uTP9wXHtbFrDafZ559+QweVs/JeadRN6Qjm8TBJZAknml6OZOrN
xbq21PYK9fIBnBVJL/UOB+eaKjGeTNZVxJh/Hr0iyedDdsrqdhF+47zgr51mMSFowGQZUI2zz6oz
dxYfIBoP5f+siOWGRYcM+D+9zoqq2MRifqPJq/Z06M+Z5iOCkhnDXEXpBv2iCYOA0fDWImbBl8or
YqddgfMVtX1S+hJMUU0oeMUNbxuQqPkMKm6jZN/nPrhp97NsEZ/9Cpe5QFdc1s4tsDiQP/wtxtwj
1qBomKmL+yUPULM6Ivh03lkywl3G+yE5T4eXnWW2lDErsm0W87DTxIL57Gbb9H3V9Jn1l7BjMzqr
mcciOyaOThIpVzMqZzDEK0RwPtDvbnaqWvChacJpiQDAK0dqCToUUsOyKgaiRjs31nkK7H5Jtvc7
b/sB0UAGv2pwikT54FLY2fi2LnO/xSKZwaPoRZDYnnoEICZbH46uWGHyHptdkXvu16GtH3EC0kkA
KoOluRsIIE/lrLRegjMAtDDW+JGPx6bD78gPkb0i6K/RdEY7IGqlVGmizkCOneVWCH2OhXbqHVg7
lSankukPhboqafZ1HtVeIPTTdGW8Ky4KMWemiV/TFwrRESdDX1ovRKiYpQa7Blrj1LZEDnVLUEQD
Kl8wIxaKPGGKtv3JekMIg4w03ySnoBE4KOHo/x7KWhgvidBvjzvvD/gtPx+5aa5FiFPrfa8rPLT1
eN9iaFgN05kVThu6ci7nHojEjjSkjWQmnq8+Nlr95KyonAEClATBUlRal+Ycz+svcCB1IYIy4lem
3C2OI+uUpapE1Js1ZxbSW36FaTH9NlnflaH++UF1UFV10JMcP6JR10JUu0yEtiwTuWPxNpW6Dbh5
nzhJA1dA4ldaQAJaOcsEDDHjN6InpO7l90kwie+0AfW3n+yziflW8BEQ3wUi45OcVrg7wxIyWxna
J5sEg0bDaZ4qkLD1qprMuR1sJqMt2afkkYtT9wdceSfc5aFzLmNC/qLSxbneUJI5EnetE2tIh1yW
eYJLO+X3RgKuU3BNQXfyR6eH1GV2dHrx2uihyoxNSC2Vve9MNGyCMbRQzXfQpPZjwI7iFnrvDT//
YdnFzbjaKazb6fgWs9qbhVf9cIb7yePBtObdNzTCHYin3Aohh7ibrPWi95GRVjyKCe3+tN6Nb4ek
AiPEDIppcOYaTQvJ1zxzL7fxVHkNE4i36dlKZTJT+09YGg8dv1jFP8kHXMLy7EPk+w3c6smpSV3J
cCjYQgpAhbIkW59f1v04otTi7FQsRbmW5Z7PmbYqP63N94wZF/1p5hSEytFSmDJWd3h4b5wk6utb
MbNea0D7B/ET6sdOZ/EV3f2Pv+oiISahcQu39BcgiXg3TvzMronNEFtSifIy0Wk1LHl8slln79l3
7E4MTQQJFIC6YLC0T4XCDbXIrJ63Y7/80xU+S65vGQbpFo87vcwXSCUS3HOjayyjcPFxERg/dMaP
CpfcyuJhSlnW/DPLM4PChuCqoqXn/H5hEbx5UP/YPgBVvpFLNm65nQ4pEyhYE7rP3LgfQJ4cn7gH
mp7jSthLL7Twf+KCYAm+y0rVuIVYSDD4tzgEeh3yJsgnDxMGAZcfyte78JKjrV90kixg5TWa9u2j
NJdjsZYxzIcI3T+NAN4MgAmL2OO67m66l5ObFLW4W/9F+A4uV4GCrvBDDUN88loIi1fPdUWzZGg1
ADMOc9cKKe4rrU8kpJ91wJVKTds99JRLIXIajSMcKqCHNdYtZFOj/wD5tgArdibz1nF0B1SJfCHA
iYrkWFpMpHjhI+50h/VxARnd1RtYSbNjgd/8XnHs/5WPzOgfIpFlV43KFPu7yRcQWjy3o7QRCn1b
JGKnSBVEt6Pk7lzpqW9Ub3J0hOZWNKOAAOz3r3n3DnkBNpkbPKg24H9l/3xjLBe9pFc6biCKTD/U
811deq3iq4XoCociISohcVY+L9iGtpXtaxSe569veZ975MaG8mRyhP9/3Pq/H13pHIReIEtUyqLV
7E8ykvXgFl7TBA7v3vMdyZ62t5GdIMDOExmkcLBUXUyHRUa9v3OiWSrhNossReOadXkrKog8ZWC6
If+BgtRNaLbv/3RNi00eMAqyxdtu+m3ZpSPHBkIW9kZtLRdqjJ1bs3ixbz36BW9ojJgSs83fKqn2
sLPFVbPs9wWnWs0bRcl0kMIokeg3VB4nE0cZO0/ipXBz85RNt84t2L5MdEyn9HZ9MVI1zSPnL409
qTWRsY6M/q/3/5a2inzXFMb0f8xsAZ0yAe19tLdvPCQg+TCI3GzhF8bkfALOikbMWYkVUGCUeMmn
vLNympR+OSHDlG9mm1lJg1njejHVBhaId2Qb8oPAR7HTl55j5Un+URJD21wF/rdHhf3QzKRoevRQ
omKgxtKTH5UqtpwA0cfjKIl3mvSyRLR6NB430oCbTsdd68/tLDTj6uVmGNt0ptDaYIi7bT7aJwR2
Pr92+eNrh+Lk7HRZd3hSdUoEBs0Lx1vA+qBfXyZ/ctBoggFHatCFsjTrzux9JaMANwAnJvsq4hK6
Inw+b3MMg4KWiTdmWLEl6oNWNeUEzXzvkjYiWN4pg/d+RJ8j+0feUDl9AsJJpGrn2yTmPlU9gHKk
X6pNCeWx+kFc2npmiyCh+g9XJ94GZQviYXHWwLdGtSVMnmeuyxvPP2wgjA54F00X3o1uIK68TY6F
4gs62TcB9c1BNWYatX20LWRS3QAFBtNaEIUeZ8Aoatq7DmGBcT7SDxteijE27LTFQWUBRLMReUGN
RRiHE2DaM6pHCoPIA0KFj1KtFWjSJdoNcB4dV8QPKl0BqtBQLSOYl/fz5x2/+REpkuh3NX+8rCwN
vRahanQ89KkwXF+4+qqVKasAi34m+hoZCm6/U4YUqlu9HvGjygq6M4/dmqgrzCLYuiNEgbwCnZ3y
XRlWsCvE5nJIb3eTmB+wfSa0pxYubbHvEjoCBDVC0FCMw+Y1LmVgs/jjQl81+putl66rWNQ2pidK
x/Ljs9BUbDK/emOVOLgl4sbBuzyE2xQUhhVKDvdypEs19Y5jyUfP8j9UHc8ryiR+c8DNiDuiBnRJ
pkWxBO14M6dcnONsFAOewPklGZKCq55tTRqJfNUc5aC9YCTzDvelGcbddEZd5nPilUcLxsJESU/g
8wsxy+sZuTYYMjHOGh4oRkkpOF4oy1SGsmDfQoT1VxRu8Ff9Wjw6HFkXCBMPviomld1nOXo/Bfui
h2uAFJVIbzNJiyfm1H3nt4lZrvbkkfQMQ/4Lh9nxZDcP+M4EtAMxmMmu4LcpJgosa2bRO4eNa/su
KnzHbdttaDE7fCPUyMbkTYUrJFLE9/TzSZDdUCwJ8D/HLM3E+X6rpFDw1261loz+Hk9eIIbBZ9sS
zdNJ4ejb3kfdvm+LIk8yYe4ffLws/75mnOKkNLrkhx7MnM4lNsNjldLYnBHZ39qhfpprfFXFlZbh
W2fcUcsfaY/NtpDsg3vik0zliRwpiXwtLbMn+PhIpaPaTxBlJV8aHp9qn69DnemfPnXQrGn7uPBZ
erxZacB8A+UAbl3pDHko4CNMMSlLb52S53fgNjW5n+uUrgiQ3ex0/KWN0SNmba+9mAV6pCa3D3Ee
tl2cigDqKswONDpuWbqMnj6s2MIKGTQtnkbNAmUOKqTLjkhuEZec6v+RPP1T8XmaSQw4sEs8Ia1o
ng+Qt+SzY5ulbWZFOEdWsg1HXRrOVnduAUywJYez0iYhxH0xWM4nlQJljUpVC8wm5FB6novTO8Jx
XRw6p+gvuBie2yO/h3CWK3gaq+uZKcy32HvyYFul8NeVdPigi2jbWCJmsHRICEkKqEZc08o+9VP0
72G8+Uk9Lji9WO4//EoGKx2PFIL8vIG+Kq1+8bWh6yqVWWqC6xiXy/DM4B7tvnOWdiYwcJ/sQIQ/
pi/dO4U6fBFw67qIucbSBMdHloS0+YU5COzBy5XVSUvwMi7NzFITJNi1R7cCjxU0jFLO8MZp1S+g
I/INprHUsVvaKphpktA/V21PT5AJWohWd6anTAA2/+yzpXkGjvmOBxlUxumrq/qp/tqWykhv13N/
wJ7rAYzSYKeetHt2T9nVRHqsTyn/3d8EZNI2wz8ky5Ai9NeRx+eRsAu0PA5C6CCR9rUcnkRFTAii
lt3rDHke+Kr7cHcVWKrwCnBMHYEeroiC30NkNQgnguoEPPAlmmhpGhFDjuoghM+jBz+mA4dn7QUh
+XxEr3IddosfLl0X3v+avF8BN4QQWfhPaafG/beJtP3hLOAT8MFqY90ktMhYe+61sFc0Jyv6UY0c
akVNceIHgJYwne5mrrICfaRkO8ODfS1CUo7iifuiHAny2oABpRqauH8Hvg//UmK5xseS9RzSQMbY
6V99Pvge3XMqg11ATMZzsFW1RC61u2m04XC88eQXIoC2XnoWB4KRuyhAqFAG7d3042vrdbCBkCRZ
jTbZz/Cba969yCjhEqIYSoTMSVfhj890iTxuRRxZBnZ7ZY0OIkO2zo38XDevwN2TrP/Rc/jl/e5H
MC1yq7uqU05A0l/8LtoxZf37T0v0X6+9scrMvLJvZutrGJUhVhtHdOYYCUef53HLOP/ZD/wRfavN
ixETsR4zy8wSuwKYL6w1Nse+2F7iaYN0vgXR+NqkPC8c6EDW9EQzMqnOX+l+nN8l6g67qsbdhzK7
yZRQlxi3SfqOjcOmXQ+cYvxDu0367f3oW7rIciOWQiEzwpZvN9fhL+KtdxXR3EDcMFFIwFASs+Q7
1tHXroWDHUQpNzYTK1eIpoiAhTR12yg9JEMV7WNvKbdkL1x6Xhlf2XlscQBUHn7ySoEEDkL9NHZT
MQLFi1GNKJ3GBB4gMBBsP2mywJCLVdY7mqPFUfNmjmmmAIfMYhUih1xETpmxHb61jOVczlYmjhnA
6qv5K+6XBkOZl/1kkrBKMEWyHbjwDlKS15ASw+897Ah3LmoaKdhsCboNCsAGjTyEYB1YL7kr2ITF
/druWMp5Lh6WvU5Glkbta0DPt62NMA43YrjGSXiEL5U/b2k2PtDnMiBezjX6GGnwY5qKkHVAUOKv
uWzozcZgrtICN50v4V2lnKx1UefJLaQ1QS1hkVbt/OqqoMarPoGWsxBLkxIm5ZgnX7vO597Z9ue1
AQOLH0k6bn2XjfFARx+zyAM2a4PmDGRzvR6tMv1atR1cWfsdE9FWUCg3ZqRvN1g+xn74knMtkNYG
0ral2cRzaNleqRZVZQNRlf9tdwu+EWfJsCGndq59WlAgpKTmjYsfeDlo+3/2GAdmtcx7OyzpuqKe
/pH7RX2EgB0F+zR3cGD6VBzNHm84PWFEDTmHuqpH14zn29Aa2tqapSbX2H5W4Zdv0Zrv8Czkmhsu
xEHfA/ZyYUS+QSxiJcMGdicePSvoqTlXSMHPjAyQgEm4moqaGJSvoBn8L5efjwaugTDwc3rQqhGF
1JQdj1Z2lelM4kTqWGKDAI9SDTsJVaFlplnm/m404ZLYOR3CMTqdTWq9Oc0i7D4uV1zZOb1GnZ7g
cnrELfz2iOEhIZMQU9o9/pV6l14dOHw3ELb0T8JXEm2CQVVa4fm2BcPXnxKuOVGg7xcqKUcnuSqE
F83NGiBOISr0NSiPocTxJoOeYjpSBSgWfo144STfvCG1+bnSszARSmfucaeqxnGgwnBiEk++Aj+B
GCnTnum/fe6hzWX6y+I4N71ptaxhtwBYwC3WGQx80gX9zG50PldrJNQ36N7zdXVwf/dkr4U9KedA
D3aWGMeaEt8/qKij/6VajOcG0hVvc0igpaZbz6NVU3V/mODa786XlkCpiOmgQHtVbuw+RDFbPncC
kyj41UBdCzcZS6I/CzAhvCvnakBHfh3swVCdltxyPKjAQeYcXYCxOxfeAfxa05crFHnRGau8qEo0
C5NCy1AAxUiLyBG7pnwfpodd61GHaePI4FaouzDXJ4qgI7irJn5UGuS9pQmEFafYDNbBoVrkL6Om
U995KCweU9JK1xYgVJMvrS5V8foLYBiCEFPro0cs/G1Kn9GktPOcvGhPCOzXqJamMpoJUQt366Gw
it9kCmiwrhV7ZcsNlx7OFnpB1BDGRpMjiwQnlsP69+NWOhKT+BL+HmxkF1vFQAl5e3ZMayw6AIc4
tylM0HzvP8Irh5c9sn3VGhMDVoMPLNQuM1M4ZoP5/0N1FtDoTVarkwQyje85JhT4eKmW7Oq8DMmz
WJmYtpzMSvl2uW/KIf4eM/3D3M13j38k+8m19dIoSPAplaSKeNT9SOsnqdYBqI0svjOYg2hmScsN
Wl6Vjs9s1/PgCOHVUCI5C3zFmTAgME3/B/zBGCEKQwxLYUcdqHBDwYEH8zEJFC+vATimoY8byvjM
A8eD1No3gRLjBFAYZDLsJwBgzokYbHbCeVs0uG3WBoEt7Kk6VCds5YCTzeg0g2wfd0ezrG6pLoTj
iQBLIK7QcD8h3mrI7hOfjuul9zr+5/fntyKC5ALFDPFdC9UuU1TKA7dEfkA6yIMnKtXt8H/pKhfs
4tB/+5ucwgza/uxy3kMIf3HORTcSapssQzBWkiXQwdITOLhLQEJIGwqaA74hU42RsruzSmR/oMCc
+DLgoc4m+oFu3KvaNFmgPmnW18unpTGERCh1g6ZcXT9Fuzh8k+yg7Nl0oGNQeJQ7XHrcw3u799KG
qQ6mNkpV5WmQJ6je2rFhkzFWUGrnuykODhTqcB210Wxfae3WBzp9+xHMfgMbH3lQPp7xraPRdibO
CaLVdhniUkX/7R231cE2dDaLJlec1wk1MkHckbDL5xq4L2Zwu1We/O17mmLa0iAfOyjcGpAwJ1fm
Ou38mONgT5yNYv4F6noxqpuvAJ9UeRvOIci/DeJc6pWTHiu3b6OdXdhh3U/3fPIftbGjpD8zgaw+
JOHR1yPObQUvK5GQ7OoQap1p9ZhsAgaXwjqQj5ijdYcSykutDvlsw+VSgLz0p6XEG6AQIrkHDnYb
K3K1mYpcZoHNAHamsMvwPGpiN06pBkdrbd7Jd+zWx123IrFjzQs93k6nIrmOjnUwIsjkeHKc4sbS
13jK+sBzkLcNydG+dds0/cOKL9bK8oqcDw7G6vjCqzhYCeOi0FeHcjNPdUpgVPxai0Bv2K4Pw4R6
8DoXTej47GxGorVH8xspg37dKxG/8rsA5HLiXnN7wcOTadhCxPdSTXgW5PcDYNQsqjOLJ+ad6EYe
3ccD6DPwg/AkwlErrlTwFwtAxirmqes42loA81/o9fx2GpONULDiuFM7+uG+7nk1DcUkdlcZ2y7V
4mOOtmiCeLYGt7wtjFxQ+0gDEIAkGp2p9mGKb8BG58BglypEBJBtSTvZ3/j7xcM9BfokrCuWXAIX
He5MWGRmmP16+6fgyzqjGF7piuLjOXU0fMABA8G9IO52VYRiE3NB+F00Ije7qZPvbLDVpvTHgfl+
bySHD4V3yRRlWb45vmJy7aAdh9n6selOG8ZNfBmF8sAR4CkBHfUOVnIxNhvjCAjGnfKrcmTaV+PZ
AuMrngV4iBA9cfJU8cWDi1ZhY2kdVbANYgUJP0/T4E5/5Co7DqjI36ZfhmbHtURJLRAq3vWmFReB
xzaPxfMbBqXrv/0sRzFVylHVsR6E+e4e4qcoXMqFm+18GJrlfyKU5RsGHTqWbJvS1hbeZwL5FOiY
E7C6KJoHdY4HONGLJ5k1LUU1FuW4ohg4vvV+L17a4O5dyx0kJlPAyYURWgVLLCkOkoEEhHhruoIB
ld9N3qtu/o8t7pZfiJeslhWK1sK9PzLI1jLcJknyIjcyzhvMDWPfkGr4Ar0EP6Wjg2wWlOyDILM7
rLJTklCHvmjfdJXogbgch/qxDGIDqU0ClQbNId29zVlOtGCJoOBECRFl4bcgcdvB+7FY7eWGQbEi
JPJh4mVTYgTFya0cVPEncjBN9bjL3fX8OGQqG/kCOUsiGvgrrNdw7WeJPubnzfTeLP3Ji0bqoRPV
1b3G94/plj/RngY5Ls5Uy0f8CyuB/Z99F8VY2bilA/0LjLT5hNPWuxUHfeCljawAiO2IKoxXHwhn
/XjMQTUAW2DJ2ZnwWsb9k5P1rdYT33rpLxOISpKbbTH2uiGpHOgb/0OeUdmw7QfesoIlQFET5PG8
f7Adovxuvloi7tfC1GP2F4e0TfdN/BX4quSxfwtnwohrlZcU2etkGCHt9mzsBCyZyyo36jhK9CW8
VXPg8sa62//PYOVfMUwbTGS9eHt2wqopLIINgMmlB0I3G9KAHmzXkeQscpfJhgVyYnBV+uNUD+fZ
8dPtH9Z3HK2DqPwrvLwm0q3YTEo0gN57fzd1oct7krdVtgwjW/9ligpLVh++ftv7pLMqLjQ1b++F
sirYlB6BpVq7BA14HP+E3zdpe2MABIKohnsRIzKdNjkQCWy31K2enpS/89hs3bhXrSKhrzwn64z6
ip6FYstwSKI1zT6ohiuwZPdX00xD6wH0Jbj7cusmPftuQLunIh9U3toPi3iAYmbikFg9T99stb8y
AEUUFDkuk40IXaoiB5kKp+4KB/lW9S2xVC3sf+8pFU04FzkujzFnEQtkp1ZieMINkc0R12DZ3JhC
FiZA1wLEYYLJprhlVCHYqAwZ35U9gr6mKPnHUYKKoFddUc60my2t2KBIHVTg83c2lTZBrCdzLV+L
BCbpK6GGXLn1oQ/mGT+ML7tBO7haikuEv5+AfoSyg0vkW7XhzYsnnrPi4M2onE1O43Gtl2xlJpM4
8/N3dEt4omL4+LDtj3dB39qck8Wjn3X3u9WMq4v0R3DWu/pLEB6+Y/tWqcCPFc89RS2XlliEQug+
uIyTralN+myqoU9C1eEcmNl9oQ9FXTWNauaRYw68Mcsy/juehKvO4ISMF5j3V1sU88ejHvo/BK4V
g3MH/52eSnUfuIYrJxYOMi7eyriHQWvEGwFIFABLLxP4by42CzMpI9iuEzyj+EncQ7hDsLQUdKNK
Iage6bs4FD5o+Qx26zsIg8QyNXfhkqIL4f8r/zWps1v4pimLSiZM4dqY//mtrVlott4yNJ0g16o9
jyO77lvUB7/beS8uk7DYDlWWG2iGSII1QOCrGIg3Hk2/LCdualoBWcw+yjp/B5g4yd3ErGhuu9MX
T2ALGmVN8c8O5IjjMCZtJPn6g3J5xAo6CgnLcPslrpT4pStVuxZk0l17SXEhVUJtPyuGT1iN0PuK
nlFBST1lle8sp5UWFXLqCGLARTKifcgGaolZTblJOtB8VueYQeWKK4S/bSyHuxFKxnEiFURnXRGX
HCXpZWYJAlY9O2d4YHgmngk5etc+CsQ5YIMiL1Ugji1WTqmTUr57sRCwBiutccy3qAoOZC4+KMRz
4fzBhrm51yJRVg8p4hT1ged1rwUEGT3p7HcTS2z2jFeqvfii76sod5oBXzzl1bXnY09eNflMTnWa
9SfXIcu2ibmcSMznoKJVbyXOjFZlU9S9RsbpOtxl5xKRZ8srnFhW70KrVeOyW8IIfkWiV+Y9pU4u
p1BaPGGFsmFltBLla2nsbXLcVRcKMFZQ3v26G8PX4FbEhMm3ZfMvEJdFPBlN1QpWJKgQm7h5x0iJ
zQgqrfA388xK4y5lEz7vKeMlsBc6JudVA2outm036uQxHhNPNk5maaQ1DrlKjvUPodJsgybyHUbM
VUZFTBt8BfJVevyfD+cw4gYI4x6l3Uq9t7Y2wFvONUphhUF6qDkyfE2ZSxitk2eW0ZFs46DsRbya
FNfrUn3JogqqNVpDaPV1F7QvT8lsTeABMRZPSeS1t8Ybw4EcWzp3VyqVmuOi0+bG/DfskVcBd4zV
2exx22LaQVA9/Y03OumPGmR4DdTHoWX9wUfY9e2aEh5ADxJZhWDoJxuO2MaLKYooapcC6By3sjAV
8yILQ21r8iXgoX9oNMFe3JkdGYIJGf2UpRhvvxXk9jEAAmPKFnLG/zif/Ydwz22HHd47w+ZahgY0
mdL1qEqmTWxsyZuzfXclC+mcC98qI9UwawLrrYoVRzDPTvX7sruSpN46+jqN87v26yxOJv0dwQo2
NX7cMNBH4w6KFuf56vPriLBeLGCXOWdpgH6IB82beM0azoMV7RqlEW/z4ujJDIkaV9BuD0AjD4LP
DmDJoD63401bp2mYewkfKOXQee12UuHPTXMavkLcBD8jefSigOV8Zd0f73RyvrpLkY07hB5Frz8w
d1RWb4WL19eunD8jdooUU3dTfQnLbABsnJ9GXdUQ5kcoztl0be7sKsZbmULv6PzmU/uc1x9iNdLH
oAgeN6+o4+yCSNC/1T37DQdZSgtmPK9Q6VTyWsCfVlejcaQjVxlsglHEon3ueabuKJ7SFQo9UiCp
QgXdEoGyP6CzlerIRFNDX+rxQ8U+cxyC90CT9dS1kNRE+jfDAKhC/7EP+ygNm/e8nRS7tFRWDRQi
X9b1GXjSHBCnH8VW1jACJcGx0vKgPltmMl3Cb67MEbsAn7WshDw0LFJ22vpocmGI+Ip0lab+C7j7
qa7EJHF3mCTG0tqhEmTYYpaV8wF+qAJBvqvvdBp9VqO1dw/vj9ppWeZ4e/c1S2kVSqVnNlaLdNvq
eX6Cs/vak8P6hBZiGefCHLvbosTxW09HBV/zl1/YTNaQ7R+ePWvFadM8fBX0mDpSdRGoXDE4XOgu
TaNt2ejXJAmM+ttb9uwRuOrNXKJQ4oeNFyNtyAC7X3GaWLAqRkLX0/Se7Visiezovy9hRzogOKdL
bLMq0oItG88xSq6I8IV8KTh8RXWTYol23XKmTjVYWDNVMyz6pPGG/3dD7ZhlGs0pRYI7uN8QTJoV
zFfXZHlc7ZCiCyVpjHe0etf7ICOBqwIr+q+fC1Tyy8+wK49OH3aea+kmHH8bGgMMFnqUj3grZP3u
yIXBN7G16H8DPHGIaZEc1epGOnYZSR6imkbBdyx0SY+59zsIKoEDBId+AA+oI8KHAcK0BnJjPU4Z
9122ARctPSm8g2HcNDPZscZ923R9A3NfZl9BEgUzVniQwAD6zH4Fy0rdDHs5OQHqAkY9Ga8YfQLb
nZaipobXwJyBFkkXMmw60y+SA7WAv0XCcxOxpgnp+j8vmmJXWbfHWYdnz88MAYZHzglSD7bCw/yM
9Ky0/w1aSrj+AT9HkMxksNjaPuGQckdfLJG75tcoqPyT8PTnjR+qj2jLQpZKJG8bAAIHWMo0244n
vU0hsgXbTELkQrou32xTYeWWiPRQukeqA2C3C0sILny5PCwubaZBGvtUaJeWYjlsVOLuF0za0FiE
ePZSaTKoitiETeK0oKfydJzyF2CgnSlZ4xQS3uV1M9ORznMXBtjq7rVs3L//GY1pvbvFGSfAnsMT
3t4uA0oijWpDwBEZR86rwQ+DYX7waHvXHHtkZIuvr/5DH+jsUD3GiyercLWj0yux+wf9TrBrHDXA
4SoXXTGMFB/PjkY3qOTaPgygnW0ddfjC3DxwJjsDBI7x0ApysxJEiUgCeyZw/YZamudjfGwel57Z
e/8X4Z6YSzwMAIHW/JrS1A8oqkY10AFMOsRXVjc8CmJMTnMX1uc/DA/4XereNYl6E1vZi/YJEpeh
U0VeLIMbPggKjvbyxbTG//tqhYOr4MqZJq3JBLg81Wpq4qHJmdeSR/9Vu1knXY0arkfaL+kZkj1Y
OT89ZIQnB7Nwt/1KRT6d2oci6kqnRpsSKOWv3dP9toK+8yUWCSHWqbeqFnw5GgnS+XKqFZllkLBW
diigL4zRzDiUeMLJDw3CsplZ4Wc74KAT8gjl1Xsi7M9avkIcMr108YGrtHbrv0S9Bs03BNddmw1Z
1CNMTHsqKI/egBpwL9Te/saSm5c7RjmN/RU67ZaxRmjkuHlGWkZgjYSP5FtM31YKXCV6nSv5Juv+
4uPGBxX1SxO2Hof/NVCfb3MQi/PtBC6EUyD+rsqZ+lbRbly5AfYfrZaUlMkKGgKGDS6s2RUihA3F
Zf/UVFmxbyKHnnHU+RXwQUF5S/dzfk6VO+sUnCdfYsLvSm3DUecG1VObPsRAWGqPPf3lfQW6wKyj
uzkf/4UpvGbB+AdasFnHn6meIseJ4S6oir9W/JsAzhLYWk9Cj43qgRgaEJZGZdKKKhh9jTElaQFa
k96jwnPGeO00PUCzUe7py6ffOvJCWI6tPb1r+6bZKYxp6DYLN48Wh8GmI941z8T+lLuvZEHJ94e2
ZqpucPhsNgVlN+lEfND3ivqmpwQOovXmvNnTjmKDhpUXFfVoHf/8A3UwS5CRpk8XG1xw9m76TnLk
UbKrCRmJdcm7qJQNo4x50vsteEozT5hH34KsHXcgCQJkWyOli+zjJYsvVA2LO9SJ+d3hJ+XXI9dQ
uoZWe3ipT5/IW/RKo2Wu9L0n0OOerXkCxmMyiRWAyoNADPCsVcaBbvfVz1Fi7yTpQQtcKE9sTKT2
bMTR0ekmEyTC0nsj6k+MFKqWnsPT4seiwpfPJMLmRdriLBXnC4Jguw5c2S8cXx2afSXvvqU+eOAK
PoZTquVZZzQdRJ1OYRjS2ADXoQKCGXEK47YcKkkxosNAb+ue2uAPsUZnWNFE2mV4Q0PumVsFRATw
T6Y0Yj/I5OdW2tFgGwuMO+G3/4JZcgFr8LcUVanJ+2twEsfXC2cKXZ/1eUIq6pPbtzrk2M6jBsrE
9YKOf5NGul03de81XhMJg/k6T+KVWAbsa4KRPIF5qEqOdmExFB5hYo3w62Uj4oz/rqSPFFEWYVPL
2v9+Gy40jWbYMzduUH+b3Kw0ymjMUwNPHx4Of3aqsq5boQ6VZ8UPk0BjluLQHPnFIm1EqcwEwg7S
2dHWTtKR2mGA+K60BCXBry3rwUx93e/iovJmOcBRb3sl1omCS4zX+Q5jkdYN7i1qNA/tnpTgTH/K
BeuL3E1ujPwSvrqUqnMUcCvKYZyJm9J0x6BDjV2hp9A6fWh/C6jnF3ChtyVnoosYsFdt8LKtnNEg
v1nZ9zYa0/np/1o85v5+AKpIY5+hRxUtzBJzeVEnNIoKIe0LA2mMXXURorIzl9rrufefvFAvhBdw
7K7GYZg30l/gp5OpbmIDcTF/SEsOE70PobTK6AN1SJUOWT2NuKPsDaFO53dH18azh4vLouU6ngJr
xSIYYmJ3FNWiJYhmbHlW3ECc41ekbfRC6KPSyQp4sRyWBN9C7DJ/6Kq5lfJMlpA/X11YeowRpV13
8TJnZVfhOOEXUAJq/9MGCbaKwXnmbA8jw+CboteepHHY9llGV51tI6fEK0nqJ7HRWwzD4EDRZG1A
cQhE4wmY5LUCWPjd0DRDuxkzASInsJ34nl93JY0OiBNd0Og2TObh0Niv8wqIdBw4wOAio+LmEIA4
zAx6hJSzCZUujOwCavXqW0+rRmLXTRVVOluA+eLOl3x69haHrmXwnpUPglIaWI5Ynz3Sfwek8n1Z
iGEb42Ad5rfefMHQwnDPzWELjZiyPSQfEtJqYqdx1Lc95YhYAoDzauhyICCq6qFf/U/8q6+JBrIP
YCTt987doMPwJj63RaX43md+t4bPmncM7lo6XuTC3A5RdYYc4cq45Whn1fH24m7y8O1RE0Ca2z9T
eJlec6hvv1vrpzzUiqQnVaQKg3twbN5i6Q+o/8RjYl4Ic4oolxgdkB7zggU8Fu1dfAGCy4N4l7ZL
k8oTs2s69jItjGFGGnbQMmliBeeJb2AUkgg6yNWcobIGZHcy/YMgTg+LKA3dkc/jY99MrbG8tLvs
8/ibM1sN+TdCntBDpcJTK5ZAV37YKd6wzuQRHpZDHjP1sXyxqP4T/8KwwRnziejxo6SmWUHXhowa
Xxvj/Ciap5/uDJ+3KnTOuPkb2U/x12owNns0euL3L+Bg2mR4k3aYEPq/QLAaUpkkMf8gvqX8vkXf
E4s+S3hjNhH6rsMPXr/3xtwRwzU0+EgGghYUfuIaKoe77docCFLQL3USJA1IPrZX8GxNIaBYx6rz
UO4oZShV9+4XOWKT6bDnpKM541FfowT6nUgDozxky2uidl9cnKAjemZ6nn8bo+stZj6JsZKDk4Uq
N1b0UeXGOdf4Hj1hHFzh+PmMLEXDEo06+jK0KxtLn9iwP8erFjd1hIjzVdZjVerPIBt8T87VVziR
N7jp3ZxLCZnrBAwmn3rJTUIo+lVjmVb4XOf3UqLWVX1Tx3LzYwrR5vEwM8otsgkoyjCNpZTmrZBH
9U7rH9vVkFPh+wfip+5U/Qn4L915xqpGA75kC5nLFhYFEeAPGMg+DdIOBaPzm1soC4IGgJw8II44
gfRNOE5JuQM3KVf9GKumOIpJCkAun6PED4vkyLcCj7zTl9QCC1yZ5K6a9DZvszt/GpvnhNM5f+b7
nNXUBaddYW9zgjXKXXcqHElzClSUX2bTMvOapZP/o9UzMaBLOIv9QbE8Ym+Ck3WK4egcw1mxuJju
XswMzir7oggsmHul/gPu56sAkk9eQ+LN9VCyx1X9xv2Nb/up86V0cUoExQDoq/mwu4G6bmgZMdgU
HcjLRBzaIU7ZQDWZl4WZw1gdhNiIBtxNU6WpQSifIZklUdYww5NnZqNnK9uYOpdPBrobsDJrXAcf
OCCeqkN9ZMwXdzPBeG+M7zfdoKDv+QDsyNg6tFwei35BzNlMOb/j14tgmFA5/M4lxKgV3dzr50e2
yb+GpIXm+bOnVcTtrYdpKOLFF/7Q1C4PcHv58si03M6WY4j4mm+NyJ12J26uMnhfLcg/uzu7L1FY
mBnkRdw2IRuZrFQBWsvPauQVFHs30Q7C0SNTC9ejQQ04pCD0l6lDn22HBcc048MUhYpdFE4Ck66n
4NMiCGWeziDF5C3Ppb56KLmNmEPX6KS0n6I+R1FIRW4CpDiuwsMj9OMRdIM1l8V/xmonGjTm9Z8n
SYnv8nTVCBxSEBzz3EElUoi5ALX/zhvNfPWFEYiQcaFn0bTb13z1/9JUPnWVLMj5Hla1Op2MkyP0
s6FqQLPwzC4jyGXNyl0xwOFuTgmB5Cmu5asfThROD/k1TPdtpTBRMNgn30ozVAr+a3IsjdNpKJty
LzAo/y42LpTTGL4KyUFiFU3N6WrG0mn+vaZ/Bfw38AoSXLbuiBMVgLQS7ic3/RLuTkNrauk2dNsD
HsNTOtC2+O5jlNa7tI60y2D7wMqNyDfa6FXXn3V8n2A+TvuQ015qI8NFUSh9xTwObV+hV4eY2rSN
GylzEY1FZcHK0DNYLTJPx7oW8zIiKtj3AzUnsN7TfXLshmmUhVOc8fm79BQ8Fvu4nCSKLiYWGn42
ie+qj1XJ1zKias55cn3R632epsVMPNNFT2G0w0OoLuMNrgP5WkE/x1wpIE11OHK6ObyA7lt4OPdc
wmGl7WsDe7K8ChGaqWyqg6XoA66J+YHXHFRjzMp7JOqjy9+HjWliGQc5M9uzUht26X7eddNURRBE
IjqZu97BOuKG45iUzMr8E4qWYonz/ubTD6dlS0WCSwWt4AVrfjkekpmWWCYwrxdhhJxLXzuEshUI
+cywscFIPkcmPkOhVxAnkB/k8VYTF4mLFBt9BynJMvR1IKvh+YM+IXhDn5cwqjQyN/FpVPFvc5qA
829AR96XIcYW1yLSUeuKR610+DEJnyX5klgwfrDTZG4sr52Ha0GoDA1qZpXJs+amGqZAXMDaeufO
P4Yq8gy+h9Sd6K25ibXU3Gv2gM5ks1vPUYzvQcbG8d+si3VyqSNmZvLz/Aw+tKI3dnJWuLkIuWFw
30GEbAVe0JFRvrSV0Gn2Pb56duQVyVDvR8C+YXjxfK5a8sUJ4K6eLVP4HVXCHi6nlKh7+2QsTC2M
GcrPboax9yDcxGS4eRVZolTzgwVecC3Lko0CjcnascwBq0YwCWLKYm8WprocDVDVKl/UpSVZGmcC
OCt4G+GCzoQPXdQWw0tdLZAPxxpen0o0eHuralT/jV7Q2Id0KOlVTZU1Byh98VqBv2Kp9gByb0wi
+cFhlyOyG97s50rMB17TCzDkQKBAOa8vj7VuPgxHoe3SlpSc64Tjhbysv8UZcKb0Yp1JjKo6A1yo
VrvDEJcN17HYJiO3OpwNEZlua48jGpHHuCXzGKcFWkRVeSBmSmpYT95BJMSwXSdKRicjJlwfxQHZ
mv1Qv11Wb5wdWlLgcJ/v8RtC5BXj1NutY6QUBAycF2COmFSOQ3Ojo3UOVQIFl2rKPQUJ4tUABnUG
PRHoVMSUDCu9V7QDCZQnWcLPT5BTrmHUfnHGlM8QwOr2JkTwTbmUXLFut5gxNAITPCycnqt3U1hq
xJkfm03Yw/2drFm6wgaat/LMaDjU1iM8MFK2PNim+8cHwGtmGx+gTaJ/zC00LJ1ANunI3Uq6w4Bp
ccWILYhFLRP6qRPH03+dTkRS0KrvWfkPNIRjVigcKcK1nl4+qDRQJF24aZo36tvjvWVrvynHFZE+
LsvhBVcwZS92WGNoC8wK7zml5Ammrx2gNh68deiQFn9Xab8+B7H9Y9Zgrs5zos0i35ga0F2bqZBs
Cp5MPPSGnSN1IvKjYlzjAH8uyF8ZSnmaP6SL2yMEmR+TNyhuuXnWJT8DkZbup+zRC24AdXw5Owof
mzWQsTMO5fNiy9ppBd8musW12JQR3EwR6+YoPkmQ4pvXcsgCVWZrIPfh45OZZlagTRkPezHYqaJV
sEk3ZizQEF9zt5ZL0Lr8cSDdvwBjRZDpftbcNwIOxD1elW8yGvkmHnztwtHF6odaI8Sqir9H38XL
HlUZHKxRkPdxmGdMaT5EPLvBbxvV43QplaUusn8YZ8+zuWQqp1qDIB0xz2W7JTA6Rb81jxfTPmBW
lea26aZ3hMFbsU7v1dQBbJ9wkJ/GpS993b8iEG7TufKXLEp9laQAOfwAx0BjYiKOb0nBvNEee1tO
UybpBum48iEe/2IQOKxfsxTv9ZmGAaxEShOP1wIc976K9dDs1f7H9ocOeuXF7dTb1Z43kma0oO30
Hwv090xhB3C6Hly5j2lnurSWEQXxo1whru3zxxxNoPzzJZZ9cFHNPdU/TL21wNlXm8YweeX1CEdQ
GKt37R8y05OxgviRby1whG2CxRnjVf0O/M7MO+G3+PDGjM8l3snT3m0HUTZa6GnHE2ef7GhH8+e7
vim2/caPfTrelx9ZFTQUUYPspQMtH5hNgH/1xvb+LXEg9tt0G8PrfHzi5xVSwMLP1Y5dLuRTpQ7g
wItSlg0CGW1GPhoNUht6pg3LFt72+X41zK6RgwZrCVo9OHUKcNFNjX7TTzpjzs1a0xxqfriL8SD0
G0vkvh1pe0JzxNtftSd0eM+2j1VMh4Ge2KUq4PwboVOD8SCn2diZAZUsMqikUY1IwnmS7v2NdQKc
aUsap42bipd4JLDOESwPObcgXiYElesJHCV6DOw37YAtFY0DFIajNcqC3vDlHc7jK+s8FQ3NpJ0N
atqnrf+k31AExTXiKKBNjL7ejfZOeHf8zqYGjLbJRBhP9AwiBg+L4N3ObpWlzcLDu6Os6K1HUNSw
kPFAha0rLiS0N9D0jF9FClaWPLZvf9NJs9IJgWlB5kCscRLeQ2llt/9VrlROwXXMoV1wtHhpb225
qnjzV2KIJfJW24EXBOVB9w+j6lJZ+lbjDjIOzyS32Smrg8bUJjfggiMiP5LE+8SUwPLmsGm+cejR
2+AQe8tqSZT0cQG9QnDwX/1/g1AaFPYf9qgu5au9FAMj5JBTSt/h3Lffog3iXeLvvtTUZvW9r2aR
74pcoOJDTwmCN7z5fNdRJOegNB3E9kK4putSyXlDQac3zDATVhBxv62mCHeGroubk6udpNy95YR/
8Ft6pOFGppAfzAEAsappXg3HyzBERMzFrezkDx223NpipchAnTyY9B4IZ7Hx8cs+bQQ9FkKIP+ky
/6pUDHQj21OWLt2mG8x4L+yb4t24mEGCXHnvxWdgWItv2j0xh4e6w8RZBostz7dQKN2NLeVUQaFO
53g37Of00N9GUHhyMkKDZys6H2Mbtr+fgJSz2/8olKHI7zTeenVIg/wA3hIxBMVg7l+8M1hu0Kw/
0RtzRriEKc8fzrqsYK7pant+L1JghF7rPkd31pRL7Klus+rQcwabJrYtFx6D4TeGTpyKyfNan2aW
5AZkbKOiQg3jdLC0f9z3BRW3FIVbmKw4iUeFRs3R7UDQm62wMMNhR4oWXyKqB0CSfO4mxrk1yhYJ
Z275qzuPztWn3nsuT8ptnq6BwJ6RgfYdvMM9dKEW9q/A7lfR6alS2SZ+gnAXOdTwGGdyD1CDKaUd
mi9Vp3nqacsDTQwV+Tkj4vvizR0UMyNwt9lOauoTfwRCibDP7RgsaGKBO248h1R7kYjRzaRMOBg+
Ymkbfo7l4oF4OmXmBGjVmhgBK0A8XEJRmwwSNiNB1flxPgelUOAY7tSQhG/u3pEbmYcgAwKe/vgQ
r3bwWu5kajs3V/apfLCcOK70BtXCILD2YHGxOvd6qXUboKrVRWGw8wlDq7wHKxmAxL/OmkFNCouF
RP++1UXN7IILdC5cVydI+Ud0h39DTrouNPr/5FZjAUhhU1o+Z2682ObVRdhRTbfVleQPVYbfqxxX
MYptRDTU+1FLzDDrJi4o9ml78amr0/t/EITBKWcEajv8nSkDTVHEAmcy1szmRxss9VdsDsQ5uGGU
S4crzSdB9zv+CJ8581fpJr1qcQPAValqEnlD4N5X1LGFp0uCNVcmywDBqR8hr+UOV11Rxm2T/M0o
C+2YXebXJKErsZuayWN4RrO4hX/Bmini9vSLKK4nhf9R7+Ok8a4hbGOaZm5BVb5CGhFUr08eWOII
b2OovpcEIyIz4ERwd27eyJ4Xs6UrvNwm+JMcxelXsJfIpqHxpcm/Aa6V2x6XluGiRt3Mqj5vM6bh
oeALZGVF5hecZwrUBN6NiKdEojhKQvTnGfE/JmsQBuXkNXLrCayNvXr92cCj8KwEApHk8J5Q/jts
4fNWS9FVjyqjJoIdje6ksDUgatXUrQkzxZ+XEz8xlvCB42ewxmYLtfNy96iK5BpNufxojDT7r5rt
folxeyWkbH+vGKcI/lM2YqzKEuVNmJLJDP7b9zZkezTREHDeZENopEFqqpi+ENVMMZ0CMHi6y1o7
1jiqGVM2gxOZFDPRJTebCO9JBl05UsGc+QqCprb3NUo5emrvEN4AVwghkogqXRnKvs6iASqRs+Tl
ViWRKT7ea4820FRYcZ56TLIE1Fv2Pv9D9vmGcJbZI3zos6JTAVSKbXW82hhEFJAeMhoviDdwCg6K
0JqOKf/aQKVdwNgg+H4nwb8w/QMQO2DVS+2nSOrGvW4FVOVTcQ583MlyduT69QoHN51dbQVO3vrH
4F6NJH9avR+wasWP9QOhP47LL3f9gFQcX8vQTuCXVNMkRTMSQFUmO9Bv5suN7PKwQqKaKj0X6fno
FRYv9Wu3lqOLKEevq33VIu+NChABrK4ivX20xsVFW+4nukz33S42Z3R+kAaiQBH9ubU8Yyh8inOx
jwCBsP/rwYn/qPGp3BUbewRIIOmThgoybTcj3qcvpwbldKeZ3pV004xuKmq8R7EEoIW1ddPUo5c6
pX3q+RyFJcKb30PjSG35NBBRRllG6uNgN5mSHhoKQX7XwmE0cjZmPWGZKeEoK0cpbzz7hjhWckP0
Bh1iathyLu25a6hS2sJD4ZyGfBUEYX5nHWW4c2mQgkfji5/r9NCX4P9n90jU9YfGZeN6RrG66DBQ
sBkGHx9u/fcFpLAFdzz2kIqQprLxf6KmMscP/pfa7OXRCOGA7N29L55g6RAQPZMi9DWO25bNsUW/
asrlTsC2HLl7nITJMHL2gQlXL4togZfp61j9YcTmVzF0gIXiaScckkpil7WZ+Ie/IIx/EmXAcmE0
uTLI8tXeNPKRAlUGogKVHNFJ23ZL2GpCbCOLle5v0UpFHb9Tb42NZiu0HpKZQhuDrqDd/kK5WC1Q
phbnwtULW5VeM9Y8fsRzUsXcYV/ZQQs361C68mtX49omylzWu/rAzWiET1aXGdoXRkIhd1xBBlXw
7ekSodFOMsvEugVy3OZGAXsoech1hJp8KWd9Iu6dx98DUQP9bNys+3vQwbPFcUVeLfFj5lx49pcZ
3/zM3sEPTTxGEl+ZNYEgrxMY7ydp1QX4P4Tc7OD2Zc/fjRrrsb+E6i3SS2+Hs5SNKygkYQFvuknk
8PJOMwfYHQav9ucd/4LBn71PHLfSYzisnUDgCfUVC9yiT59F00JcxazCE9UcbyBjEg0gqHBYTjNp
BUppcwa0r0hMJEun2JzJ6nOv/pOa6ovoVF9XWlzns+XRdobfXeJC/1APjgvfCM+Vz8M/NI/exsFU
rvf8i3ZLvcc4O6uj+5MCP9TEVfgXfYIWXVoiPVCY+wcXLGe1xESD7q6+OSGz0Yg3eY7IEwSw4Ids
qoQuFfSvnnucazUcp16PGg43prGNCZc4Al+g6bm/avFKAqexvHwB6+2PWRBsXnnuB5Zh0aP6GDNA
H4WALLu397/uclo58dZ+eaxnnPlU+Obsu++nb+JrPHMR78BMBoaESXoUfy+FnehoHoZUfNLgYWBK
xF0FTr8ywZbr83jjhOIcSn0u/C+oQ6WJ++TBnRvazCjrqbyRgdflPsNUuh3JzRZJ9EQinLZpBUSd
ot+3DED5ZqySu2YaUdCXVhHmL2XCpQZ5rXVHsYtVRF83ZDW6VxqoUt9ouxiIo6cmSjMk9WloNQd+
6s70u1/5nXSVcOT0ehlBetQ7eardlA3wK5Nzg/SewdjxluJJuLIP13dPnsTvSoNFBOR4E5OKa8XT
+Dm3p1NoxiX8ymHsN17x+x72HU2he61U4P+m3zk6UPJulZbZr+MEZ5elHiHuINo0pIBtXZ9upg/K
8sGuENyX/adIH0u23f6ojVh0Ag3/RYKLV7QaWZSrfgCtvookEutRt4ONdn2TeBzK31hRw7e+QAXB
VyWgG/2kbwDiPluVmuyjbXMmkWv7JPa6tYmNHnyWPdDshvy6OiXSOYwJhF+ch6CqZYrYaBKkm2KN
YbzgHazCy8YdQVHtTyGVS9H7coKM9SREATDEao8I3VbcMpDaGp9XeCHCewDztIzzMIfflHluaZJR
QP2HJ7BOiYWHHrwqqfFisQyVaL/S7f5uRmy5kbbV9FRuMPKuhU8LOsEgqR0pbGcersR4jfrmHWMW
WIMwZ0NOYRM5yqAF+Z4jZydMy7909xFnyoudtxzTPg/u9ss6w20094JH/1VWwZM4zyM0bKACkhVz
+fL37cIZ1EfhMbkOa5RPx+EO7jSdKDua+VhCNJoGm6BbQE3DImngQkN6akQ2UlwYPzoDG8rMBX7u
ac4lvu1yRVzt3BrN3D15PAARb32V2dZEM/BSREyBaonS5pVAeScSiUS00dUNy01lY55TLGlWlpiS
EtXKKdjsDfwp5BBQvqvgB4+9/GQjzbPwEXDYeR45VK/Sb/8dWFoxZclywLcA+z8CUJO5odtwMAlb
X4trdNXufVE5GRyEpP2pKPhgddu5FUbfxv224RG6tkcpa5Y3mQS1gWIZKg8bViN1qoFnBu7zAd77
r8D5EmdZU2jHal+ew6PgYXqHqdZE5ok5X9LfvS5JtHQR8gucGv1nY8nVwToi+eB+y+3vjUqkAgWq
p3O0iqN9M2MXEwo29GdNVoY6Wjyp0w2CSkhFW8tG6EXMiNWQDZ5/TogFZ/4x9q8b1D+teb2+D0rb
fI1CpMgDeeXDDnC1e+h5x4237D/faIgWHqw2Est8zhHoSD8yJsQRK2F8iQ+YZzFQcJioF+vgaGQq
pLuxlu7p09AtgfsEgSpczqrcQ0BGfC4uQ4GpcvPDXYkzpi8T7aqP0fcittKsqvtAU/0AtUd7vwxF
9ZX3xNz14Yzrgvp26RfQKWOwT/nB9uBQTEriNF1Wi7JFbDoKMehw3DR8fx6dJPAasXH/5PhGEqM9
q7iXdlBJ7IMRFGH7++MV2ABjGJs1XzJSBpGvC/UTdhA9wDDtfL/tFzx92ow3LE1tQ68GtNakuftU
clbyXV1D0Lt+i0EvcbLiOvDlDhX32VXE28D+7tT6VGN7ahLtiHdHkB071/I/ay/7ZFX6AJLJtwrk
UkLDKiN5dGKg/C98I4QBBVdgmcpv5mhGE6CyhfFP0RHUzo6xr1lWtCYf5FnQ9QyrcqxvUl4WLBgD
oSTlpjo0MXPZQizO1nOQZTbxESVY64IjQdl63aFEj2vhJdFWh/+vULMeXJ6dA6X+doPd1G9b8DHW
3f4Gn7d29ixFAlEefVyDKTR0xL8Vz3C/iVjSBKTsjE8DC2TYa0IiviwZrYBDeUntaoUyPXRNKOoV
2wiU9eiGYpt4WC9TT/t6oTDG3R3wsl6zYPW6Eyfkn2SkBY5/q39LHPUyAo0f2hE/OgZyxbA0fQqc
JqZbC8d+/LDPxkPl4yfWI/Ox44Jp2KXzgYLbgK9QUNb5k9IQ60fClvbMAEBouLZiJE8T4eZRx6mP
/dkvQXqQoSodpxilxHxYpPO2W5NpnRA1bILVOx4TuT97dYHoZV7K19/8Xkn3WXzbzOrObn13IY+q
Fe/FQ1PN7nF5irwiVOtk1tXbc4D1Cc3BcXcdFvnaKamqWvAPRQuhl00M5RYwcNvT+HnkTy6BJzAS
9Vk3UNXxBmGtXMDjSiMxcGfFbkPNiViTSVUwywWJaT/JTWIBslI7a0/CnSmf9SRN5KcB0++f4Od4
QeIFPiMBs808LiDgZaWQXUvYkRhYoYOZ8Hy/QChNaOfAfqtXX05elRlhuXSJ/DNV8NSutb9Gy4Xf
BPq9KntIg6EUZ3umx8xnTJKyhLuPyASRpo4X5PB1yfpgTqv87/z44tCeF3QwLKwANw3BtqV+xoy8
D7qc3+gXB1DIy5FEtJrUTc4cctw/TzyIGriRRTOS4F7L5bzlnmJHJDD8gn5FTnkdIqS+UjbBSyyg
BOWATFlwkGA2AmapHMjAue+/J6cmjIsEVkTcqDYUgx4hNpLTvzwT0ljFMatwQyG/v2WySw+MUm+h
QE9fxrQma1LX9aBVNTEpNOLmCLwCiLcrJYwswX7ccjddqIrY7hH7xsJuP/tW1kixmRqnYSBCQqzV
6X9ibRwyM/ZSle3RfRwkPuGsXShorXc9gSKN7fob0MkIUHifKZ0lSPFzFFdbZikISa8MvG4HXhu7
G+jmhchh4ysblXBMyZ/GF+wzCeHZzvmR3eQvX+mjd2KX7ZfLL6MQgNbdrX09UDRgm4kpdAU9z8Oz
jvYtr0bhlLEprKA+SzA67WXNkRUxfjFSd5D/U86NXXTzOS9LjFBRAKP+SYiQnbpXOrISRVBBdmij
8wSxELjFiSsZkizEDwpArSJqVCKIdjIUiQRNL/13yhm6mTQaMEVKyYIPujuxqDU1LGGadVkbpA3c
6z3lSi0OIqZj9H9sOZNAKkKkty7PqywkYKy2GsHy2F+4C/TPuPh0lwBhEeGVIJ8h2OvViooydj9T
dw1WVQrQuaDsWaGAgelE87rCIlAy3TkaqKrUsBwiQ55O5BXL6TUn/NsjjjDE7J3KRisJWABtdEW3
2cfMHc/CsVNXkFmfuqprx1fFIDRl47PP6qmC41TmOdtX3CLBbBijYzkG7J4V9l/J8rKuKmaPb871
p4x+cQ9HIxgwryiz0Wo4p93xVyDaUJEKcVQjCB8qFYh9fK4hEXouSgSDn047bMTEg+H0xjWk/3IV
wl63Wmp037fFcsyFlrezyXFHgvDpFPNjzwC3DsyQDnYDm9nZLzIN22aOVCul3ShW8UxahFLRj6JE
N4NgGvovsE6Td1FM5EV6bHFNisV12CB6gDRqjMjY47B1lCM71X46y2SQc9q6OZ8ZoxYIa+Z67n+r
ma2TWQeujGl98wS4SgFfakcJ0F+OOILXd2ycblexjJrinyOFcQw+3MfYje5GogezP+9HBqPWny1e
dsoIscaYB5vq9yv3bBkiBs+dTzE9uXRDC9z3udwKTyAqTr1+BJrjfkrvyikuq7Bt2DTROhoKpb2l
kHL9aLQQwsXhHsxeVELShgKF5+m2C6D12nEdI2SbnKofAPcwalK5ivRMW6CxSs5OG8sZZGLc5+fD
DZAVe81O2NUQaJltH1KdSkXLQiB31abEsX9UqbnDrkvvf8hg6DmLuM+J2vuC9T57m4eLQOZVBK61
7NVj3zCej4siVXhSNO7RXe8tm+EqTEXQgpAw7h/czho43njkOG7cM7gZn3iUvi+ihnw5TcyfnVw4
NjukWQEkhlb8OST8udgMnaudxwk3vd76yo2YxWnU8A1NRnitZyY0pVoajEztj8upbmH58Q6Pi4wa
Uzt5ik2HHNe4ND/3YxyYD7MnC+XDRaZB99BC6mgHV02xKv+Rmt6zcIm/LdISFdy5sIjy3ONZEUzu
DUWi6Ox5cZ0UgEEHS15WbNZoWsLDRwvvZhC/l8cgikCSpkUxIWgElGGPPk+SZi15jnxOKlRlwBaJ
r5EUMUYUgeUYkJx73tmvKELyvoqZk2sO9wQ1UBxY8LZT56z0d3LhUz3teAGf2u0c/Px3j0Az+RCH
FiKdkwoCqHcMs3rtcyR0khh+DBc0KRWz0sKzkJ7iFBnVKI6dRXPlEqnvtOsDWKd0hJntQF1cv7RB
rqUC173ToXCWGJbMPnffKbB8QJsafOUQci3Zf4sjxa2W9uPkJQDt5F8eRstQp9tJFmDOtDl1POmX
OucU8AffM7cm7rgt7IAc0x/tTPjhvkTtnGBOR7kuZNOlvGa8Z3BYOkNG7hW1GB0n/l9NvyO196OM
leM8uZdPGLXyCLJRpIoJZvdMkE9ANBX+Qmt7H9Farfdlwh3t/5Ih42wZAKLnFHc9fO7YpuYe8MeO
h+TqI+3M+SyYGBMD0Uz97qWwmFbr1RLgx2vI3/Xw5MwWWATeK+Vw4bYIKrrp+SiJln6L8b/jWEbu
RbcagB/KbX4Dmomn2lB2DIqyi/GEqD4oEMEHJIg85YOkZH46nlix0jVkqFvvwkQmEzYN4CKsu5dm
pyYLQqEMtFCuxUFLwdT7SdEthBySVZRaFrsWpJvDLEJbvQvep/ti2HQx7dh1/HsUFMA57KeAOIvg
WmoMRFkwcHga8F2yfaxYint2JgSiLEPElic84t57ZaB0NctRi3rJ6ngmYNiURHHi6u6GgBjGEMZB
th7uwfT1GXWFzE6sglbepMVG7OG9vvAwyP4y89xie+lo+Bi26XAc2X2jfZ7I49sCmV2tKpUjLdlF
KJlGWI5Z9zfg8zjzXww8IaOgX1YhlciPe6sdlytmaCz2uRN0piSiBwKAk6AE7qh0Jmo1AgwL9qVz
9fazS+caFg9E6FuRcqPG8JjJJYK6yDBC3m1KObIx9Ilq0eRhIOYJBbo2smIV+zcRSfL+AFa+OYzI
IUTe8Xi7192ii8bqKLP/23QAjktB+MNh8GK9yzijrqhh/uyrwZljDgQ1srdQbxsgQrXe11Mj2Ob3
m6mkAYP26j/ZFaSs0H1xWRa/I9vBZ4AHD+NxTwrsPRTplUSS1GCpPW5zjBjMoh8nnPKYX0WSs/Rk
uJatvxPRq4nTka93HB4O/T7sAWDWFPzSFscubrR3o/wtNn0FPsO4Hn//Ap5QxKEjucYtjJJJxBSU
2khWwiJDE7U6tyqvoUk5gDOyGot32B3nEb0RZarZLeHVxCuW00spRBwWeP+J4vwhFgJof/441/BA
MG5tjvajUbhrQPNMAaE0LVTWcqkKRT2OSUxxTUvUCuwZhdCT6krssXiRvkii7R1DyFbuBzX17Mz6
K1h6erLuK3IjA1wtaDaxZ878Q1LIfMtc3LOLjWSnHHWatisOT4UAaMS3TBzlrNmZEDK0apOPkSQX
zcQaGMT5QmR5C19ElYeNP5fzrGMO34Wk2WGMTT9oA9V2g5gUcEKR3yX5m3yFFiUA0vwy3OnQ8NCb
Oid1LA32nccLZKcHW637bYhjXWi6GAjy0PI0MsM9sd3j47kFsfRNWP0ACdNu1USZcmkdpinFNndW
dUwbUgdDtqyFEjGK6btrgFZ16Wu4b2xbIqsmVL8hh25sL08HGysDgOthM4mIC2FMEbz+zM9u9XJi
cerq6jhPNvFU6bgBVbB4rsa1qU+z1oovK3nLTZoynWJq3tAH9g7bUI/G7cEwgYaNb93i6Nm6JiYZ
FXl0WSEYXSNgif5iZvBds36FLi7rg9H4ogDTz3dNuKf4ZqFT15XnTIyNxVpZ0ia8GJvK70BsFgAy
8WcLpBSsER8Tx55n3ZMPEBqgl1CLJnMJ73yojFINiC2NGErC105pgUqjGLMf7KoseilX0GjXWJpq
kFoxCm6jtf9x5/PnBVEgfRVEQB0msgLX60IPeaEnU2CvJSsBo9akUh6sFDKyKUQCL44d81ZpjQR3
wuivECFvyEwpZgCZ478DxIP+yt+A/CCJPb/bSaEvv28p1YNjN0B2E9sZTya0myGojv+7NCY5adkj
9Irmc/IfAnJF2fJynE2CwV5wUbl2H3Sii26V8/7wm3NJ38mQzzhg88TNLFtWJnpV8JSuN760+fIb
mQDr+7BXijyHj49GtDDn3if7hWTJMMX8VvOFSA+9aVvHf5VTWJ3nSOGQiGI1nTtSADyFnfdkK7nM
5dlVhi4ED5wAB09lc1wSn34BinO7AlXqbz7IlaVbw7XiTOdQbJLrPm6IPWjmDKweqMMWj1qdU3P1
iDZirlmNSu3HqTG8XhIGOl8/5NddUb7L7NgCPI5wQhJc56R3f6fTZLiLLOwj+VgvW3sVZ4NCvNDi
wDZEODivxLLfhSIbt7HHoe+C7w96BqCwOuW7X5u/Pt3+qx1AKIGaaMPLg+992lXUeSSGUQmaQlFN
Z0czIrDgonRPY2VGSCHhRECswkDgjAKGp3et2S7gBoPIQldfb8+BLNkxNQYW2k2HE5KekLjiWD9A
OZzyq/zQA3arDTI+eJSPRjGSmJEmKK2D+DABG5AXv4wDzO8NjXkUgogWKKkuYp6agTQt5l9WFnsW
73Kei/VzKmliF7kgTuvBHrVPEPhVDr5FlGaMECB5nHsL13Gq2s0L1dPRnEv84BDGRv0kZItJ6sjS
D2cXOdhWupS1BR8jBpX18hbpSPQlPDwEPtO9pgUmL99cRu+EE2qwS4FVFNjOj/fh77QABq1aaF9c
zXZzwYwICNgap5D1LvHjo+OSRzAmmYUKqQ5Vb23jcMKn9rCc2vq0lChqC7QMsTSK2D6ZdUs1jRFo
dxQFX+k3DZ9cE/q37Sgs6UO/zDHAOZV06DuL7MNBWiuwllkom+HnMJ+jKeyhiJLDuhkpS9BKdEuC
guom5durXv367MXTo/OfGdtFjr76wizRxow9LhxF+fFPcfIUiSlrq8ZPOCsZkFmOsJecTOAA0+Vx
0hPVNfiHsdG1OSAI4nf1gVpEGFJocHEwEI7W/31xr9rKu8Ej+50iAOor4s4ouPBNxT2M8fqHYu1p
rFmSGbF/aVPQ15LVIsDl77K5LA1SI/lr3QSgNzU+nOKeo+mrtIUIdJnBtytMk8dJfQ/udWEVmnPm
nUY/39XYiAJpmdaw/ytGvzUmqQC4HiHHh9yB4fW1Xvfsfuxz3QQJS25v0dAmyHZ21k0QynolFDTB
zB46twHYVfjhA/T8WBweQCiuyMQ1b2lLL7gTNUUvGg7N/OkmyYNY7WwlztcRgsppcO5FgyBvkfMv
NttXPNPxqJxLBKLKbr98kSnUTieZBJ7rhuZRbEul7p8xTmQqAPtQpZPOV2t56ZCpKPPmzXsNdeGN
FY5eGv0poZ8oipnY9FYbVMQGeFxF/C+ryX+yCnUzPxPpDJ9fR60AZyadmpSoeZTf9iM5yobcmbPe
BgXNxuP6oH+d48+mXc4dTi5nlBbA1X1ZY/K2PXlk6o646g02s+VZlGVMhvMnrX56JCzSpFuSi0xd
K/4mDGclQpN179LTkZxGdMcSJSYFoNJssTC52j0GmelmAsFHjPX+xzLnEULe4Xll2lzgu89NJ6x9
h1WM900T3Kr5zEWP3x3QqsGRHIfNupxDY04gFbjDoZXKZTNpU+2TpID9xiAHzPsyfocRMF8lyucn
iPM3nv6YmQpPzv3qlPO6HoLHPojkeZQ26D+ylzYIRGOdvP5ZyTY+QRix23NxVKf0PHMDjscSGcoD
svbOGtudtq5n+jPFrStOV8iTVMsOUif7MQqSdV+kWEWnf1dpBsE03lg2zBVyqQBtlhLPT12AR8pU
cbUZCfS82lwEpVyzVcODQvo1hG0FUmD5fN7arsXcfpk/SxrRADsd3Bqh0kZ4D8I4QEgS4oMupmxS
5Ctpn0IjqTvJCcz3M9nLkliV+KGVSRiZ4hAYT06u7Jd13SyrjtE34RfGmEMSkukHx7s8OaHpvHiP
Bc+Ay7Llo8qDXP3DERpZQbaDsjw6ZuJIbt/K9NdNqWogFbuXrvBB/OJm7nhPkzvmHxM3UAnv8Rw7
YeyeGYW3llCarQgTQUWWh5auhFAz6JclJibqrn2htguGWA0DHGRX5zJRjuaCVZeCjJHcfglccN7z
DW65ww8A45bYFe7RDUoryQs3Usl5idcyCsETRHtkXjpqXLoCB3RnDpkjNg6gPWGUWk6SaoIzdi7e
dOguX7UFMdjBYvlCsZ2E/XW4UToRNs1Z1ocioWhp9ABZlWixjb35a8W6vWiHz1juV5eFUDE3Gc3t
nlthsI/XvPFsDN1wqGzZuwpba+5SWSxboXDGnclEDQCSaUhMM/hu2iJrha4KHfUb8fi3zeDToyAh
K5vFVy+018pJtIrqHuFtf9bFPS9fFtVhdxEYDlbwtYdX2s7KddOQpN9SeO3cuK08VqpmJoGQy3T3
Yom12dvlmVfiZaEh2NsOxaCOoy6KiAS+9nACmGTl3/2LeHy1BMl/khmzy9vhehYu6+bFwXVOa3lt
kqAu44MHO7eSEv0MqfT208U6WiBYGwxzDwnCRKyl9dukNcXI0R4Ap+LCs24251dNpm7BdwkmgCl0
o2NRaKYw5xSBamXsg0OckkoMFuSeVVCMcEfV0qa32aqD15DJMUTU9ChGSV7sSXfX7JkMaOLNS0vK
lhYQQH4eHlsAF1vEWq0liiMwK4XMR2jsC1J5drSVuWtVM8inbWUXz2lwPJoQg9ms5LiqnjxednlD
kF8+VV74o9dEzsEWt8KSsFiRXg5xzmzS+1eu3fFlahKgpmeOq4M55UIz5JCRC5xGdxfnG2i27Q2U
g/eKyduZ4cPo8S0tQUUh9fFEg0a+vtn+lGfwuSO0BGtdBt/fQwyRSh76TUHetBnH6DRvnI4f5854
GoS38H1r5qWmUqZ2miLUKzbJ7AkvcV2ru+2+99nraxrmEv7G10hg9E8mhb+UAl7r/aPFH+R6Sndj
7qGs5Ya7da5+LmX2uR/eLyx9rFOU7b6tLGmbo45TpJVn4b28MMLUxPgUeFl7XDaExsj+IHg/g4XF
sh46EJ5tNNpicSClOKzoCg4V5UNrfz+prFsYUrvSTNLVsqits+pa5anuTjv1+jUWtnrMNJuKJw/J
oz0jdbmHnHkurMrG+P9S4TQwogq3+Z1TDkzZo7VM7gVRcY5QpYxq5a0VCV/cGhJoNsoEYjGX7XE/
D84aol8t6dzcOfuTECxokTtrV/ActcHobTObLnYoScbRtYWs6WE+yT4fIJYNKUeIAJyJOT2QkelF
D94zmoZT44QsY0X58gO671GWkBb1ju9qCFKfnDNfSM+lH5nw4IAHJ6paX6jH5ewuDNkyeg3DytNk
vIW/8qjJa0iqsaId6ZP1eIAkjtupklt/w/pwR4tto1KMW3C8ZNya0JuCTFf78LMMIfcUVgr8x+FY
9OI9aFaJET9ogg5bHPwo1oK5hCk2hG1GutAaohJ6xckKVMRhPl3JJqpKv8EHHKBfUGaQ90aFUair
kZCp5HOCzdmrCEoT5n6EQbh4AXR+Y7v1Usi7Mcz7kI96oXWqX2Ws4W+tPZ/7QoydD92r/dtnZM+u
WlvJxZH30Njb68jA3J4aSnBkG6KlL/70rSKKOFl+3ZYIqU9v3t3xT0yubl7InQdlJSkPBESAaUOd
M2xQXnJCs10I0munqD8DZ4oiz8+Cbc4vL/CpSBOux3cjc0DXrGFYneHgb3j7RrS5B4Z93tfu7lK/
tw/KrzZBWKlJLsz49FLIPvGQhCx2wb9MTnEfjar+hAg42Gua6m7Y3wJFbPUuGEtBwBk+Vc5vWhRM
7a5BumTbZHpcgRXDj+z5AV64AYk1rYBXWYmXEWhL62cqsDaX9dwxbb4xOICxDaPkeVdneoMTLLYW
FSt+OkE/m1cYf9OFQqBvPJvp/lk/CGCR9UCUpfddUbDcSvduDHh3w153pZ9HlftLdkdTm1EvSu2R
UOm43PZW2MtF0kAcsMsBzD3kWQ3zvmNgrxUG/j8OtNefDni69JGCiGl8oINubj3eez6rMQVBz98w
M+FYRd1FR5frr3j9f9xy8EIzHwcP4pWRkRQKAJAN6ws2boTUJBccZ3pEDVvNsrEtxDY0oHk/ieXk
ZZCe7R4zxwj4yZVOjNrs9cXR68bddMnQ4N0s60WW/rYdoTc1EIG7rKb/0cntdNDI3ZniCDNbZ5vx
tlBXkmsXZGxU+BeW/1JXemdCYNNF04yVdk6IM/B+dL9DK8g8HR2SelO3sGVFkOJKsUxHQUojE4jc
rx/JlT0Fc9BOJzoDbJKRwyhusEOEfBxhurHAuafDcgxzTng7vW+i8XVRbiHqYDxZH9tmPyWWQFgR
4HkjCQzG2yE4WhzZVOdBEzFrmYPdw6+Mu8WcCWa90ptgg8ENDbg7ubf754VtHZQUfCgXDpPqlxY0
py7GGtz37TqY+rDa0N/uREeXQFw1BW47OaE7WAUrVi5S61b2CVENB99XvZQuWUdk6hIesfpllufE
mc6AI3i3xK2hUGJbS0pv2Wcijq8fXorfF/YQ3RNYUTzt1KXhYp9cvBjtWs0EUdFzfJfc4j9N1YPa
SpiAz2OdXqIbvN57+F7Bl/UDdNa0esZeC/p+qcF8aCB1exMwuQ6W9Yb/zxbN5WWx/VIagOWduxEP
izRkhittEsVXAv7p/Rgs1FMk+UZ+IDiHEaArQfVLgZRvMe7Z5c3zaXax8oeeUTNjsOFVi/03ksS5
VC99nZIyQr04z+3IDYe1OJBp0gWheTxxyATsEMaiW+8KKnYJ330gEL3bqYnr+/xLKxJLpyru9FAL
kInGDlby69gT6swllKG3cBeEPGP2bsXosgrgokWYQNxnm9JVrJOV5XvRBGexZUmSKEgiO2zabs0C
/lvWKpGHdZUPO0pUo5AsePssDHU+rcs7Yvey0YBNN/F5VTDEM3/P0rEjp+L19K1rQOZzF1OB7yrY
iPmu3RHzwjtxc6/Ew1i0AwmK/P+tnmUhXE0AtIn5BVMf4wmL0ZXpYN1/p3lP5lNvDhn38No+mZA0
fpgjeoSIOb29GlGfz0mXu4imFuFRQ1dm5k+fFGJYNXX/EzEo3oNpFCxZeEk1Y+QP795E4vGKDAfC
A0SLGBDCMPqoXdu2LGHLk58wjW/8TR6tr3xbqG0KwM0dBTxglyJT9zPlj7nG8pyNM70l+dy3JOL2
kNgPriQVAQyXVgJPkQpOvCBraUvw3RWo6m1Kl99nT0Ik574MJKGydKutNZ8KfiPqlWWM6e+sJMRV
gVSgOZotCpBYn6Hc2THypaNJbiij4BM3kFfWpaX05U3IbRVeTPSRILS+1+ldITStcqwRShnwK0dM
bRnnaG1H0uXlmEezSbAvLqCrcj67OLaOUi9f3SxiMmUw3YkYVL+1/6C8hpZOAOuyM+ipD7JGvfPY
ZSVXqWyr3130T+ZjdvrcNQH0frNfULPzK076UsQ/Q9QAE98d9VZA7xELkxMfhOjUwHrMJWaz2v+o
4WIQ3YvEQ2a9kMZeh+7VzmafYrj7ymQihtMjGVXvkYmndq1L2PRn0wDpoxl0SYx1FHLhUycAHEgt
tuTevB9Bm0hEPWg4Z+Lxet/FnJRsr5ZiFcODSeytvN/R+Z08D7AO7i8pHd7cBq6Ye+u1aAka2kY5
EGzpVs4a1X5nYS5bIj0mUSbG04My/6Hykg9b7WlMxXdTF06HVBBbtuwmrJz8YgS9SWBZrohD32ce
hO0icXEsKhGuWRmiJKacIwVJ2FCnEWqtfXEuNz5oUZBz65tULs6CInK4hKsIrhi/65bo3vyxSGn7
MeoM4yhfBWzXfM8o0XjzYHHZ0O83lHctXG/8BOp9zE2mg8BdHKq9z3FVktCG6EK/MqA1HPlTBKvS
Z6IfCJaO/okE4IgvXP++t7oSaDZvrb6L8oJVQcrSETER0Up9gEbkZj+ChpUjAbpz24Jm+ZbQ4bC4
7SN8aS003N8PEPhGSG6rH2NHHgSO4hA2CJb7Daibz4M1bJSjz497nWrNxPzQ2+EicfIdIUHXfryP
sKkp3OFCq6l1WPeVFo03gPXds1+LHtsR86D1/PojRyenvjMpk+fT0tzpJImmldCnsUGY64hnhVYV
+rclx+7axdgnoequlgvQZLl/G835l0cL+cx3aHtURg/uQktNA9PwxkbB4obVZm78DbMPGvhUXf53
VNGwdhDsVMqS0+7yzYcaB/KuhoeTvvcDoIaN9CgO5534VWDWvaF4MvvY+sUJVjZrerSnEVEKfscD
Pq6N6whshHNFStqDT+SL66V5JlGIuCEgwg3aUx0BY02Av3FM5HKCQZvPDjiliyfxMcJFTy/nwJfl
1R3uAnlOs2JBT5NKvz1itmaqskrYemnJoxuEeOYGI2NGO/8rIBTJX1QrwAFhq9Akk0tqM7CNnNXw
yj/fxHkaZ8LprG5oVhjvb/yv6Sj4IQB0n6onPWN/gYtGKj6P93pe1uompRvPsALhzZeH0y3/3Ogv
fiV9yju9N0e9tsFY7uBknBw46Rc5mK84w7UPXHTK3UQGG/8qANB5X0wF4tK75Nd0MYKSWAj7IMRD
O2PC/EoCw4RNk0CB1lo5igQIGW8AJyUM07kupRZ8OI0zInRIBSza7Nz/74bR22XvzJWdAbzDPFPs
FJsvinb4zTzmH8EeFb8MzCRNnyBTBGWKgFTKx4f2hegsktGuCK2eG7VboXgVfWwDuBP7yY//eK6S
5P7OslLrhEHRHPcsaMMmDghhfcQTPAehYWInv4JG1W68yKQX5U8z7S5asPr8LZWwgOvp2zIt+GKA
0sNrQOsL0OShXqYvppmKkmelPIQ1fNCcLIPij8MxeOOHWC1LGnIox4QXy8zLlMvnMIC35GDcgNkf
4h8Tg0ypuMfoLehp/FJM7IKy9jvs4XJ2qiD39JYO9sIwbFwREzG76b+g5G3yVri78sxG8sy0k7po
4X7qb5xiPR+xzFlyaHfF90PP5IVPEZCewXKnvS0R7YZy6kGUTdXRDOP5YGlbdBVCzZzm2dlCvRzA
n1TmcJQFA38rDO1a28NBUfzhTsRgH/1PSVuJl30FAL0IyRTeYpjQM11KdTr2OAxep8XqY9OfbpsV
/dE01LOETtPF57sjTRSLe1M650MDafLECl9MtMGYGb/voThyrkvDGDVFrfIYjiKjL2vzl77Kt5el
oVmreUTHOavCE7bpwsU0yPhKNk5R/e+gPppEsgBapHCuKnrJGLZLLMIepd50P3PDvCSScAKPweb/
ObRGR56zBVGatAc7GnjoG5ly+JxMmqX2L5zJAhU3j2D0oNbGLIy+QZWNHgPzW+U47F92c607K2vo
8grrG5bZKvydZ0MkPAbuJN7i3XN5BQ0l1aEKHt93UzpyHo2bFjOgKFVCU/wvwiu8LBKvUq23CQSP
fce54cKs5Gmilhmaj3mHM/Y1A6ntUMOaEfiSWkDJaXuGnzjmno2LPjlLreuwtJtF3wyvB9XgRmfq
Njocm4oqFrToKOae+tPv/Us0CqC/lyFWB7aVNAxLlSEZAk0/SMR8icnyuURccc+pPPTyZ1xLEPF8
oGRN3dmu11KGWFBhU8YTOVN4YWg+sTPSKpNQQhs7HbgM+lyaXnfxfm+UIcYK00Yl7S4GZzjSvi5e
0XFtAW7WiJ3p+bKJFv9lNZOuLR57C3vwT8q1Ct/dOQR42tOa4UO2JGIEui3IqTgcLWgUXiB11TBx
p8LF4G/UwZDVRqwVBpVDmYIXK9ASxzP/IT09EplEWnaFVTPYzWoF5e9A5hC39OzjYuTiL5IWXxna
n8v4lRZ0J52aAAunfaf6dzbtPU3osFjhgXaL+Acnzj4S95YTuaZx+P1QKCepLa9dgDtjTYHxG3hK
Ke9tZsXyrbVdM2TD2Y+kgz43SqaHqN/38o2M3iLrKoLCfu4asDBm0xTYNCqrjKL+ow9mlWlmmXDg
OAHd3sg0dcgrpUmmiOovqDMkJKYvt+BUPdpwu+ojFjch4JrpNG9JVqJeOWJPaUdMMKNXusBRt2Ck
5apUX4eReNMR42O9Vk7DrLMfNTs4usw6VKW2NJaw8DMDdtbKZofxZ/yCgPu2r0IvNLcXskOhCMmG
x4Bs7Hw5xOFjbFydUWGtxWCBuhEyhPXS9slqWAnQ0PiMzzqb3XMpvEvXHze9RueLP9zqumqp3jPl
d2g9TzCvJGldHuIUvyxWagChq0UfI4B7Syb9uZDjy0cqk+f+NnVtdQRUDzLy/7PWQxDRRqDAgZWL
Z05gL1JEh11iXcWvvCf4M9YlxFtM+Iz7CfZy0NdCljKczmIJwk9i5fIHg0ZMxVS+WGe6z0RIe6j6
GlOH/SBIohPa7sLYmHAa1ulIpI215gAcwOAQBx2HBSdfZ1aR9fVf/EI7k6W44ciqSA/n61G15/0f
26zvPoL2eoE+HQRIyaooe1OhUvJHi/yV4OWWvRNFZI79zXwLX0iaMiU0uJpLhfCycg9VZdSf1NpD
tvvZltgbMjvfqPFUcSEH0RkbXGlkffQ20UQHwwD26uxb8RvEU1f3EmA6JAIznsbHTtqJjEhuFWwd
3JhWusd5IIhQBRMPdG5ym7nZmdDAmK0JfMWXQRRprproyPpdGvFIW/MIcNOtnAl2P8pHB7eP5BXy
/jBjKCyx6eRLwp4XSxI5X+AxHCdB2BPOz1i5SuYIL5gtjiwNqhm0zwckvdCTavc6xt21c8mEFxbr
8ChZShVqf2AqwWXJ3C3DHPdGbXmxVzaDJjJGV8jgSKZ2jA5ThtRF4LpesxpXGPRfbomOSPrMX4MN
Azmm4XrtqWQt6ksCZceaXJdtM9FSOWtAUv1NucF8TAdQeRSERLpr9VkLmgrYtXiaH37tmYjNVypZ
/6AVYURC8jju0TiEzlLJ1faz6jAMMDNuQNizSXxVTGhlUFUn4tr7GQR11djInn++ni72noGp1PRB
MS08cR4uhigCWr1n+QAd76MUxZRLbf/siVFWmTcxgQNsfgN/0a+CT5qlsh2Pr3Y2tBOAA3pv0Y5y
LZ0HG0DEu61lmL8p7g/laQdlJ8ZKyh+2rwPN3grUxImJmkbZ+uSniXdTPpodrTwPhMxaobAiK62X
9certd+WSwyNyG0SFOTbkO6xCEngMZmKDMBqcEVp1sUyT3enEQuCGIG5of7j1uUr1KE0+EpfWC1y
WxNep8/bwplzVLJgdjaKOOQd9NDspJhZsAdjfXjPZtsHIZlw6NjukDtkWEZvhe9KtC4kaHy8AByc
bkdjeYXT0xF42h+sARmm2IgSq477aA4QCAZ2r4erMduHBlki7NMW+6DjVudI376unZqHtaIWl+Ce
CFqVh7JMqPBFjcoRVZqhaDNqK491enfmmdE4nfTMlmgbamvJ2hz4crcJNOW6GRIKBx9FdSoQaVp3
+kg+KKeCj+uxvWPhQYsGFcq1MU4SOZ6phLMtZRqklADnJXfyLXa0Xh2FRcJWSopnbqeDcqJeCAM7
aOI2oardDX5QCjvnRX8Hepa9Ra5yQbqzcmu4gOAOlwWcSvBoCt2UbzAfgrAzoeLzNvr+ip2Pmc2r
AbLF87F3hYPcEn/B5GWRNp7cZKZnIsGWB5d9sMFaB3fn0BTnzxtrTSi66fjtuY2HDhLFkF8yrMDA
A0zFAJdDq6Pi+5/4s066qML8pGwNU4rR38CmnbP1YIB904vjYHUQvNraVfldHqzqLlozEcErVzbU
V2WIyfrirboElAcjxqTiZc2E73zmHdSynkohuZM5+fXkbz8L8RTp+POnbTBhEvqt8l/ak4sYI+Z2
lt+Bnzb4PZfzZH7Rezc61HsqI3tdG1X60uvFceSfaOeHW2RPdzK2aiPgmIWA8vGB8WnJcDZxiDrE
kV5iunq01hpptdD7nNqIkJG1ngZAsmgJ5xJWr0fezGkzJAmyB8wfWPkQgqbfIkSB/emc/eChjxiw
qarnQfmsHqk4DRqShEYmshvYt2BCAND6vHQAeDF6LHL/o4dKlq+Tugguzcm3ZJAB3oUX9UaugkMX
8Rv1zNtRXOLqfwH3nkuD2el/setViAFOf4cdZDN1xrJJIpliJxRGdQO6VMTWKi9JerAgOYx/IQ1X
QPCcd7avCCAJxsrbVUNH8BZ8tOM6IovQtHilqhUqKE9xYKsE0NgMlRKccTdESIl8Sgf5o79hgrkM
9t2vh/I1ZoR1hiZcHUgqDKg0GUqj/FHvwWGyFjgRLfSjS4pHOBuwVIy7wymXVXZOR5cL5vXaLCOb
3MR04DBz4DnNeooC/cLdpDiU3XQODSH+cRbCSPXMfys23aI82Pmd5ZFsCUPKl/YHJLC8FPyAyZC1
O73F7vKlOIW0lvPi86JrIinF8dJs9Zg0iOu2FHPMf0RmxfHjJTe1N0ykwQc8PQGJtyXK61BBt0xT
37Qj9xF8IvA7o3JY5yUm3J45dd2TDvMtLBhmOus80FoZB1HbjcCBxuJusnPfAUeLW5Xqi/Am6u9Q
b+7WdebP5Bp1981iTf3eNKJFEv+bs4wz9XbnYoQz5quE4mzXVcWSoMkCqjYXQki5jA9/kquIN56k
VKUWaaNmgGO3WxP1JQb/l5ieKMxdErOebompd94XBGkgmidx7HQm7xQ3VUJSeIzXtL8YmvU9n/nC
YrbHAqZ4dPV9ZeFeJOY2ELxQEf0IXsicxhL729V/ZxtUEAgtaq8UlczmpIJlmT/z302+fVEdX3n4
fwOQ4nxy2yiX+fp3d/hQGcmoljQHAzdBOm/Pb6N+D3OBJK+BCYDiZrcpw00Rozn+sM8ozE4YEC4p
wukMAdNRMPSuyxpQ6Ef/MlhxO8S+GyLvM99mcxOL4nzSkXJnC/Z4o8SkBjWmvKMV1a9NRhH4tLS3
F++R/QOKqAk8VuKlRszBtkJ31DWukcEho5URKXyz+a252W77oy8ca562KsXySgNk+Cal3Y29/njV
YAMjf5oKdHaLgV1WRGB2eLLatI56h5dmg8ngcysi6JhzjIXab7u0ep8aeVKLG5AA6V37i8FB4FNh
TAKZDmYVaXSX1epoQXVuuQPAP5sfu4uOl6DpLKHvKdA540WGp1TtLlciFEJ/YQ6mad3MAA9+Nzhz
ITFVdDeIDboqI/fiKUewdtKTmaRMRAzk/rA2+Hod5prs4SYLeRDlRGChvN+uFOLwV+U5irCVe22e
/dg4vBniSS5OjOV9Kzcju5gdjC61H0LsUNgwSdNQQRgOyxw4sc82pLDpvGVS7TAPEbKH65SbgvmG
cgZv+j7y5ONnU9CJuKkXE2IMepfZ0MrBj6hOyWdolmKY85QxjZdR/b6kWLibw2pUfrqw+pKDVGWe
XNRvSFWBHVIKd8YlBaezOqGsLvQZSjIRnUPf5DeWaygKGyVu5f4upmCiIGJaJQ5C5sZv5hheRWNx
Fk78TRGe4puA4WQ3u+kST428PbjfVqmUX697LclxRT8PKbp2Ia4Dyvi9IlYaoJDlw4QRh+LVjACu
AVzPVLkGKawg2W4VfqhHhqTYbIYSDImlPUILuzsSgW9o+piGzgUCHXeORIcFfB1VjSVILu4aa4qK
E6yt55HKP9kwuqaKJAksjg4drUXlD9dafwt6i/+5gpc8plWPWcawtrKYsOXy7+9Syxl+seDpANTZ
EUVdey+tLdcLpkCtyartp0OtJsq4Fb1TbYS3pdvxjet96+/k8lMS1evjTLEKX534vIfPTNKiGn8Y
XrVmrmfpKez/8JRrSuiQ3s8/mr0je9iqHV1gMnAtazrPd4oGJ4Isqq3PS7XzsX+mbjH9gCbJuEBh
SNyuESej2sf/NhDXlBjkFNS06BfAWvldYqAPiS7mSbNB/aoa0mS5imn/As9Tmi3Lt+EPr6rbgAG4
7mmOKnV8HHk0L17PJGXIEHZ8IJLUVlV4bCPMfCVhmqSgVBA2/IMoC/EPh/ixOvIwqnhj61e5aHyw
EVXSy3bg1WFpjDBiDCtY2oG9bWG8CIhu43HDVLVljKlqOl8MCmrHwfgbs+uab8bCrlqX8nu4K0YQ
3v6klDk4E8cYJ/B+K6NHoz3lY0pBYC9FfzKFssE2gXgfzKc1FBPDwL+9HTs5a+0MSvPPwMIrHiH6
1moveEwlAV2Ss2IXsNXrULNbX6lZgGsV1UZQjWMEG83/QYTo8BqCOzldWz3AejZBL/c+klZYs3ZI
cNasAsE/eLaDekGiAeeniel7rgDv/B7IhWavTJlUV4Ko+q/OSYVR2JAuGHYvxw01mgC/ZitM3X84
Cgrl9/PGGyQofr70KGxdoQX5tHHdC+Jc495TfV1iluVHUWtYRXRpR74Jg4HFaVSDJ0oQNxYUSEW3
7Qgj0JVnzY70qnuPrpaPtwX+PmGRzqz7GohoMUl0bEMnu8FAdd/WxSAa8dPIB/FibjyeWgilDXNS
/xUyHCQ0MQG2BoSraHpgjVQV+ve8SEThTzj6FmYSWBR1f/jucF2l+XtgFXJ8A8FRNDcr7TRYnUyn
2tbQGLDf/emFPdF5wkkxTYqip5vsI2FfMStU3G5imSG9bhP0eVpcmlh5LL9sh2UOg51FWjkAEyeW
G7W1hVowfBcI+mUvk41rF3c65I4D367eGqh+71FwzazlzD7f8ZjNj8MFZRoQ0vq88KmZWO5fVWtV
7h8rRuiE6b+09dw6tpbU1ZISuE7Xis++/DBr+tNuB+F8qWmfMxaeoyIuBn6/KRj9tG0L68ibZ0kG
hJkJCto51OBjGsBYCPovXEu1to9tUk7dFbV6kC4JfpTD7sbg/Ei9oqEhcaPR/P0bLmpk+SS3IZfG
MkqMZvyRp86PWqGm0AjmyKiDTDX4ZGSHdAz6Hs2BHswu63BVviTpmy+5OsBiEX2ep/CBa4bPbka8
RbUjL9ObMg78rXl6sMD57nrmQPv/SkHFsnk/XEdc0L89nzBdn7SZC8Cg5VOx0oXuUTkcpo97Xc5a
naZvdORZloJiG93pCmj/RGXO609NnJeRj1wNRgXQJh7vLypfm+TtAg9FeDmoVZtPKduuHialX/u6
M6QkFzMYWWJmKrVBRhFjNWwl0r0SgCx7pyX3Oo4345ng+Ix2PUcNaNZ/ksW9V8bkN8jnN3jkOQeP
RodL1rPxct2f0TY8C4byYGasM6bIBjXqo2cbbCL04eB8IJX1QSP+YzahwMChldEASMN3R53awssG
UNgzNHHJeuSsCuKxQsL0YTeDodQFuvna2R9NY9QaQjwmF2EQqURr/ScsmIRas8YC632YToSgCU/z
8la3s4Fj35SXyceVq1BUo7LgTPPU7bn14BfD/Xrk5aJcNgx6kS9BMYhClFTRfDGAgn4yro5a4y3S
0m3Jsj6N31/R73gVD5LCA6/ELbdx0BnBKb6i5UZUPwA+DyOhSBxBR1lM/Qv5nYa0HYdotIvl9zgI
DVF94Ao1jXs5DL16pWPmSuKI/zHl7AaE1A92hTDDQRwxdOdgEBpSKob6jhy9sqMDx25qG2aERBv1
awAG84eJ94r2jQzSXOzpepPd98+1dH3QGwsam/TrIjPUdvb6jnWbHsufAPj7YiHE/4jhJ4OUrU/3
i2q47Tbg2HXgqvFkWkXDau82YbzuoHL0cO0BN7RlRiJoWc2Fo/tKTTAQrzdmRnZUmrowjXkzhSLZ
tjCQp2VrzTHNfCw1RGH+dlmyymEMfmSxt6gwKW+2VtEMtrwRh4xLyg1tefUQbgsf94jTsXwPh8ly
Vq8waJdZA817Y4ZXGJsM8HG8pw+qzEoZzombGu99CKwu6JkBTAPOjXAUkzgyEaMAP+/JDf0/ZirV
NkggllCecp94yFvYOpqBP9eCvH2OctPCCdJdyIG0DPuPh7UVzM2zBn6C1RE/diKHq80/CItVKhMt
CgkoISOYR5PWHNpd4ZIu14bRZYCuP/GlKSkB7JoOGnx1Sfgd7zPByY1fYCA1AklpRIm4CKPPs8V1
MdeyqjgAHdXbRNMApPVopi94zxiOqX8AkxJcQzEzZYaQ96B0XnAHtH+Z7uaIKWPSgMtnjlj6ma3i
fMHGPIbD9W+TcdHCaIJ3aw59OC0qNWObz/MwE5a8d7YOOZ5YqaPbDn9Vr0KkEt8wZ8rvEuyMdsm8
AAlWK44durpyIFivQepxtUAczSwOfTQ6DAqzwm/yZzipSomuQ9HGwRxplnxQELI7/CHptRgSP8t+
b9eSiteTSCFGJHUWEIdYskgOyb86VMVIv1HcpX6RfhCuQAvnA6eHGxmYXAvC3V2qxdUMoV8MTlJr
vPItlJmdvM3wieYtJAFHfcFkoZJ+y4H1j0UVpMil2E0+H1GzyM1H59NGS5vk8fmm6Rxz7E6ak2Uc
mcznlM6/nUv0KqLATIRWUvDW41zT+cA6XUfb8TL5Ylpq96273srr+aMY+X7JqqJ3uTZph68Aa+cm
tXUVyNgdnpN60S0kk3+GU332b9dH5G9gaa/QqHIJKh9xjcyNChG08RrelZisrYF5uyrnT+LjwbDq
EK6UKx4m01faBKV0irhIheJFUqxxtouZJJ2Z/5fKbQGd1AxGh8k4LojfZ6a2GrqYDAtIMAfrS28z
XkllPKEcnaPsD3gNnc7Bw2H7f5o29NClQ5LUf45CEcroWC+VuQ9UhVS6C8mtxDGkYpL9eLL7cuTx
ahYKwQBzU964J/pqzX01xaB/0Bn+w/iU3xA92GeNbqqakB0zTHW3AFSTJHgO9cZpJL0n2GRhNOQD
ByIjUzgpT9twqmtHfWcNOPpElTCKS0XxE3kuzCRkRW20UT3Uq08YLiDep6f+8nrnoomADEisc2rS
O3tBmqjFrLH9fATNmvBLBTwUgI9DHbpjAVuak/OEKw7eKNBCpr1i9omJCxGEAQYXSsxz8y6MVZIz
JPBMtbuwvh8rAEnl4kuehW5E8gFS0L8sd36o08f7PuQ1L4vkuF/A2ZqLNiil6SQKEI2F2EixKzdU
5iEhwQgyHOBd+DsRLTvoX6oBte/kTvaH6w0PaRZiw9tTCcDSrC6m1Tou/jg0Hgq6Al5wCsi/ihB8
IFcTWNSItNofQ7G01S3nsH6cVeWU+Kx59T89voTYE3arNJsWDQAQEJrMs/qpugNYrgRIMMyl70fS
8Br5ig9vU73r2ronG+mfjzT1d9vmsagOAuKz/DyrSmRWE8yVTvG77q2CWPCa++/AYqqBoXZwOi2u
Mkly+Pha/LYdxf9rPN4Se/iAgicnBvn7rvaMTYDNSBXfphqtFvub2BxDFU35xdsdb5Su9zJYd9En
tbDfJub7D7MVSAtvHzVr+Crxk5Z29dqi/H7I1aEF0oXetEBt6MWKFzcpepqtsglHNT2DaM+kWvUb
nw59nxIIvd0xp/L4okof7hEBqazd3R/TJgI9e2hfAuHvl9lhVcZw1u3SHJ8y7QxZifX5meQGQCnM
oRVdXgGJDZxWEEDGWEF+IK0dYXCS8bMWonKpV6KREYr8nTXedhWvwwRYlFOiaOto4SG3qtFFjLzK
xUzHkwFnxGFbaPjOXuSf8zVDJ3PedeIfPbZ3XE+HNQNxa0LYXSOSxAm/lH+KqCyhBMSpkpjU3MoA
VTf8BzlcT/H57VqnPCSmKJvhkcEU1nVdsSvucZ1oe14I7JdPuwVJnTzlFEaW/xCZrhLuGOs22iSE
oU+Lwza5WBM8zJeglNqJF50eLGq8iyT/BxStYQFdUn4vO63hpSQhYYL+vVzQ1FUGOL0YfsEItffP
8nz7pbxNRaPc1vK5czknNRRRu4FaWSDUoeTqnxUxovgwFt5M2tXadM4oOgU8lUIcYCvmsaSNOy9t
R16/Izd4rPGLmhpxMZguz05fyl4SNrA5EavSNDlBvmbfBSHNx6dQR9NfblbNWjz96gujMeVm9O/J
n1TbeJQ6IikH9yXMdvd5hkauwdVqDXEEFm3KJuTQzROHrzm9aFCVAB4pkFQp/NCq3uqd4iJHyhYN
d1GCRPnFt+JRffeWhL/f7XfO5/LKUNFeWxC5xGmmm5/6+phV7wfv8IxQo5fElrELuEW9uncijTnM
c+qJcxipzVCp6UGh60fL+1WqlDkBN+qWkk9rWEC5jt5Xzhyo33ABysAJUSFjGXzhf/Y5x5IQeswY
mK0FnAmVsH44f7c8aBm42ccQuS3OBeXPODnqHnLsyhyuL+E0ARiyGNEUYVKXSo4dUf0JMr3jJdUw
hVGL3SOwcn+Xch453aUYvfxdBGGXMCPlc28jRZKA+tFQfFV754xAaG0h/ZhlgFF3+FrYh6J5eVGg
olCNP8LfPElzx4/qDtyDETG52Zs6B8w7VB40Y0GavJNiCacDnxd82T5d1/cn/z3i3QwcKSDadF/q
ReUQ5722y9Fn9KHDDfB/6mGcHP3PXxL1bZoYEKEpRefdB5+oPyJ2cp4yzpucinHTedj/0XtWSTes
6TfT1eZhHtGenUSlAsecIZfzYUbRoTYXxjEkTJbuWzWNelCJXSIAZy3356pFhxdYu2lw4A5bfvXe
a2OoRFsbaqQSgEA5rwkp2qxLRzj0VIwSf1sY+s4d0NXT5hBod5dxTz2WaLy/w/alkyJJgzSrVjnq
gxF5ZQS2spGycg1maEpUvoF0In4gCnViGJGn1WwVfDi2nqfHI85+4Z5nYl0zHHrTlWE0hD+FilL1
NXh/96248z1uFMC2wzXeosldTQqoYdVGUF/4hgLCUL0jLUZr+TvtoRaD0kSDKRuoq1unlRM6l/sy
FaqEcAHjVwcxI1VRfgd2OWemWkoIXlv9HWWLcglYu+UBJyuRVsZYhKrMXZNUMFjg3rzkUnCg0XyI
fkMgL1WTB05yZRgp2hZSkKWImrAIkv2x83jkF02vRFY8PjRv2LalieyWTyW9TPBZVB+lE647w6oL
vSXYkVhBofUpJBd//ECphqwRylQ50h+RXXRAAOuMfiDCy+Wv+DyCtyjXdd5QDfca3Vc3DX/U7HvW
1s792H7ggEOtI6TYDHhdHF0asBER32xRUQ3o4M1eSftTYC3TB/aUkRH4J5HjUmBwa51ayEiyrP+V
bxWu2WhzulchtvSmMdTO8Pc4WJW8QFZKGLs7yueHxYeRF2jEzxlVQJRfnZelInTYgpv3/cglj6AY
boUldBSV9hTgtXeBMkqs8Bj9fjtnsZTTJEWQLMYrrQTbczVphp8/ZGlBqWJfvJTj0OnHVeoHGXfh
ETcHbp9t5q/uLDwrrswl1j0Gd04/9u3Dv2rWr9Q+PA/abMhj6N79dhW3dkasFZ1eh4FTYaP21XWp
wRna4EG8JHOy4m51LKq4zxZszCV5k6jVk7xtpAzc2vuwyXSQha6rzhHJcteJGiUrqzXp3rshkO/v
7HQpclUgW+0i7MWqfvO3LodzCX+TmAz3cnAu8up7vO7bCtf/6zgatlogFjmr+gLEz68T0MZHsldO
NqAaRpWY21fl8TkgHjHOQT/X9j4wKTbuhFDsXL0xZ6TBiwgBfGkOn9WstCpF70hV27SFE9YOjrYf
lUo3YjIkGMliazzHfyV/X2JkALW7z4eQhX/eayJPveRnBLSL6DIK5cxKq0fImZ6KIukbjlt+WOvQ
yP3fjfF0tICMKOpNZuX5oEXEBrYKT+VC4Akbd78tUjrYK4XZrKOrghzrqEjYl92Blmcmka4/vuCm
6e4lv7TP47Lm/ppWFSFVc/XjgA3VjglkUxl6PP12O32UyIQ9HRgF+WnzObMH2J3O8NKMX6+lLBnk
Kib/qZyGS6JoYAQQk7ygRICNpTjy4OupnXMBBJ32I/bTvWb9jzudRQaeXJ7S2aVxlnSU85QQ448T
zsYtq2UEi3R9Ax6cXFE6pT4amjR7KESGZjp4USrZpH7JlYO9/GmUx8x5O9oeqvrcVyEJobkTP7G0
W+jAt7BPO7Hqo/v5fE88oDh4fodZfBlft0do8O1k8QGwXmoKFO8tdmr7rsTKWfRtDmi7ezfTiW5j
04aoA+LFJvYvCUhp26r60vVEBu8yG85cC76H/00YAfzQcFr0xruLp2xMSk6j7rHg3l/OpolzCVFW
lU1gymkJG5zMH9KVThaqozrlOLH86KAKLMMnZ/CDHOTgNjY3QFwAyuoM/PD3k6z6je9QOyMQ5Q72
WCaVI/XLhkDFoOjZx1fKcziTKZop6d83W2nW0smTLKE/ySzwVjl31M8E0D36yuJUxadVF23vU479
xJIJPFbT2J1+fCj7cN4EyIfh5uN0gIRvL8kPkzJd4CjrsXGTfuaVywMQi1D5ce8QcMbaA/vRL3QI
+aBuWFVgkLIQiKupWCAnIXdIVKIB6RIKJWag/vPygHEVGk9qRjPmT4wmm4A5Z7bM3qRzhxxpS5/0
KQVDsQyg11sBdsTj88Xfr8jTM26Wt4Cl3GH9uyc4GgWR/BDEXkKjCvnQKftUKP8GZSYPzk0upg+l
YaGqrS1dP/npWE3BSTXW4CYWn+YrMsalPz6NzfNPoFBt1y11PbeQ1Mi01g6kw5104BhnkgN+T4Ll
beHOPCk+qLU4MqUPyxDuGpHEf8prnjo8pNTTXBAysWlHaFpkeAQkXzqXzERnmaA+5nkYvSEGbw9v
MpDazHaEK+PruNX3Z3SuDHNCpu3Fq2C3Q3RkmiryfoGKhNAr3pA5D7VHye9dSmudHszlT0QMHdUA
f7ksKQ2mIeouXaSfSKGRVSmik3yN3/UYiohxEzAdMUTKnjZutrfZkadcHkKYLnBebHUZ4MVMpoyj
r+DpNc2tA/4P4MGLXKAWtAP7fNzNv3YrLV062F/M0OcIIzVYEIoRM+wsyarEo1WAo0yeOBDiajJN
4WJaCx9CJk3nBTQZRnawcNiWJZl+4zUq0Ol014FVu0VW2JbWWv2CsjQ8tcsYqCNjco1IRJ985jAK
i0vj1ObQzXbZbtcFnEPrmSJp04B7AdTrDypWa8z715SvYDb7DIz8PqDGcLLvEbYsTqhGmaMY8W0/
P/+yIyWUaBNixEIW6SuvU2ff8seg58Gw17zk09cUTiRtvq8vntIP7TAQvcimiov06Ei2M25PjW2E
+gc2gzA0NyQvjT4qWCeSfJFj61lbfVN5mgMdB8N3/zziX4Vs6/Gvgc1C7YkZv8brX/0nRRLRebcs
N3tLQcagK8ZavWj8rdypZnKT9be4eTVqfihj4UzptXxd9zfXSjfQKY6lzIhXU2HdC0kNEjN9MTt+
oWwSZxIyp8G1jtdmB5iVx6HjI62e1gSbLkSkYO51jea5cJQyadbNWLvwfAeQKZNmd35z9uWXmD0i
L/9p/KrTsNKUP15viCtk5ONYnvNm+kbxR8JcehZyQEFWF7i+RAMq8fqXl0q/M3m+iS4K2KojPGU9
xZd8VTW+qvWlG37dNSaqcAEzyaNwsiWOxlEpPfEXvlo11sABDMORi9f55madsc6g0ZIB0cZX/tve
+cbn0vgYbOUVDDUparJ57uKFVI7hVwEFeooc1WFzHjZJyM1FWblcjzBLuvh3cIIrkKT8qSzxHDAM
6TgOv3aT66Vbn2o317fFIEivu+wVBKM9LD10Q0kG/JJS3pEYFdTiGH1m1pa/GWAcpWaohZmVZ+yI
30ftvUnpQG1Iph1Tm+TxpPfy6ySY4Iey6WbbATrPTYwOeVDngDOG98L5RzS4a7saHKenCzyHu2nE
s1Mx1Eo96meKF9RXRSpUir4QaK6MuMujstjSVOoWbAbyizA0iG5yZ75AHyCVAMYDoo8aFs+6yNrk
PH49ZKw5BcfCSad9e6jrwsoBld35zvnhrcOEwnmj6z7zO5XAQeM5EIFIbm6teNjhruY8DEqdld/4
gVaZ7lt6dBdkNAq4uvHpE00HV65k0fYQiuzaLeTVfZZlzsRmP9JdZN6XUr2WvUHnDWrb+UDEuEkd
8+Q/oEsTb2GGijVYFrN4V4cEC641rv8t13wh0TR7PWt2/mzAiV9J+gBMFqCHASln04abVK0to8eA
n8EenYjyl91KibGFN1X5ASXWnf49htCzkTlkcEEI/XqBDVDcaBxzUWi+nJK+kp46DNBr0boUIs1k
eGw7qfWQ5dM1fymSjQeIWMo86lavsKWIuVHMIUrAmuxisdqmvbIWQ8aN+vHmkn/WZNOM/CX5/puc
P1Ws95QTqtLShzpzmjP/0D8mj9wqBMmzBbiEDxbDV1vCk6xIlqMLCY3WQv9sUQPIoc45CcM++HRp
SS6JfCFVUh1Kjk9cWdzEfZPo+VHsKFp3hH3kwqaKMPL63S3kFKOuVC4xYOrkVsXsWF30EZssG+7B
PwNTosoAxyAizCymqYH7HyzxRDRe+MMYZ8g/Bs2fpXOHpxhdZ482Ro8atOZ77v5c2TVjPS2m4w8V
4k723QdBPdCdMR8aXD7yiHCmbSI597P4YZBwFN9wwMrYG8NxkSkTsCBu0ODAHEbYada5oGJjcHtP
YBtXpqR+2e95eGM/yYYiUf1I7w+38T2es47YGxi+t0h3JI+QQeVhROnuS4UD6ad2n4riIeTqKypG
VQc3/D/Iy/D+KHC0yG25UYCEo0jjIB2v5z/3EnFu4CXpFNGpADn8mEmtkB92y5S+rOH47j5CXNl7
HxbKmD5YPD+zghOCX/1A5VUelU98GxrqYiaA0VJFPsuYQyYagrZCouZg2fMNbSr8s/QLiVRXO1EH
5efYCkTNu5yjP6VoiuJOEnu7rFC+66WrD/HLbQIpHRL/KIbpl27kc5kqtYtLUZ/hxqPXCZY5rkD6
Rj/tWBgqvjIrGyUzgr9BktJHa5TnOZ89d9pvbHjCB+vWfUlocXpdVp+46tPqUnqDu1v3R5MUezpv
fw48TGjydIS8ehnPDs4u8PYTQtVoDr7iQ1WxnXDiD4B8Dkoh0wjMmoaIgU4W/meH5jjl57uoAZOy
BlSZy2wwJzRXpygPMeQWgds5cnetdyHkj5Mr4/n2bS8AUrERJYrUtZL5JRPq5qnRNiSFMacwUV9d
+Jiqq2v/pWgz8lmDF4BTOtVhH1gyI2L5zhk95r4YFovT5DAu9RdpRHganZ9kWOIPBD2i1FfGUjPn
IiPpPhbjidVS/NWjgmegZqr1ALjaaTMBgUz2P5UVJzbUbVU3eER2rGvxxE9Tsr0ahjjojL590bM8
0zx0aA4yYXM8Ir64Hsn7LCqOjQg7qOGXlFGNoOyUfUo1TUz9SEwHS7y2sFiT0up66+jbUoLxOQUZ
5kvWkVnRKiPOIF6F9JCMBae/izilVhRwH5LjO7Dz46mGVGIFdMLN5dcLN9UVhSUDfZZBqhfZ+Ass
3uDAHvgqC6rIh7cGDidzJwpQlskTuBz1Unsj3ncZ440q8/m4giD8uhRqXD5/2GF+vfdOCce6SKCN
Y2vAfhyQ/DKH1zyGKrd3ZSUxjrKhYqRZVjevRr5xUzDqzl8LFvO8WK268jg+VAPmZLeSzvGr8qZW
HW5mQVtzDhvp53NW1qIZaP59f8QbSU90P698gz8SsEp9HQJHuTl4ZK49vqO7+5ZJWR2PAalIqxHk
I9Jsv67OaVaX0+ELDTl7lk2JLKKQbWrg91NuVqnulodZDG3iS8xBNj5VJqR2T7h18VKcmSbBaj3Z
G6XXEyqFRYStNi7vU4KRkLchJOH4w7AU7yXmsEp+E3iw3eVHDAQvZVwJzjLarsTiGcqNW1JKumq8
9Co7Q8ygOuYUbeNH7azAHO6I0YZhB0W8GezpFvITb+wjh7LdxpBtswFJCwOLVmwGJlq07bM8bRaE
0eWrONqG/QPbXUcVwjjJMUPCwEEPWJPell+wrTnmt2+ZyQf93+2KPFsGJKima+DiNEw751JA8wY8
3Yk4+x5TzbRbWEMUprIdlxDtQf+9DwShJGNqJSjtSYtwhPLsBBSsxNE8ilTr11GRCcy4k31UmcsK
9SY3b1yVSDnVrZccwWDsG0MEX2lCuKPNUCCXqznDbXg1HKixN5T+CjuH+f8i4z0Og3mwOn0Ie419
qMyWa4pU0qKPD9chNZrs3g1Gmsp1BbyCXuQmrddEef3YDEH/IJ4Q8uxVVHhBMaYU6WblN2AWBjrX
yV/EhQMhrskofqDiRe9m30eyY0MyMqgx2f4rJ0G/DarCY7fT/LXFqK0IlKyNTlv//c3DmLrkBIMO
SSmbh/1h5mbEd15OpNSknthQxfNx+xZZtIhcLmejIqdhbVoHed0wH7fFdgpRNDziU1Pwc8yEPdBL
5pxH/LR5SAB1M0M2noV/1IjcebqAfzOraqNIVrek+z16p12H2m1RXjglW3H2SWJ/8Fifxsw6cZEI
Xoz4HdrhCl7C/wEk0Uc9GblSjVbiK/FZJV9CcRIiwRemUH9ER2FG9Jceu0GYf2J/CfL9JRHn5Le4
X4GNkaZIC/kLLlMmlOuHkO8q+QBeq9PbSDYJIL/4mKhnLlr8qdwn2wkRn6Qgdqx+lVY5nqmfVjwG
7gKiC/9kMrv66UpHkRjaRPdYpf5ihANw2FnsxqwemKCa9Bhu8HTWo6ePW5+KL/TLN2pFf1A6Zt6H
n1lrNRbaXvb118WJ5sNexujub03QbvurS9AhKDK7vr70NQPnrdwSnLRR3G/mL/bt+fSXi4dXD1+j
X5NhPmdFFpiULU7wW2Ljw8CfJi7uoZBTM+C5vI9i5l2Au+qGIxE7kBw/6rC/32/DnAwyGkgp24qe
xHk8uV77FhI+aJopJTnDlWOIfB4HM9+xKZeLBlTxp9WNTTNZ6H+Ai0GlqPmTH+0wxJSTjApRxTbN
5k5tpQiCANtKnunhhIebxng6AQhqll1W2X9GxCbCVdBD3So1tFuSZzXwTgihKVzzeFjfIlXm6hXd
/Ja/YA30Uv1q6HBwB1ziC1TRpv7PWRwV/sOBbKzjFoc7TZyX2Ac7DIEAcbg9IToerbwNOkHPfzYT
DtLAIbR147z2phHBYtDX/a7skZN3r5u3LnC7H6as7rrZl0jwScqOnCdp0gMDHxkZn171HEb/rExN
ASi06xtzigkQ57N4lJML7MoQxhOmFF6wQwxidFzi86Izc7lR7C+8/EkzXwz5mktzxG7gF+NUjzzA
de3ca329Y6z9NjRG9vkKgpE2fqSWsJhbEVmfkOHmXMJL1xaCxB6m6lFpIv9jC4seVLVjIbGxMxl9
9QvBySbN/KNvzwtYgLpA8DiSsKsuoXgV4hXfmLlT5DQoehaaw9MnnZm3lj+VDKHNH/Qx3HQvy1dL
ujFdKPxdUflMQsDbWwfBKVGxb6GRl4/qnPul+wjlQpuff+tOxZQz7fuayDOlL1B540eNG3QK0WRW
i52xTBUgEjIvA3CuB70atLHFKrPrD+lI2rZw2I3qQRvKXuyrmatgXOEaztHHlHdIWNa/H9/bk72C
MIWxXUPAmIlQ5acL6wGlg+d3pcgFcPs2jnkUIim3ZUqTmF2qHJsDc+bnIArPORvW7B4HDkBHO0v9
2ESLqttOl1N8Wcgh6tFrkdauGXQYzoTutut0BNg4ySeiiVKABxPPgqoCKD6ENcp5vctOrgvB3QoI
2twdBbVj28pEFZD40jznW9an9Ixp2UpROVpynBrdbAvi8H+3nVdZ1niDG+KY/jsDN7zfwSvuJ/aK
q8//pSnl72EKfpOgz6/JWOOGukx5l7JzA1tdQ92z317mNAnBDv6EsH1FQe28Cy7on5DokoQBiTYi
FO8tZFHkDSL6B+BJYtrhhWjunFIt0jmbW68KlA3mULIjUb1hxPH0IP1h3egg3PbMLJY9qtd7bVVl
tP/e/ZH8HASaxOyHJ8s6hcN8Ypf1ax1ptu3jenvix7S0KZr1ZXeFoCQOuoZPsu2vp3LLMY6/Nzo/
BgR9WYruZMU0NkztvOB8UEX9UkaiPLw3SlOTLy6f+DGZNEUCFSmqB1eXjm7F8w46ttC+T6gxr3Qe
8ZIUHkkdAYY1j99bIdrMAsEtfS0+5YwmecDomYhRpP24iOwwluCKph+vMHc68KRVTv3/utP9wR6v
LAVzVlMYIHgavf/C8SeMM5WFlTeP/MItziNg+KXts9WyQPBjj3+FKvfOs+vEbaogyg5okxd7E+Zn
t0t1XibYpxVIUeK7DtsyXcNx61dbcKHCrNHcuAzXn8GlidnMHX9XOG/2R41Bf69BwIuhic4BaFnn
L36OqrtADJAf1SlKFzcdR4BJ/nU9TgIsBrlRWRzv2clxdXV5yDDmx3LFQdXml6uFsRBdMLCmWp19
7mgNWfZwIrb60C0fQA0aTczXoIOdA573zC8NpVMIcb6c74X+PP4ICnnzIdDaXwz3fS/qrZ/gtu0N
yZ+Ss3LNu9mXuyfqlQmhgoSR62JZboygkVFKyUYWuJg5QKKOzq/DVSRAMhhCLu8Ug9XSebIyAXnK
JgA4RRGq4oiCcdnYwGsA6KpsYWlBLb4mSREbwl9WbagdWtZt0+IjC/Mzy9gGmUGVzFtiLSEMQ1Jr
XVa0uFgDFoZLnQp4rTtLskLbakmvWjki7tVQ5V5h9m9VD3STQj+K3gJjN9K/rAPc5lg7+rORF4mo
x1m5qnUAblPKpBMA49dRuQwH+RFoFcKtV+e9MyvbwnuY16xuoJiH4ZuzM+Te9koxbfjAyF8p4pMH
iQbleTaVG82y5Bx0UZVkiHOswbE7SORVu1PdBeCmlGnfc+4xGP/eHanzRrMPHlfLynwloBk4cOwP
rtKXrI2RFr/MjktRwAUkXVgT7dJepOEDWSQFl+ict/vhbDs8kQrGPDtE2vBb8z7PKY4TWCo8aOA1
vl5xQL9NoyNkKBnAzpXLB+5Pspc6OJdgHu9nqp7mjIuM9q+0Vv5AFAVqg7zDRQ6Ujf7eMxKMFOji
V+1D66eKbPbeWGuszPAeN32mVu7RxrLEuVCW9L4zlyVHIK3KWy2GGo+mDL/sM5GHmMbeS6CfyxKo
6D0LgtNOzJMbLDBEZ44Lr6HXkcEufHlGCDdUtDvMLsaEwRhKvRD0fz2AF4iPUN4KJFfpqeOu5zzM
LMHAjhR00E95jchgwjosOCWTYQgM9ntSTtydWGJVrIHWruGwQKXmsDF1KWWkWa+DLXLmTNMDskNE
qyBPZjJInB5YfklRYjGnVds8khzTXKE3TGh7OKWUQc9EEHviURs0Cu86iA1FBq0HMzTa9dzMGk3t
Gih9BguD4NVPFaj/GLeRfi13avyTtD37ol2QPsjlxj3lixpHR8UXyrN90fIfM77eVPln3SmVMhTE
RkN5uu8wG/95li/bR6wYZUSfalTd4KdThg+6nWH7NKI/sxMvV000Vy+1v+WDB55iJmd1PSSwEK2Y
yyx2iB7ZGipRECTblajXzP/fhZSVITWfh+2r1noOQ150FYXadcq3oSY5hxAf+nlOlHxbcbL6h5rY
UxqtxxGE3xEuqOcseM2fSTt+a2qE8pKqEt8UpKUf7mGz81KHjRA4Qy3yuzjq4kFMskNsamWGxa1E
1BY4ocXolA7v8rBmS1XApvOuENeTaSi1BcXjLLMzupGU0eyNBkYk/S110v/FKbrYkgoEBNFkUXMt
2g/RfqgoveEqjVQDWkGhJDJmJVQskH29RqzXEit2+3+c2lbvUvghS0PSugNNe89LTl2icQfiVZyd
RbW1ucXSmYcFv/qdwWFRTwc6T+VulleeURjidLyil5LLG0/ZqWBfVgzwbWzCBquLmcOwwBkWzJ0c
3lBzHoxfi8Tr1At+ilUesjyZ+BKMleVR9ryCEHT+ELN/F4KThmZw4wUXH+s+0mUKyytyH5K59vgt
YFG5I8H4r8Nu7LNo6kf0rOYwMoGhm1puFnoJ/arfrI+YwS0H5ReyCSbAnMXb3d9EmS4lRweBf/HY
LHvamGgNIlnIj7S1aYtnHCNHDwmZK/z98tsQsxZyYAmo52I+3ym2dWRuMyeAOu3qS7YLRlZuUti4
3Fhroqg3EiGydOsBCqXUlZZ0aF11cK7n5p8afvKVmLxcIzzm9XJbwr6mFb1eLvLGNuXD5hl1t+CB
bWRG6eEu5xE/dXt7mtZH6273fIzWqoihBTfAs7IW9UsUXsL36ujbw0mQhg+wNP2YWGoJMxx3APKN
dsrXtIUKmOkTd/IZKvCFoNXbuWtfy/7/tJ4ubH/0fh6ASlmwfgprBAOweIOPD3l/jIZeb4oU2iK5
xrNgTnSsVpKwf7kq4KsAmRwSigPZGa5Gz011P7nR6nG1uT6MOLb9hQHVkgg5w+qhIqj3ojABMkMz
FpewOv9/0/K7FMX0ClxeRDX4WnjywVnck65s1zxRgM7Zg+eIpum8ZE4wqitSuE7HMzvQ//nBc+Ur
4PDtUQfm0HlxWtIZUBWtCyUkPz1pdMzOm2jn1FtlzxOhnmZC9EdOBu0vTQoay19B+Um4FWARE4NZ
3/bZEHkf265AvCKws+vytxIVnlBg0rtP2z3Q0U6qPNLxdae00MKIb1OQ23nN3cJBrvBR2rfwuQZM
E17f+VX3tfIhrJKJGxfMUq3jPMLACuuSmeK8zGk6C0nTjZ7Cu8ggfD+jR6bAaBh6RDff1FpLBR5F
7XyQrB9VrXxV83Tr+uj+3VLwFyXb5DApkX8lvRwJXmPK7TQDfMtKQegXNCbZG5lf7XZDBOZu9iBQ
W2d/rbOOJ73mXmc2mPLDUd5e73MmgQ+I3RbBbetDOI9j50GnZqg/GonrU2LrU1K8d3qlLpohMqCl
obhqzaARhBYf52fkEz4CstzvM2Qn5JMOYGeoleB6uj/xqZiyjqullYZyQ73duF6iP/hl+s2Qb9Xl
tuuZ9e5y2Bnwu8w2WnNhvq0FyRMA3ohAwFB+rUr+Qa8Xtz6wYYWHQ8wF0rk0b9v2DR1saY//31hf
qmmX70seFtoL2VVYUswlhBXmweJTCAa/kpHhDkw0neNfltVJOQxp6EujKBRsEp5okNYJpslvd3S9
FJ+bDq3vWSUrKa6z/NM2EAk3h53qMaZ2+S4zfPnT3vK2IrFXB8/iG5eJkPgI6q5/KkkhFlPgmnYn
l85IK/5N3oj6kbXBIi+uHbb4ThuDKPGFeJRdVfvVK2ivgn8rG6UAf8tFPIGgFUIS8a9/wiCZhUMr
rCaKdWnCyMTmWnI/fLlYJomlqrQWV1C0HJiOJxOlWIrKAvAgmCSOAfNoJvN4V9IQ/MEHwl9mv2ZN
d3aB1hHzWHFtOUs0lPlifV4ZxIKuJTe7yFJo9iw/YBnoApRrTE7yZdub9jxYgXiSbTcgefBVOf/e
OgVpjOpxYzM6AhwHZZdO3H3FcC4vz25GzSbIh1dTYEEpOl/068E9YMSdJB3FWlzZKRDu7Qq3BXIn
62/RWE4N0zpu3qNEwthB4HiolZGxtcJeVX86KsE1UhIU7Tnf/h7F5iqIomPY2+KpddmVHJb0RZF7
6VslD/V/RH97GDTOzOFQTBydGfj40RPjjDnCuAWS1PqQZZYo0gMaU/cq/Nsr50zQNM9kxrYSwlqV
YE0ZjbsrfjX1F/KMUaIMTE5PIKOirMaO0pkIMT2tJVyysJOEsJjRV5CHbVfkIPaILfstS5XzA+iq
FxOEsglsPdk/LziRknpmBSrjOACrbrfvEXiFzI9p7Qc7XgfkIscB+h3SN0QGGA0VArtw/xgZTeUe
rWkDXbQ2kW+22YUZ2Y46YDzIVilMnq0WxXakahqNzO4Bk1JXrn3xFvUJTzaDVGoCndtfgXqEVK3D
LYint+LA2KSzusbScGcz6x/eYTbj3tq6Bd49xQMkC3zgO48BIXVBMsxXMxjP42URaYpNcUxek+Cb
7Mv2VWUPOJLNx/aHoF+7OX41lJ48e0QrcQiTzzXtkGf6N+zV3xVzZVeJdKPfsKV2jJI7bgEEJBHn
sPM75Ae1VBMDSk5TjiHcnfLYvDalGcaioKTYp+Mzo00ny3bUegdhm+OyUH0L7lg1AoTVS6fmn4Zc
ZV8rDGb5gozntLhFVOJqFCp2ZVfNUMW9wR6RwC0/WjL3Tooj71pjiKTIkuV866O6dmYbBWLk2Op/
2mkGih9MwOcLMqwOhid40Am4NHeUaeWBokZHtm7UeHASSl03B3JFSyF9rgLynNIIrpNHZ1+p5Z8Y
8chKwgzvcl4/Y/vONTSacWW8s8b9rDuQQPDlpbbGuDaacQ+yg/SMlK1SYBnxwp6GpFR3QpzgicjU
JmGKrffwwjC6YpLY1RCxgB77zlceKAzVVtyZzGF2t4oq/9LKS4vtvs7xmemGCY4YdBnAf2/775nc
0xPRQlHfaPmvosm6D4AF2OlOtJHk+r9EklE80wQBj9OWpsMtOg8twK4Mwx3afb1Q3J8jbFyF0E1d
+Oc9YW/zvSypV1lganJs6XLjwmgTliq8ZrACnKFwkz7XMG79KhLVfpxJ7e9Dgv0krq0tAZaROV+H
wrqsRH+tZfYK5Zs51R5UU+LRV75rzcIRdWe+Anxnd/Lt4MVPhJcsgKfSRAhhysgBZsCq0hw/Vq+7
Fvaydkqz5KY3CAQn1r/8yAYTC7H6HjQeYzWRVO5V2REIezJvsPeva+7FrYVoepyIeOOgCW5H3u4C
qw9fFmQ+6bZavtKCrKVsf0fRxbGq9RqL9GAOPQw1+VWm6yvsgNeo2SquqdRhPebORWKMNOMWYqgK
Ybeo3aU76/NCvPm1LzGj8w+dfal/z42YDYvVA3PGnbb/MNM9lucJvygaiPRy87wkbXwu+l91iZT5
rf1di1B9NZDEgkOiqcFu/w7hnSU1xLb1fOyCCltDCTvamDNTPNR5fG7QTLYw0W2PisQl/R/+iDfS
KVtoufpq8Qm1O6yCM+SU55Fyt5cX4M68QGEbbqUqZbrVY8SYtLlw/UBu/A3ei3iiahUNp9n86WMW
+1CMSUcvVggKkQz6cRcSg2dWnI6GO/hMp7hkD1VhP+RPQkKK/EscC64A23HMfTjOkiTChTjGWdlh
5NVlElON5H4ZngszqOMQiY7DupZzsKOCHMdA67eIL1A8XVhfT2rRhFDRkREnFTEACNFMnpkzqG9i
CgiFYVdnlQO1SgdDM+4W5C4Z6tWiIbaJ9prkNCOUwoRK7yvaoCibJSkemPrIfxFrEqKm7qaBhNkS
Mhspy9AZf+UypkQ202mz0O3p9CePH9i8NqsM96XZ54h3Jb4lEJOxYN3rIfc3yV2KtKEkEiKAR0sT
k6wFJZM2iPXxeDvMi1in2GMo47WOkLGbLejUgcXylI21r+sOwIBNlb7Xg8onGvNnTfvxIyikEAsw
L6b+N+GyblsekECn1elbaDAaxN17gbm15CvF+DLvxf5bOJt4G90fZeUCSV85vslw0Kwt5n9yEf35
ZtqOiXTrSE0d0DI/7XCA6rDgKkYWlknbh0DnyAKd9XA+kjtQPg5VGhAXY1t2je7tbHVfmKHh2Tb5
gabuK//UqUh/3pn1HeNulxGDcRKnbAp8zVIgtANHhlhhoZoOue+BiCUXgLyeywfveYAW14UHv4bz
hKZ+c6RgpNA4VuTkfVAgA5W10+qw5GWPUDnPyjO+lJf50zlTAWdutx8G2kpZG+HfOi1fQg0HJaiM
XcCzLshoVuzSMzIx3a9n4IEIOpJYRSLIwrMGN+DqThuYQPbA27Pi5vRW2LTCCGpAH5r9FnKuexnK
ldBK/75YbUUvojk4V6efa+tnVudJF+MmzL8egWQgjaCs24IGHXeYQ7aEBs6/lYlwo54Fx3FpxSOU
5861FN4WerrGpbWb42xJUPTQh2DxSqPfsVQl661f+0V9s+d+JeSXNeQNDXaVvpsti6Jarz21NBrv
ChCXWWjbPipZflUShxWG7lK2DRwpBKalrBObzvh1zKFBChOTiVdLFf9UN+ej3OqNKuS+alHaofz6
TDeRGJJwDfFA67ksj1XPVUhEQXcAY6OW1li8f0cYMLeo+JTRh8Ff7W7KV+9onA94AACXjEyqbqFp
rXzc9LEo5uW03rpU3tP/AJ8lTOG8n4mxnPY9mYfodQ9qyftyHrfgKkbS4LifOxxvlPRKpk4767Vr
A46TxDkFZ4lsdCQgXatpCHPtaGQ5Ny36d04HnPibqP7RW4LcLnWI8jTcJHeYL+5uedTMSx2UKUuQ
FmV5xglRquDYYiHtrjMlxKZdKvKaE8EIc2YyuCKq4+fMcgHDSbWfsQ4oVz3H7ROxCZdj2rx5XNPl
N8VPlhznB4h/ywQr9XhdXCF4I4gqoUjQ8i1oXmKYFQKS2LkPlOKzilYVP7VfUXxmbsNFeBBtJ0dH
p6wkZF4AV3GGMat4z4uBMMd0I0W1KyFccZG/eq53w4ncusUEr2W9lTsQ911ejuOsjySEnufQS32A
R/1bwcfuJ+/kFu+UD9mCOTVMAlL9Zp3CrfSgeJ66TZbIYssjNUk9eESTI7cQzgNcR/GaYyZYhIpd
7bOiqK7RmFS7h10X4AXO6l+cHZVEj11UcdXnT3RNT/6knMRjyynblZVG2aX3RB+3HBEVhx/LIM09
IQkdnGDiCFumBh3FFvYNQ8imatwI3qILWftUrk802afNy31jMdmIOGBbTDkNbV/vArNACqRcpMTi
Ig0ErsRUV01wdysApJ1f+pP4mQnkEubpxnggKjShr49nAijJUjA+26zwzRDzQtlvZMkMTbtgF7Ld
I+rxqogg8ZhpG/jTfVrasIUzwHrcgdyAtCJZPKkXa4fgBKiuJ561EF/aksz3sWqfszwa+neWGI+l
1nBB9fDtZtcVRZFMD5uPubca3llyXPCjbhRhqXJyUi+vjUXMmPoNejCbHcuP9vk1c8AkFZPk8OSa
yZVpabYXZRIUyxYrLs3nuuqME+wYczZ0UdKPIrPSuCHFNV06qYrTVyF4jplDtw7jzluqeKv+dLMb
/xGkyNIpXvWbWra4SCa9sK9hFB7usxO8XeWpD0lh5alCD6vdM8w0wawhUc/NeBeAlUsCyc7VNA9t
P4MR9+wKNEZRhnbX25WwaQzOQjHI57c+3cVWzirOLDbl0u6AQohwTBeDafb2gADvqMOYte0ksFzR
cGQtuuakKTGKbD0PsEfPxQ5ki4LRMoKBycaNgiaECl8PCc8zqD8tIPTGxVwdj/qobBW2wdY6Dvr6
Dk2KZaLWhpo/Lkg0CgVQExS+wbZ9MOo2VMzPwLxQH7vC6O3rheanSKbWaY8tRDZdIWtDm5a8KbLl
TliYTHd7qw1J4Vc205sdLOANFkaZMpGCKvaGjdx5r5gMeIjJjb0vJt9o6RfM2ynoL+sLtkjCjo3i
I3m28dFdRVmKB+VlQ/WJ/r+HSde9KTTGjY8skcm7IQhJivHbOwa9Afz3rZrh6o0RgZ6/LU3gjvLr
FOw0TKEc+EV/Kwyz8IQCsc+dpJoMFFyoZ9ts4AGeHlo/kC8Af2g9kXicdbEEsCaA8WSWlrVrsP6y
QfWNuPfg+ODGBLkXTwkfDrbLKG6zX6pZddTFwf+/BKa6xFRhMIIhseottlA3W8X2gter/YIiR4ZW
XFwPufmmv06mHTUNTLXJ2BdU4Wj863oqbxjJ9CTgLJJbXekbETP6yG1amqJgwuH87Zwp47PG4p6P
r8k9SBC7kTbmYHpdZa+WZNhIBacGBim6OLpx53UsH18Ipy/hzbo7SSzoPBv8WMtDz4rLhtTfmIe0
m2DyEiHUorFmTi468w4pa8G1XYkk0TqwBWep+PQKQn9ihyakaNeF7Ddhq8MCvxwXsd5Bz1v8AoKt
BAkDNdQYaMy6RbLeVAOxP0dtUoUzjNc/ibHdgGvQ/NKhUw/oghwX3iQGFhDAWuum8azOjcdG8vJW
/uS30dobtB94QywfLhNCikIXoNpaMJa+mQL4eXrLwIGeRCOXTayxQxV+qkwaYmVSalanYuSBV4HK
NXHsBmCKfyCBYapOJ6Dzg99ooX5wV07eoaxSsnWxD5tdi8QA25RvVOi2+snw0bJfUk0wCA2zceQb
YIr6zkcmx/0FtsAr5W9aoMX6BLyQDUQSNfKj+H0rL77yB4TgbDeZKthwfedc0T3qZ4kIGah1e4iQ
60BYiemeolAJS6FrcDWvLyZtYbgTlrF4igbHPyRK7qTdCgDqye6Gdbe0CWAT7mZzT9yE2aRqrsOa
srQ5j6bvVLk0gUyXCdk1PFVy1KqlV8SgCdvmimIMp+wKSIS5tpj/+LSZZzVNqbAuakXHG7vuEWnw
BRT1yUOY2t9ZTvZhdACXWWt5FTMVrbO3ZJrmFg5dlA3fuEs+YkInkXozPp7PpNZNnzLBj2fFtrsk
OuUdwoeugn0o0ry/nB49IY3ZL29W71H4F5g9k5qmWvYxHqdhcxSTkZoj6xRXxnHwvgq7XaCvguz9
0avNDrqT+Z8bm2Z62aajFqYjGWPTPt4OqHLHnPBSQ6Jwz7izMxHAkSkyhEogorH521/8nDXhWBMT
0GmwG/O1dsxImZdZczE51ji6bwv3l747QF1npLKgr5Cjn6jgNuAv12X1AflyQmnpSj7SDGSPZF0A
Jk5Nk8iCV1RPSVB+ItvtQ7+iPm1SFMFOfUHH6hko20PYzt+uPs9VQhHJ3TYi/AZLj8lPoOspJtdf
f2INXLNrBL7T8ldVDr4588tUxpzmQv0g6IlDrTBwyQlbWhxgQwMZJKlelLHa+brYt6tYEUN2mARO
MV5BwFralpt5vjWoTd2jKlQdAF1ZfYAxB/BAgDe+z5D34LbeFpW/KW+0JrJ+XbNv5R86GWdNHc5e
6EophtXt1q0TqbrfjIauJKbb8jQ7ySuoieZsT9kF0B5mNHDeixlK7hOwkM6nk4yP/TgV7CMltHDS
z9wp6V/MUpmfuw6det+snwV4jbZQaUALwSRqIoqQWvBdxTggMTQ1ALDI7fhEVsne4SLRO+FDUsGV
dSPOATX1a/R3XqN0Ch//KGtW+FN64/yjLlWr5QpNGAbHsTkDtdWN+6PrrzGVAp5RU5QfRAMCxgN3
elYGFU2L+LNFb3E43SFfo8moUOUyHoKSPITMH/iFZuR3S1NDnKPEh9INAP6p8cXhOh7LYPApUjD9
3sei3TL3B5fv0/9h/cvumHD3Vv6PR/a02A01rapbnkjTXOAwqv8wHDnQsAKcbiM1r48kF4vam7S5
ooEa4/TrJs+YbzLloxSrXiVowR4lwYNNON3JVO8dApMJsAg2FlLOaHRN/n5aPubK3/LRv97kPqsN
L0npH0cBj6TnVmBj+d4WT9fQj30z8mo1SquyzFL6vi6u1L/3p67Idb843KWt396zIqkvPLXrgzqw
jrO/8uvxkYWbGt3w/75eS3uUCRoka1TLYj0VKT3Oq8IRvI5kss6sgxv7DRkeO+UaMtelDV92SkW/
G0QbW1GGZwCYMYBenn/JSnpNACVg3h5wtzj6+9v5+fs6z5XCJAlk8GyYvdQjH/jMaeNRUwV0aq0U
VkWgKjNAmosMj7cKtw5b4d31xpypKqRUZALvDrhLQxUJImviAB2qdSG04GiLyJsRwy7AnPpLBm/t
0HsPizYMzJp8qnk3qi5LDjNWu42qcRC2mOF33Ozq8STxaE7tkf93hUmZCE7XaXQ9HxTTMaqS4rst
y8Jl+99Fx17BlP1/KxIPbwZbd1oVhQcOJzzSJriAragpLqifQJIcqby0e3Qv2eLD90FeuruIMzja
oq2oFbzsn0qj+tfZTtyh0v/1iETr/oIothbCQtl3O6Su4CokTCZTPcWPmVVX7cRCO7OHlFBFRkE1
GVQ++zvpIwzLjTS/U5H6GpP4NiqtgeJ66/j+HMEI7hdGUA1eE/2A1Whu989s/AXXbuiHuy0DBd+z
C/nmdUwZHb+l5offBWnRCMpTc/6QrdFGvTbMLUcvVXxnihyYPjejuGg/JKwcgQ8zgTvSQTw3P2Ku
VREcCDHAMIfVo0fa0Ywkk3C5fNtR1OeD7TICXw1nuh+E11c+czfV+LwqJWnPDM832A124kf5I7hM
I/0CF56TCiOfuCQUxwIMxdmdivsya1mPRKFfkAfqEXEFjdZQ64scAhEpaXXc9AOkADqgzkMBXtR7
ybfwbyZA1oI2uv3XXGiDmMV/lhSqiwtblPMGOwXoce5ELFrybvp3Dgy8/WZ4tKiXbC1iGC/kimCX
xwxrQkfuSU1DtS0GvuNU48ZXBRCsbsOzKYmCaSX6ble3+EjEr4QK+Vkn6HPv6z5ahepqHgTMOmaU
W/Pyl45iYsUBGl/rZ6tqe+jzBLZY1mJ0gkoiMeSBr+wezGtXyztXDB9YENHZxVR209Dn3WQ7vKfp
V3mJlZsZHnQb6h+ueOswsUyySTdSZPDGER/qmwhSEMNcoqfSS0i0BImMdvkDaCQEuPPi0ZriuzcC
Uom+CVfkS6dBnZz8Gqq7bo7/QBfoaQlVhk9Zlx3gnm+G0sz+VXVd9/wL/Xjkzj3kai2BLICC1lpn
j7vuPP7hWtKqSxoRvnbXQFTWkXfnrKiPWTtMpnDwhXfnWH+ux6s02wzHuIh1BUoVbixmNKl18ujH
ERm+oRNXMuY5Cw8fkAHtrNzCZw4ITSkpwdIwIB2wv43getcAx56HKs5sbW4AN9rlnjLJOCnQjsjR
eMw5aJQWRcDnw/sy33qwBfVERF3JoafM7eKxIcfwzDIS6zcU+zf54GeJl6444Jb+nQMJgByPF3Wj
4gQ7kbN1q3/PDOuHC6jxxj7Yfmz4EVCsAl945ftXktdo0PMJ43CvNKhMQtP48XUf690UJasQLPkr
1K5R3kjryR7BMBKN3VZmaq/9UTzsVEgJSD0qUuVVXaJKv4BkI02ZkJ2BfvTflDJ3CWtg4bR1LtI8
TTWK4eg3xS9fVbZtUCQwU5tX/UCi4jN3hnRjy8jJuM/dl4gxOz3pVnQSfnhdo7kaL+f+WwSVXyco
NKe9Jtxqh/EMamvFfrczVHwpSfeOgrmuSWGnphfjJmRKEmd2YXwp1GfVNopMZnefUYFxN44k4VUq
4yTsEfI+XqWM5EiAOmnS4g2WD4XWMrqbxbXDRA4SlPIVfEZoHOBfY7xd+fL3DiyeO7aDG+G+OKwj
HBmc5KqzxGhhEkoWNciX6D8AZ0LypTeO8TpTIAMU18nrQlDGsyH7h40cJzTo9z3vHP4Y3m6dMfoA
pZhKRbcRvcXqxF8Uu4pyjEZcqFgGw+AI7e4GcIp5vFI0IGAGvPy2zbiW4IOzIeQOJ4IikrKwzVno
6LTJy47YjhlUc2Qb/40tvQxJi9yFQClqnn2uk35M0q2Tj8xXsOZsl6PdeI94hE0IIxS4VJeebw64
zV0WZzCt3nCdH216x4VXlHYtLlYMFSQnMC8urHP7ZL4zj8qTSu33AGj+9NHIUzMf+rQ8osVroswV
yJQuR98oEAACyNuBD5vEVud7haUgH0v7DZU7fT33GI22IrKGhvteCTbS2R25HVolOzN1ObSLERCn
otLJP5dmKXSDN70QwSacUi8qjQJkJJ4DRQaeok+bc5hrSrWXc2CmNucUYiP0pFOaA9CASjscg3kK
RuHvZwde7/ATdt+fTtcabzaS9HD6gKw3gNdHSTvXAOw3RV9khTgxYIUpu0FB+WRnWNKTnwf6DHOj
ewKu0Gj+Aai+QI3HXkN1ci1C6OkHGNy/iEn3hRxKB/0DcIkrxhCwgaqVOMvPAYFpj2J1PF08p3US
PRpNqSWqmBf7QOFLri95FJJWI5S4OJQfglxX6QnsShqdg/nPJucxWngmBZmxlBhl7OfzfoK7x6b7
v/bnaLxuazSldDVCrYPt8xU/AAGWpuOAzFs2k1W2K+Cau/ODx28sFGL9ao4Q2k5niIGHIoV+rQ4I
MLkyj4fuorRjtri3C0DW02iUpm2LT8W2ChFS9RyvgTcyQa9Dhf9hPsCqtJhCOhbs9tiDxG+jzgdY
x+XaOUtYJqJehoWtagBAZ1PfaBPG6M2IUywcsd3iCCCWNCWzJq9+LneB1k2xydhpWlLaeJjuIKWz
PootKUTLhxga4132YRDyorVBQeVW6dqyvSijjuc4uXDYH99jHBXVtBfen36fnujOLQQinBq/JWYj
kY9lyy1cXpK7yeZe35fYW7+c1ISP6/WFa3W3bGdaJVqtA1HOhqL2gmdKhdvrEdZ3nykF4oEQCpNS
nfheJfaFVCcvhlW3pC0VUf61eTogJ4QGZEEWpf7jSKEkrsGkLcGovgc175k3gxXD1gn9Bb2JhjEu
CjA35LSskG2A8p24ANzVwHcJPn1+XODZpben1jCIae6zdlzFc5C8/cRZztmCVEpc7ct4MLAnnuQn
/zPaADjU3hVBOGzaXhT5FI6vMy+t+b3VvX7WUh5w1H41tGBonuzpW09keyIRfyvFm+e6CuKN8L6s
GFAPRUhNGLFd+mQMf6qnJem26rG4NhT+xUjngH24zjLJyQFfwRGkePP2z66BQQzcV9VMS3Fr1om1
/6RPL5aOGS1eYa848YGeXtCHQPybPUlclkVg9eFOwm5YStD+eYClhA7Od4lE4JcGFviekSVqEToE
z1bKVZHAg8/Dz+h63lqnhILIN4uWhvvyigLyimjLwhQ2PKR6MLSMswQrg/vznmkgEE0Inuok701K
99xvtsoCFubJ+frAst2N1qNnHg2TY1ud/rZH8Dz+1xLn0OjhW+kSt18RuHJZrrSAH596NJUFgLbV
dYQaG1huGVuptDEd9qVeg61l57BKAXwFXYl+tKSxNq0Hh5sOIqWfosIo+9fFXwkLAcCcYb1WRIry
gEHrEyZ0+XyB09/yCtAniFA/TonHIsDQh35xbopUBhHMx9reS92JbCsexLEbOC0GTsebBm67EuzD
T2lD5P3IbTg9EsQsAtTNbjNKyfMUZOkhH3H6O6gk1e548nWApZ7Rs9RGiTx5EOPdgJi6JOAtLMuz
u0f3S/ov6cWdWag+K4xxFBANpIvRpgbVJoDcjp1zW6E4yNvvQJ83LZw7LSDOoNV2U3Pl3RngI/Yd
RFRYc9lGqcUUtpu6rgYxcJT+6MTz1/7jPMD5kW9yGtGGWGnVtJfetrmmWxtnJghbUIkySlRxfu0E
t1D5qeL5t6CVYwleziP0gHCLP7Dp2xf5XoQzhmzOo3tTeRzBLveUkq6mCqscff7ypOvXDMf4uCRF
FGjXEA/MVLFkm6cKGR6glKHQaLOm9hz1gPJOcpkxwOA7jMFNeP22HERxXRQfqyDh5OZPca/Yh7/G
q3y5/LOMABKSnlp4gdJMCEo4ERgNXaNr2spKHyggRBB4B96MqiU4eB0rEzJUTZ8P/vKf5mBydcI1
DAsHU2Q79WZlT1T9PTcXipc7bAGR7M/l1xRngT4B8i75JJwGLQr+OHenUOepBIXtt/JRiVSX0/Kh
z3j/UX5gMay1eKsI8e/eiUUK8lUieURLcgKON+797O4pErQucn5PMVURUtsKFXofVFpMRQnOVSxx
EouxOt1ysRY9x1PA1Io3IU9+NF14RGjkvjQv9RmlS8NElrdPvNYaV9c845gA8ebzjDy48gItz0Lt
P3Ijt2wT+UB6LtXLcsXHckD4w/3xFP1ggGLsHGVHbJDPMzRvx+FbMWhv39+TYW8zw/TnjVuGIfwz
74aZQJqMXAbFj+n7jigyeFga2sGhY4PqdJKAVR1BjZTHCvLAQBHNUcAJdnDlXMsfiFyTPzI/9Rha
JD++mMCy/gXRpFhHRVmIzSIPdd0rv5RB55ppir1jvH7h/vWRuNqmyGU+ejwpxZ0uDys0LDoY18X9
tOraYP2oL8Bv6bq50sYmrfZSI+vtV9uh21Sza0BtM1CrbWq1cnpBE3JaLWj/VbVtt2JC0wkbfVY9
tZRdZazEoDl5Qcz2fLI6MQWoAaHabUgUG14Wh1zkWJWWlDtVnDUU4RYVz+Hqn9Gee7Xb61K/O4wz
YUrD8dQEv7Y3bxzn/em+BM1fJ19J/HRxSFkUU9znW8+85WSAWIYyTQdsiltmt9DTG9l3EyG0vgmG
XI/thj0PxFnT6o2wMJnNG1qQs6rjGJWgcswDzFwR9sn3O74OHUzUwvztAOv2GWuTWEyh3uN4q8yd
kuRA6hNZe54LLyXFpuDbIYpzQNvr2mHN76/btnAfVmY9LBMhPFeCTnBdNmOzSfVu9djvs3LKvRrb
PXAYHNAkCf1rxe7se9tZTqGqDtnWUEo8+m6B43BMo/0E3727iSAFCFwEgrVZ7Qj2noMPPKc0rKn3
ReUYUr4tIMQPhrpfQFUxD4x0pYC/zh+5miDhxBcJ/A4KNrN4WJb2O2oYBHYJ5sxadbFig6+64Pbx
heGq9a1fRW7+58djSPC8rTTXoN6hRE5qbB136qdMnN2f/rVkhJ8ABjPjGneO6q5X9FozlDqr9N/G
JGhikZr2Kt/KKSxecyQtWjE09ATF2WD348p3hzs4s8c2xmOv+P2nBSWoeS/vCI+xExzzJ8IYx4rx
249x0XbYVTt6jiO+5ypdRqKV2NVdObfan7WC8McFrgHv3GbNb8/sTVxKhDNqI1FV9E2yvpTRe5GK
e/0zmwE0C1AjopBOfgalARpRWmeoathcotM2UVtP/SvugPM6N8j4J/fngtc84Jp/2YnOT9n67NhA
gDCOMP0Td4IR8YbCb+CTDlF5lyPNed+JA00QqC7ZPEX3p8445jSL1KIhrvEDEwsX6mvouUx86gm2
xZgnVGcfBLpFckpl23xPa76EaM8XoMe9lhSBYbsgngN9EhY6YynwkT4WAa0qfhHtUnqjaA4qmxlF
1yDgdQBkXo/yizb5UlfzD+3/EL5Cwt7i3ai2kTPfAeyHZ1UItZ3NQDsWqfUaR8ug9/7/T3a78uKn
A9NQWxiaHQsUzv1U60VD6D+lQuC2JCplBUIXxyXHsiHPuPjgWGLWWtIn+GX9BiaiARb20lg3mp7e
Qdo5WK0lse3PfpthC41wWHPKdtUTlkjSMkSBSnq3B2o+Ftaeja5Wtd87xTsscfzL2YfEky47LUpX
08aW1Kgoiarfn3v7/I08+qUaFDCn209jtqjZBEo/iZk/Onlgyt8hRJPy3UxBNvMSErlBdoP9t4Di
tOj0GZ9e/SnaQuIsLq+qtxWOuUkf2TR0iO44qUtWDLqgb/BIchfGh4OjeNPq63TegoyMNHJElLV2
y8+/xgPIq1omU5AzKB+eoQL0CqkzUQWCRCjfCjuC3FKju8qMJAKWtntCCcjDEuysb/oQzeKoG062
+9Sv8spBkIzcu04hNdnQQd7g8gSYt1KchwIQaqQxnmyB1Fo0f5iGNt5IdghwqSOfOMYDcrzMxbzx
fI1dwcKJAk0Pc0SjYkQHEl5fTKCkP6MV4SuNjgxDkUcpUNLDy3IkWYD/9PzcVcVoUITl/SEbkL21
xRDO//3tJbHKhNOWszXhn50YoRnCeHFyA4+i4Pwn577wzqfyuHgOVouf0wDxVzVEFnb0Q0myEiHI
VUr+0xmH72o2M7EHvUQ0TJcEgjqnc9w0a3WbJFSN5Fp4Z3LBa9Kx794tpFQf4YvhL1OtOt2Zwcin
KP8eI2UMIK7SHKCrEylFpw+wMVitntH64jpiF5FU4FBj+bl0zAV9CXoTp2s1QLbJh3GRg6pY2w1r
sRvhJdJLk6Q+5moRa+qBFH+0fSuNWMlj9Opvjm8LcQ7HnK9ioQeih9/NPkgVnRk3g81kvs8Z7haI
SzGTV8u/2HzPIst1FtwaVnHuJ0FHgWoaoz+bce9e2xfXicXnTUfm0sMHivURAa3Q9zSO6thA0Ku1
BjjCSiulvUA9xH3ku46BvG/cFo28zomLjltW1L9/zXLMuvQ5ftkl7RfAbJhNL8A9HOQ9vE0v4cwD
h5jqzbT2xvR+WE7/m4IGkz/+oJ0MyiPnhzk2mY/BYjMT44oRmep7JMy1KAv4Xid/0oRotDi7QwTi
L2/eIpjXwZNP6VvT9EXOYgZD//+LrCIow5ykQ7RC4IgVDkeHMG8bdZZZs6pL2TpUQPnH5HmpAHrs
4HozmBvfjRd7N09UKf7fHJSnW+SF0fo6Hm5QxSgNnpkLHRg/rKgn3C+OxzA1zQKH3+QtjXh1xZOr
lTMS8ucghweKxsxjRUOJmev1zMv87F+yD+1/5XY9P/mHJmr1Xwc05zVWZPCuT0r/fKF+ffsQdNTJ
wYk7zVK63+WC951Zu8wJAh18PwbcDKKIsUN9LvTY8qRo9/KlalxguonAsxw5HdUI7s9RPRBKxjHg
LKGjInhgRkWzPrVM9Fk8V1Invup13butlIM1x8wfWqdGeRMEYk5rsd9ammY0l4Yh5YBxof3qUIal
P3ULO9YbW1U4fjD71CLoNVm+hNFbYBaoTcixu7TJdLNnV6qllfzEE1wxbFWn02GUCv2CoHH9rdqR
T1sq+KcCCHVAnKSzphoUvjVA9kuhDdQg5a8VVlxO5lBmigdW2OXHR/I9e/elbI0Q4utm92byOaX2
w4S7KkuQ2XvR5gvHDY3LyxHsGtfKjpUFAFwd472fn3kfFT1FGp0Av2rBRyA8kjEUTU34tlv8luHL
hYlVZdboLeEz/PPRth3eCb1iUqywjHGKLztieXseIGVJaV4VeGhZHvh2Ge9ioQw6kX6Bhml9r5tm
O53V+N+cnBynLV3h0RNZl1aidDUK8ViWOt9h4q93XwfANuJ1xG9L+zn77Z4L54jpguIaFUpIFfZC
U0hntU3nHgKjuKs0U/3qs8hbTe+RgZS0WmA49GCIp76g+poWmtyU0ZTM3bkTf8y5haxv83a81k0i
cWunh9awSEThPLDzEocwaCH5RPUf871IJS3ugS1yWbxkBeme6GRwJytHjjDSMLYuHC4vOgvxYfSY
tH8xLXYUuAw375nbYdZM7h/DIanIC+6xIf8Mt38L0Mv4BxpMlUs5PB5pyxWqr4POs5mnQ6UiI98Z
Gu3/cGJEid4q56QpYV9z6aOuhCHW6tCFLqg8pKIS2218lm2DClGMvFHOnQe27x+99tW4T0KOCHNp
f0t659gENvFOsFg2QQkBJ0Ln6UOG+IafRGhrLfXERulglPZHAZOdVWZ2Q7+Jw017rj6GOAvseQkc
ctSi/3zYbXvGOcu7YvyBeCWCpAMy+vcP4bGMJZLnYBHd9/0NkUZpnUVcOSUwStGTUimt80gE/XDH
Qr44mKgg3wDt9N3/Uh/cb3tAnZEWFTgpNOmz5vOjEPqgQtbuoh7YWps9XrA1wW6Xvmsmj0kaUtoE
4zvXxR33iGdUMfbqmuqubKP8C2iYmeYFHJUWflzzUsSzacWvPX6ToT/aNlH55IbztRBTka1CvGfo
dhJqCaXyzCqjuYmGT6zWrVm6XqXM1RqnA9aWqvQAeyGafvHejB05SxHU2EEfR2gqKisXyOLueu6O
gvNiX9XjEfg1jQvUypvub+h6o+X94MJiNnCqZH/JP+wpIlYIt+UZVSAUMHutLpApzm+erncK2kbq
UITi/BqDChMsQJz0eKqAvGFWduhZbJEfGqWSMLTtZWQ0ei5SQc0pYwM9yzsQDs0CYcTWRILxvJl1
NrB/jkuirsXmmxBC4P0EE/lSo+bjB+IMLtebUSZvW5scLCIshZGY85+2p2Q1U+JZcz9YhhWCIZSL
tUGuqD28Ujb/k/ZR3ukRGg5KZEW6fmVfHJmucp+1M03y0h7xN9IkAgqexO1cwFee/W+9jQGeyZI6
T/pCed3olIrs+IFXo+vXwvCqm05YAWhmRb/mx/UXPlEQYY40iDHJeVY6oRemJ8OolNHLcnGG1Z4t
isNNoMFtON7AyqT/PZlfrncmjFMsKdcaWo2Cc4Nu0SOeJBfzMCI4l5J+eOdHttmk7qgTT3CARIxo
FshRw6dZI44eYHv284uvJWwKm+UnDkNo8bgpTCYesbseZizrd1ADnIsVrlokIWZAgkPYxsrBOETd
k8sbHRcxmrvLzdbDzv0obSW5JlhOZYzQtXLXKWUhKBtjOAkICTZHGmXjabkbFejefIQlyHksPr/I
Yffi/cSGWhrpM+MfWcAllc33Y0sNasab2w7f02mL824SDPd7tvwcO8LSIQvoyqINE0CNdcjWMaVp
pVkhCp1xe59LHkb+Vo8uF73yS0HDz273ff2cwyWwreqlKy372e1esUYG71Q/dUE//jF3HgGyNGYR
i083E95P28ux6na6GHEnpjWGzfPVVB3gP7ha2EznHcjpqIVXrwrb9ZkSg6e3vvDSOwd5LAc8O60V
NExsI8IGnHeQqtaf7W+kq2GEJwOB8RUHAwrBkrgGZykNkA2wVfmlusaVErI7Z4opK2eyrrxnh1n3
mUUWdry7Cd8CTQKm21WtFR6TDpzrPZa/7HhdgRW+H/ctuIh7qen6I7Sa30acKw3Esh/vzEUxhsxk
Fgr4UaOF5WgDsJvTnE5OpL81d7i8KV3E7y7PapQXnoNQ0WdgnsX9ESF5O6RI7e6/uSK+bg0swzsE
7P9XTh5FB5bd9RAgDXATjjiNQHNPpUa2ioX+WHQN/aMMQUcxqP3PnoTM5Vyi+QoTS4DXZ8i1m6jt
dwSi4fKjMIL92uou+mvlavZ4syk0DYt24wHG2B+dfsYx5K3b2Vg8KDbzzfSpNIAPH7LT6WrKYVsG
mRZiR3aaPihz9HFUtqNLlR3/6e9EBpbjw4mM3p8xlqFKjsysJwtieQs/r8VvYNtK+K2aHwekIyBs
EE3m+hwiIdvJpoYvEYzev6zzqgRj+fQtjpboWn3zjyRlI7CdFE52DM6w8hUkTc+rjakOSq4T58KU
0gG86S5+6hEjenaBw10vX537pbK2DDTRuLsxgiVb1dhWLr3+8G+bDG174A+Xie9st7Eoo1LdHXZw
rDg3JgHxq3otZD4BlfqMyV4nbIuTqUbDGHMqROeZ7gMrbRXTknXvsmWHXdtBawnHOIpveMmK/BMh
PMfwlwUQ8EssgG2GTX+1C68pr6svFOUCxKeFyq4X37f2cDSBMwVTauYMuUsei72wpa9XCmIITDxj
vkSm0+SHLCh/JVn+8Usi+ZiRpgHdfzgazefp6GtN6olKFo6vryM+KY3rct18Qa4BjgRPvwRxqztr
cozC2u+qyxl9kbQctBE9hOxvalT9bAAtrbOk9LQYbgSnp6TrK5EQsWF01bH2tmMOFSqelQn3i8fx
YqxS5ngikawYJTzYPEOXwGj+aHuxdF+VB4qltZKjyryubaDdQ137ocZX8CM/9hO1NPnfh5tG2zf9
yUrv3/gPTv95szFb6OGG9zwuAYLc/4EvY3wxH1vX62hYrSCqxrTJDr5RYz/SnSuqmBNCWdlBeQZX
yq8jFawLspOp9rry8W39eI2Om4mip9qPtzk6328kXN3UXx7+8wgFtpYdL3Z8eqqzLi5ezpt5CIhY
hz6MJFSCN8gd9PG7Ev7kfH8yMC4rc04/LDwICxISos/3DjoubtYMFCNdOstqwe497Ne46Zbobg/j
gsPf4uCF3SsA5irm2auMHzssXONPM3H+SdV3kdiYsYrasjcEDT3eeaW42IuRDuntFkDbmcgHwxVR
Yex9rlnc5IEmZiAVzfyKapRqbjcxs2Q1aHXvaPIXNxap2i/RD8pdZtL7lguC8kSFDUtp2RzwsZO5
SrNvxEsdt2TS4dXSsRFY6Q9RLlKp7oLWyt3A5AVZovsiztPIlzNn6fC16GSFfiDdbErWJRul2GtB
yAz4yVcf9rcrt4W3m0A4eWTui2Y+hFxsFu/MjCdFQOl24jX9gql5O5unGqSJaTw6Rsp2FJirLnIB
b3Wmvn4QyxIMZazh177Rw3CDb0QS9WkPwAML+H0gvyUExROO9V/Z/yCjKnmq+toOlN7In1AfW5H3
YPwd7CRJOcPHchL94/p8mlyAIXGjdyz9Qolby+0TVCdYoNqyAJbIxjVnLrgxBk4jTonGGnaH8RGE
mCnz67sQIST2jU0Jqn2q8+IGZewA7HzRCs5RnI99SVVoKcZNq66xTMcOFo8X5cSlNNchdmy8Lb7y
vFY4iY9KrZhbG3gpEWeOjNiyCxUqqbLr6c+O1xdc2hLHFV9UwSfesfJTaUD6Z1vfeepNFEy2xkmo
nkKxU5/xF6XeubXHI6WZEYuAh0Do49jIMMAZYRzxoP46szX/p9XWszDEBtF63L1uvWW3p/H0lGHH
7uNL8WOTSYi3N2tRLNdPejQaCnhZMKewxic+FT8gqBVsOc8DKritSalwXp8grb8n8G28BhlvFFju
8TEVtHLU85H0JTY70QMyOSInSgMT7NNuBlwMHH3R+h2xe/yzv5iLWhoOALEe50Q+EkJCMKNDXUt8
ztaHTajeyDwoNkNB1YwC+BpL6Z038DFAwMlKsOdvBzOyTekXo+NdkW7Rir2Rn5LW2IqGz6/+Y5ww
3uFpfHpc/1PJrHxQZuzoNrgNX1Wtos2stfpnJ6laJh0hD7dhjS8rO3qJvG+QRm+7+OY0BtENeOEY
RXMdCTLRDyW+FlaYsw80dZtGkUfo/6/0IEPvZYweq9zTKTGoewQIAdJVm3adDuGW/lCvYzNS8kZ7
nvaUuLc/Jnbvv9N8y9QiMvBtgZLNlTeSoT8R3GaBLFNBvQuIHJk8rInVyxIwFD3swRaweGEcPFes
kcvqFWr4HcEPV7I+AHM/fShdZHKUEz7nwERKP6zd2OWQempN09w/WJ7imniyokbA37j3iDZilRJh
UpZhMlL0ZV2T6hdlSLbThXZgDDsXH1AR/XHEMsFhfKDCOh+URpcYymkTQdNb53mkNiZakcZWZw/V
4b5Aj5vbTpmjUhEm0L0e1G8gul9eG+rInDK3rIaiR8WtNq9xeABOlClXuJYDkmAnckeS/DPvjbQr
EvwzN324CFdpEtMArhWspdg/4IOwxR/9t+dWr4xtf5vLl9muEG9jGC856SfnAcewHPlZ4PCZeX3a
hi9EM6hCBsf3J6d9jdOgynCJkVBVZPemy/cNQm3Yq1SIAhj4Qw+9ut2he+TdCUEJgiQjiChDzy9l
grwNiKNnTdo3b7EJQx23cMGXXzoatJc1fRky92SPURQR6+d9RCaTLFY6BM53ARKOZ7At9Q5wDmHU
8tuyTCWGhr+D5Jdgdnwf9h1oChQtmyjPKmG+JhDn3HWeyQHNYaH9hW3mLs9dwkeuA1h+vpfW4Bin
COVNmdki/fgfrwGKtpkvC1PBCVDQCwFRVtS0dqZJ05LYvSAVd8xE4Zv+TCO61JFU6kf0Ys2ckdNA
uoOOCOOr36RukOeZTIVGlcF6IFhYlmBaaOodCv6YJrn/sUMN46bJb68xb2MQIHq26uVFh3ibp4Ov
zqkfieDLHf1Run12MTfz4C5baiRih07TEfabguExmT5eUAQsteROehyGupOOMt7uVRpENP/SzjdI
7u2PTCAwhTlk4Tj0N2yBiqdxuHzh44sEAnNZrHAuc561q8ngNFLPD21RHFWaO99T0YRo+mlyD1bP
i7n+GQ41NAF9dXwRmb/Shiq9rIUudMYSXUsuMF4J1SEy+hTCcjQkuQ5KBcWoSip9FqGcsB+9Jh/T
3nCgLzKJ2a13V5tVEG9JXB4oxGqDqTHOGmVVWe0LJg29T1J04IR34FYq+KQf72Uv23PKEIz9GGrm
AK7RfUP6JWkPtdBwcIVj+DTyWz1ynhNLukOkP6D2J/ZQMeacH2x+9wT7UdhhJrTVFaGKDLLj9tzX
sSGYKRuyk9tYJW/QhfX7UKq3hgYmQz93KdhW0lkfdqzPtDv9g3pI44iTjCdJlnwQ46KpJMmIgqHN
A38jLc/9bEycpVy11+y7/Vq3P+HhhmUGQBB9F718uRV66XXQxs6CbORlvZ6+XtNZqVX+pGy1b+cI
nt/WEniukYLP4ao6RmYc7zcZL/nL3vuYnK3JArLwtwpvzqsO19eKRGnGTLBM+il+a/TNixJtKXbo
J0CvrNBZwCmEuvh+jMZHM7XE1+XnRkGL5iLHNorGpPJ7a1eEKsC0iWXYazfEmKwXRwoY+mi63WDr
kyZ+joYUIkqczDMTzgVRVDr3fPNXm+oi17E0M+GOgOVnd0i1XFIUoHtAFD/jVQjAVFsJyTjQkMeH
ZuioaMIrHCUJWZHFjsKmFwa6bCMB6jwoojssONkejlSJuDmCAznFKUBGEU7RgyVqQdO/LbDkst7f
Sq47Al+z9nbNa5+YKUwzl0hs59RfkFP1ibcz1gGAM6Ning/4UGlxRh+SNGLs9nuAeo+i9OgASVpR
X8dr+D5sSZs6mTbmhUuiKLtnX45xaSIhwzAcaYWZN4V719iqLfqTReX4bJNse0VL7NmH6YT5GHcw
Z2zg633hYMNwKA+M64Bu9mBiJqdFQe9okLpA/wM0u4bcN2wuHQ6EgKxDbL4BnH6GXKP8J0cIf4dR
cXCYYgX+cHiSEVXE0egXCw49YVYDVfqutNUTFcFwz9hRuRnYHjJTsXRFWAfKE1dgZHa/eE1mKnY+
FHKOSnj2pfTtFR5px5yu/eUkibT1lrIRSnrXDcL70XLmrpg6R198vlF8hz+01c6a9JLfyeiRi4h1
YAbojMncZgNjIALB/F/Uq83tMO7U5X0WFeYUjuHRRT8/JLhR+jBATc5WHBVFvpEcfzYzMOqrv7D0
AuAdJ24fu35aZ6E8u3g4GhHSyjEvxdSSZjyqwavV5CX9/lsvxT8dxI0WqZbiMnpkZCGvt7myFErI
M/egZlVZr7kKb8OE8uf+o6YXUEml/dZwp0A6IZOdxLgFp5yJJnlmXum4rYc+tA0pznC2Ieu0/RE9
OBbUWmpOI3ssg7NsnIsOVuErnDeglxY9SitdKIBMGNwGlXcZ+XnjsSSfGoOXNDXIbmvmMkuELgv5
ex1zdtqoFI1e20dmCN8c0mmsEONg0YZml0cSeg+T7CQ+JzTO1byFLvsjepk2EbBzcQaSxEC2ARyE
66IqQp2VZD+hni5M62uoIx5q0IYLNUcJz5a/uUfmcsd1ClhDpSIA+c/Mv0IJznDKH3LdCK/dixgm
CvpouWlNyzXaP8iUccEBTK0toly25te60bMxL5ESzROjUfPjYFtZzBgbbyoHDZg/qbrQ6lrVJQ/q
VC5s4J9rgDMB7x8DzRzeIcIvi84zmSGqiDE6p2HMLZgcXs0y2r8iEITFgR9Rm4oVlKcYCH/fntMU
qSHDE9kGV9Cj6z/1YOsBIVWnqWkQaVIVWzh1jprs0yEaT1tp1hFhjNVt+tDu3dtFm1Lk9ovc3lTZ
FZLptEf9NdW8VE7MLxzOwuQdhXqTn7QTdrOUg91xC1TRPzWEIQXknfF3En+CpGzLIyzvoN+7vfyf
znOxVYhab/QHcqz1UUglLocOh/K0LZNmbHbkQjB2oaoTAhU9wRB2gjnp9fVIt+uUBUJ2TDnB3XMC
N6kXhsXv4QlZz3gXx0Uq8g+wTIK/K2A/Mqn0krr4kGbiJVKGdlVBTcUjEou+NmF/c42Pnp44b3C8
uQS9BVpY4LmsJgzJ0o/8r46PQB0eBLnIIvEPlwYF6PnQZuk5vXAN6uwsq7IPtWg5LFtuzdciRs0V
cEGK621G/ApjHGpKXB7lscZNnXdkrWtpZJsQmR0DkRRilliFFJ2Egd4WBnuOLEI9s+ZUThig+xRJ
LtcbBiUAJBW1d/vkQMZiblOZcAne2HDrkTW6I/rkwTxCRppjwxj/RfgKWbUxlKXonkdjarE5StWM
vue4xV5SffP/xBphpPsL06fYIS9dhsy8xIGDC0IN6PYNJFYMsfrG3f2Djg7O7mVQoNGaLTxyYfBO
0QS5s9CM4Ca3hkf7LVvMP9ZJgpKk3tjYGfHNLG+yZXvzkUDA8oVlnFNtR1vPRojwbu94436gSXl+
Z9OylZO3Ha2a8LAJpFmVuiv8Y/rxI8nThYVmCFnmvw7SNz6e9bM0Pc1se7Y+UWEuz7CspVfrRMr+
S2qWXAQQPFoB1kvOuXNp9QN+F4yQeWvBi8FcL/tR0+hmBcMt7Ezh2q9pT4gkvwe/Z80Bl0RB4nzB
vu5RKgiZtBUDM4ivUCMH0Cul7rT/F2yMOfLJJa6D+ppJHuv4F6Brbwc1TxQ7qCL+OBhUyItxAcki
2NZXrPCiN9p+cTrDux5YaHYVrl+V9xV8u1Y+TCE38n977IFMCoO63EK+8zWMSdZk0oG6OceXQqhY
JIa+MHjb0BOT7FlNyfl/ECe8f6/uJ5y+/nMgmtIsjdVro4j13ccQtB17+ZotVkuJrQ+I4llzgM8k
gubpm4BS5WjLe9H5gGzYZ+XTHnG88rqAPyYIo769Wgf0aEkFBUuDWOu6kF9kf35vuqLUhdRT0AJ4
iC+qYpQlcY0y4dOlH7/TekZAL3a2joGqpaJdQ07tmVv80b8SLkSQKT1dlPwrHwzaDB1QDvrn44cV
MtiUBC5SkG/6caDPJH9JOEuenSaIY1kGArtoltPqrNzVHrXlbcirSkRaBjduxQCplKSDKayfh0cb
otmt7UGBE2UIr0mrdVwiJ5/lU5jpuHijWCrzqbgQ4Rnv9SuZa5fJLO9cx0BOpRdUspbTSWVW86Ka
zcI+qyAqBU5w155geSzOg365LO899tug0QAAGn05DZ3UChSTAW5p/9BNK5W+v+5YIZdCFOFG31vT
wsl/qZk3fRnHb/hZYqYzozAOi20Hdv+8YEV6DtdjxBDmeOm+YsTYXKAvUKJaZAIp3ngEZsQzdJ0N
iRott2XXHdHiFCjQ7JeIW/XvePiU8AwzaEtzwNXEB6dzhdZ0bqUHTXY7tkk1Dn6st2n4MFEuuQns
XJ1bkLLaOTjOFZVliWTOIRB41f74/fJeyLxpCFrfaRAS3DIaWFLHJCoG34MQEdzwcyTZ6pkK+FV/
hZ+nWdXJCR13JndNktJKCxtKUFluzSPWBxTArtMQn9FXA+ql6H3GKZlcOSzZTjMeVClYzlhT2fNp
tQbG/dfHWlZasAcnZq6DMmRLEylIRVViD6GFUeuPhQCyJTt/g41Vlt/5e0pDdS06g3pOfqjKleKV
HX1W4q80KStrwVcp8dwhzRgP9YKEOYbr3yDX2eniUTO2CgNyT3v2p4mobrGq0DgckJeWYI/r2uf8
LrKMVm1E63UT9NrrR1encMOeUPZmq7PwNWinNE9A099hLzsxuTSQG2Wg9OrhLf8M0MrsHq7WwfLT
jZXjgO7alyCRFdO87YKaMeKkb7m2DZJDIZ7DARjkmvyFvB5U4V1afIkH5AEE5VG4bk4+7j7pe4mL
DJ4pqU3WUMOwcE+fiKcahWpoJioVVnOJ6u9/RKMksqyun0A7TDgsaYqWDnyPIQdK8xJAyRhBFiyU
iDBPOpVCPtqQ7zL3Bfg+T3oNcimhjcg96hA3n2eL6AbpP//uTFHBq43Mdg/vJKRB1kd2mmDrGfPP
YSut+E+xpXpiGBABkfmArbAWHO4/kSSVKCq39LztlpIvNYxTpnEC+MqfD3R8V88PNym5QGr7cs2i
rFRPGyMrYUoFaIbkb8kRhD8Z04RWz8xODmIFx/2IJBi0P/rHL4jzlxVZcyrvVBWsAd2inpa2hsXS
lUVqeIYR6etORY1HjBjmt8YMBgrdF1dh0SAuc3TF5cyCKTxIp/38c9UXyeZEK4mrqMVmqJ5akuNA
PVTpcuap9ZfcAYnGMfxCujFRH+vHpoFG1hBe+7IJvGANT03oMTBQEfkqsaByY5R7o805OncG5iDw
DD8qU3obHvOccX2l/6nq7HybWG7TuTgFb50MkOslnqAh93qIaNGxfs+8Ij3s+G4SOW3ThFXv7b2F
fNyyJiO0YKy0Rp1a6jRZldKLzlNB+5vAMZg4n6suXVrtEBRCYHejyrdzXt1kuurHiwcgzQgc9Yjk
5fR3M6jtGoqeP00AYq6z/crNUkDroAkoocn/W3l/PKpl8Ak1lutZXGdOuAEeCIctxSVnN2iW4jGU
G0Sj1SerSrgOCe6/oMNG6GICl0E/kOdQt7VSB8p5TYe145yYIJbaffOHR9bdatr69UXjrRQ2lc4z
N5IxysnixxJlhFEhbBGjq+LiSUp1SBilykecTFVQFnxiD6wUzINiJHL1Q2N1AJ6l0QxbbW0W6pBN
4Qc53nm66+g8N5cLt6yL4Q7NGny3PbxW3p+lenU4DM0jihYopOOdb8PinYULTR+L/O0w7Ihx3w7l
XL4QRZsskfH33P40vFTwoKJYVYgjM/ln0U7YgEzNuNb0pdLjLFfRLN9D4Vsyf1UBJ+Co/g9Ocf6L
InZg2qocTfIJLxcl4jkmnpMHpFa97iNcd/R4UluwHyLNyfZ+q4OUuZANbYKN/v1etNZlLvKGA2q2
ejF1OC+8/x8GLQUAJQGk7uuve9x+p3z4W0egR5msBaXKMqA1HnMKkytMw8y6SLyTdFSDHVX2ti1l
7jetwm9fKoHwfhmVnj9S/ZCrFNgC05kyasiCI7Ughl/Q3iviYMdlXd4+lac5sXPvLT3nJEC2W9U8
mEtDyCpKHNHPggjMlIN3phaDsxuhX5BId5V8Iey+DFkB2OfSjkN34RbX8KPU3G+FYtQ2SeLVCWHI
HmONvSQH4K1yXTCp5fJ6OZ8d8+twezOY0DdnenVDYmE2dt6ryVb1PwRI3csiWcoRt2gEChOJMScM
4twAkjeyOFrTDfa66nsFAThHRzzuYW8OA+khNrfZNmEfAA3eyaLnGuvBZDNtZNPEf3Dnfd1/GkWI
C+k6uTKXihtSHbSAYsw0iyZnK6w69MoXUELut/lGW++3Onwd7g2vt8tBmxXYPLRFTFv37DcY2GAq
fCAwvSImyVCeBxOnzyVrLg64ktava1g0anfaaN1yqH2Si9P6fjwavQtLL3MbRG1ZJOtZbpwlDeYN
khLAOyLFccxUxW26fuushWbM/l4emw78OwVuA89Travnm5Unv9JzwRSNyOvrk3lLCA+07eayXHCw
2uC4Vg/c1wIr+fNSvK6WvleU1dGfO1JG52lhSzCMqTxTs2ckXsQiH8Ntj5j3rOLQA/sNfSBOGpri
33rsDIYYAoNTN/G+iuwi0noKjLK2CDvIGc7Bz/pKYXrzkYJPXpsRLo+AtMrlHlPrbpsorFHsLDg/
/pKeM7/JdiUsDdhrQAIdFTQMl4sd02co1reqQIeNMXhjO1zJQW9MkbP2rtSNtjHNGmwboMGaMUIn
vNYWJdwRo8wf0qIr02FcD2oyeUL6dTQ6qJtk6ZJIn9N5BDUJ9ZNxXx0KIle6M+UaAHe73u0ITTxw
tXCf4zzBw7CF8YNS80Cmz2oGsWL4FVYy0ButvJJZVEEAGmYOdx0ruLAR1Eh+tbhVLRMJXBA90vk0
pqYcNQhQHwYj9W5MiW7CeCrAqIK6mVrQjB4EpsiM0IekV1wHCyJ+EeZ9cvZORaX6Q50BcKEzsMTg
MNmRHx6d4NlHZoYDySxYrNVQ/X1pLYibKLzbXSojj8kzk/5NWCKzcRRHfC+/SmDHlsnuTwqeejXZ
r/HBO/ZWP7KuPmJzyQ3cvKZYHEK0qL825sIjPIgKsacdIaAlxDKyJ3LOgCinDxLETcKwoUtW8JGh
6N91RVroR64VMY6Dd+0yd/CYR1V0rWsqKY0Gm4kKpIjOdzWJVZShLNilXlIUaCo1T4vVV4ulQ+8Z
a1By5GjoOrApEqKWxaGSSK9GETj/rDPykjitPZC7f6GYOb8qBHE69etmKt7k4Yiv8GN2BZYtT5EU
nR6zDY/cGKvJ4mBFGwEGdzwI6MzifeysbkIEC8RnoGh4JjbwmI088VxZWbDOKZqAKIDuad+EVvp7
8qGF7jHOU2WSpI1b/0erh3emmdKp7/zdi783kqmp9P35+m0cWnQBhkHDSNcxFcgF60Kd9oV3sDnK
/hk6QdHMXAcu5uEtKgDY7z9EjI2Z/X2m2VOK4Q0PBOWeGYtdiEn9qmX/1ZIVm8M6MaxxgdkkqXoQ
y9K8h/pQx2ljjV9oMATCTrcSE1FxwUkE2HUeUaAnd06xk5Lf32ad5JD7cG+dIa8NxZePWVwrnQGC
CmJzFCWmGS1hxVwA/2fuXZRrrcnG0OtnWwgUJqAxB3CKGlEgMy10UqBw69RkWlrWVeWEqvitlrcK
EvUqtF2zfcEad4/HqjoJKWT79sTOQ0DLWQnNFoaO1VYDvb/rqjndwh2uYUEPw9dkw5D0n6kJx/M6
MquUsRg2O5bU+x+zvP/uXRNp4Gm39y+xsepc73vF+Ybj8o9gDDu9XinIYDQ/yeWpnFVDNgVsqnpV
INGLHvua221XYKMZ0hw6Ak8VB+3OcvwC1+iUcbbeY59dGVFh9VTpoQP4dyTc0WucB1eQiy5KMbNz
q+NQ0N9hQnBRk6wXTI/I2q7WhpvjrstH8zBiLycTtSIp3UOZkL/9viQjy1/bdEf6Ztbe8O3C7bYw
VAiSffPj/YaB2Hd6V22fquExElFw8doOeJSbWaU2FgD9Iuu6uhJ/ctrwm0U956IByx33r5dQYtSy
hqLabR3H4CvhoifvQHYrbmD4gftsZdVRlOSdrYDnJdIIAJEPwrIDxihaO0lYVpZ/2ouwcSF1Sg4S
0Vr5w8qEE/gND8WEPRxXTm75tTTt0yOraPDG84okYvdUH+56OOXuzKUlLV6P3wythkg3xKZoxJ09
QXEWVoskos1ZKbJN+Q4QqsQtYGsU3mijXNhfuAeWkPpaZCIyouRmkHU23Aj+Z9btjRwSj5ax+PTQ
CwQkd4HFe83PSMZrS7QUxunAAHjheCz/VxMtnsAnXhDwXzxer8ZRZM+CdcQQ5BsrtAV1iLlL1O+M
fK0tFjshfX0RK2e/UKByLrYn1kHOjpemiD9Ag32d3Gp1+GQqEmdOeoVUYKZMDxV1XpW8yjAasY6Z
OxxEdJwrstYnXBUAuAKXoZhQmrcf1RbLc/9XGK2U3Av0C8uCre7YozeZmevRM25Yo0fHatOo2E2H
6FAKmio8OzdGiIxEZ/AjFtLox3ft0jdiRD1qX1RfG3+BVB8aO1XRaHuEvku5SMwOrumuevzuhWzH
vUptIh3Bk/os5FgRcR6eXFHmzVW5i6LcFBfl166k9hu0jhvAMno6wM/U6qysln2b48OG1vzoUx+e
QDbUPhORGr5Gu2ZMqWRUpLefQ7KaXBOkZjugYhTtH72fjxTbUMpR1ZWedW6KP1ZvAKTI3Dry1iiU
GEICh2JJWW1d+hjm1lq9c+ugSgrLwo6NPgQW3/Qmbm7Oqdjf66Em+hy8Tp4CVqzdkQ+2USN4AEFn
v6TixJmr4JqVn/6LPgqXxQWUsG8dAJRc/DuCC7tw/c+yf1T8k4NnXahL0I1gdtU9SjPBWwVJSlPu
RZYYyEFRIWxttsps1ExdyqXLltVn8ty0m1+TUXp7X1yukjlPRDLcGLqC3glnLkVGPZ3nkc0u8qR3
1idJAltaGg71LN0KNTiIbLuE58sCow2vWRm7ytCbftIbXNhGhXK3BXs0U1ZaKJfvR2E8JwGgwh35
SNymFiZF9B3NpQdMDOnvh+00QTw9CsOlvbSnG/HJyXZudWzlAst+5d4YDvFMGCI192N5AIXCieoN
Vj/wapvDbp17A4AYqBlp4sgqWzYwCq9wz+8RqYY8M+tTWPZJQMmct4FfFY0GFFnF8iz0NHTkGmR/
ykikPBhIsCmMVM1vvq4lWPRF20Et5fXqFn8Lrx0bjKy2+t8pJkzMYdpeFZDjH1U+0h+UGvjYSHYz
wckY0Gr21Cg9xdLc8zYheSoZj6Nr6UyJIv8BP8YOejArNF1tUSZMJWm9piqzrzTsXInPwPvtmn/Y
sawNWcIMrg+ks6uSvki2hx3/577aXmS7dRXYeGn78fLrI5Rt7Vk38hI1qqqS7McjYimTpt22tg5S
mzdaGWdiBp97sJGoT635rxm1mQByh5MWdmyu9NK9I4EzoU/a3Zz0n16Je9/9VDijSx5tQRow0LLq
Qdb7dWv8kv7I9u579IYNKiI1UZbw2X0l3ApdqtRW0FfHzeUQKo4NqeJKAKgz+q6TkRN9vuht6KN4
bypfQP3ex6hKQmqXyiPsYymzhpxHgTsUSptUkc2qguzepU76n5PlAgTUWOLbewtKAYKtkQFmz5v5
G3WbDNnmoENz/9XJf4ftScQNuwWgKXeWOJ8/8YdGjC6ZBZuWjsFHVcb7WsBLd2aGfPrXgmY/gNdj
uLclVEb4JJbKUxvEQIRHte5pd5YHbu7GCZuncRM6/6jJ7eoXC2E8dFBvhLy4RPPu+KX0TGIyeBiK
OwcEfx7wy7jqoFm/L9wrQrlZOUS/MEp3wyV4KlKA+YrpV2NRMvcNRlPux6Zh0Qi8hsO5emKzb6Wc
nROPWXXOCgAAFFSmaGYwQHgSDzAkg/ZoyTRlbDvY47yZbdhS2EEEhRpzo0t/Lf3Fww93Gt1LUnp6
lyGhRyWM5cCEtjXfL+q6Z1w9S6A58Flc6bKB7F0uRg5Nsorl8ItmODTHyrrje/RXOxOp/2PeeNTn
0CINgfPHzu2wWBcK8BCnh8n9umaVFWzBdI0hAFTCTnYkvne+o2lE8UnJ1jHJB7DK10G570ltzw2M
AOqfuV6HGLdpV6IEVAXsrUvCVdV6KhLZFPxDtdSH8nCoYPTgya1dXFmY/KVVXwvN6yHjwZeEf3jW
dLmN0OXWhKQs9Bi+gKNX4dLmwZZZdUrztOuiv1vEC2EAlPV1a9BFOlXTKNijgElS/KUfk59piAru
/zg0T1PZ8YF4YsslqoxjD6dzVRHrhuFKA4ej3hHAdPgzg1SXZJSBPMkYvSprzDzj6uEtTkfIE8WL
F6wB3IDsalb98M212xlqEHKqNkR/oL7bHyeLgiXQ+IaQp5n4Jsp1m1uJqRSNVw8RDtyzBhYEZYfp
/atSTmkwO8qfQbe11Q5qHew2blSEiG7DsJzVqDJ9Zpw7wJq3OWdpkjiUD3nYRQzXAOauEpMDPPkd
nn9tGM2OMkqP1PGXAw3k/XzSET3qZx7BJAbGyFZPby5c3uN+GGnKav8jtEEEzpQecFuJR4nZd+FV
8iK1vVG9YoA+sS/OBA/xKZjmPOSZVHvfi7Zj++uKLzvB7/rXnv+gKY7DBQQEUogx3yYrltaccQJG
LYGpLlTkwFS77V4TzwIm2VFx5lpgua20hpP4YU0KjPbdJLpggdFcfFTk30PgiWDPr8QbhF9HGAmW
LMBusACSyxymqs6bAf3ldlnPo82pDV4boqtiSNIiW1ZA7zObMuPxUHMeSAmomNXlrPhKcDaomR1h
8rNO0bbjsyjnZgBp/nLi0rYLMhpg5P0mpLAUjUNLtUH7GhGB63TkXWs+VaulWk83xk0uT4/1l31u
QK1aGpFxr6lFSXooVesEFh13dSlgSkttX3dmfyzkj30uSY42aKTsmBQTVTEoEzuH1tatbgbgSKTF
9FPiybfzDSZZLDxHUkpxnYz56zD5yWxnPiUN3DWhKTE44RDt6v+uzdr8PIoeBZY9FlWQOjp+EpKk
3sjoRf6fJ+bUlp6y6mrHjoFgWJCrzjdxitUjBgFwsQHt19Sijj5jtJ3PgZJ7Jo8oWGMzE+Zq6h23
bs1n8epmXEOR9wHoKO1bVSxGQqzF+iNUEagN7aWSxiHPRBIUZta7tW35Q3I2BL2gz7VrPEI1AwR8
4yFFnjiHGnrPVVrFf/Cg0w2OLppye2b8iddgBVHW68JOW/EGvpH5bgUL41muEBOXJ/2AvZ5sibIO
M7OSVDW2uNfspFjyhWAidabiWIMuZpD6QVygDBaUdtz7pS5NpUUAd3ewFwYpx5UwPPDl10GndJK9
7/0W2qpZEXVj94qlh2OssjbLa9SnB5fEwG6DlMOAuCEL3taVe2giJ0dyuv0SEk/VXAYFTy3WTIQy
G/2si4/J2UE3WyDbcaJhyBG4kGVzK7uzGDl64OP+sizUL07I8Aaos+gnEbGh1LZq2EfaBnQKgYWA
3YATeh8KKbk122yvgkEu0FO6XI9bTjuRavnvjHFfOyiObhrerOamb+Rnn2MWd5DerTfiEIZrq+L7
Wiu4Mp94AMT7vC5+2ZPHxNGIKNuzkwc9wFo9JaAYIlVmoSBB5QP9QUMt9bF4ybJKN7fyuv0paFPd
2HfvhxAsUnaAEokJ/CUKwm3KDsnfBlpFnQtTEdEOvz54qjiThkjitu2DINvzsJfbP1HlnxkWKVVR
V+c6hODqKPC3mUzmcYDhST153C3AJHLwVGJeS7sJXzkOr5TmAOaLzm3giLiMEQRHthrTvvJQJ97X
eQysiEcjNn2JKCrLX/Eqp4w6UOu+ZRVJH6Pe+6o1CHspEPA189yPO1lxpaunUEqytPtYAFo/3dYR
7kysDHfJrew8QhSwx3cHR9gpXhKQCXMZtwF0dXFtOWbLo9GmaraaRi/guVY94yD5o8by4qJwn4YP
fCiT7upIPuTVtABjSCvFKqyt3+rji4/2ASVf3dVyVg4ay/VazY+wuX03PTuHrwDlr+nxEe2IBrPP
DWmYXAr4gvOzrBNFBiL/UuuJGoUkqYHGMCBKVRinjRa+4ATi78asfnbccVS/KJmRUB2FXd7aesJu
mNZA9ZbPMpKdXV4Yx7v/6Gt8S2rGcdrXl0GHTQlKrCo6Rvwavr4OM7r/852ZUS9U6SPoGZgLLN5J
Z813jwbqFJ0HgZ4gGb6fTT9LHtcNRE6Wde9wL0wujUwfRyQ7KQdWPWL0iHPNyI2jDuvN2Ae86X2u
VQEKfb1ARJLWyRdonggNiTWh8Pu9JjY+m54hjOBas2yZZiuo7YHuee3fBQ+m0Pdv9ye74dLDIPR9
XvF7pokkPIMtHeYXwwz48AvFRUruLn04snDs2YnT5HCVNzF40FJEcjePfcmG3UxXOZoL5W06VTGU
lnnuSTtE5ZS+/OJKLj26BmCxuFuTYyPun3dOPDNafFi99B0Dzg4Q5wEdmBsghMmk5jrCKh0AwG1I
c+PVBj15qaUoE8PFua564GF9HzGnkzT6oa/4jGP86Za2RAckgXv/gtkVAvMus7uEk4wYl9tOooiS
MUal5auJ8rYotIdbC4mtQSWapPJ2L0MuJi2zvXpjxJU7awssviM0zLIeVHn5P9Lnoh8eZZ0iGSj9
i2rJnP2S7aGuJUCt3VDT7C6WG8782+Wss6DSQd9sIbUD5nWXqP5KJrnjml4/SdYsy/SDCAvCIu/K
wo81v7fVdkEysZLKiwNLLKGYGp4VUE2SCUNSHKlzT/jPp1AxZEqDRbEICBPozURPKFnisi/Bkb9q
9mXr4c6Zqmq6ohZZRR3cW9d5BlRY9HQ9chQOD6Zj3ZzPk5QvNJ8z2HBQK2OuvbfyoIpx/MSX03qh
5Hy6SqlO/1GRhe0KREnfenjVNbyuahIhd9MdwVzp5E83aF25iu2GcCn3JqI2nBvSgFYjcTmNUGga
Q+EHvUgM711tQjadUlc72sVvCmx+PqU5ZB/NT0lxHSl8b+s8NHLvcYX5I+EVZ/FY4BfhsEHWZiy5
wdE8oJbrlmWfrr0EPHrDJ3xHrrp6FvEZJ7sq53WVa4mZ4BeLxOXTBRz8S09SKVcvjYsbOj44beE8
c/BSfCYSIMrsqK0ugCzz0mZoh0bTtT8hb97d8sen/zZlNNDkebv+G473Z3fe18iMqcMMzzDzoH1h
nUDK/N5KW2n988Q7pawyVoLN4iCCyfvuyWGtzmYn77BbE4GpLcVnE2K57B5ved3nGomgvqvvwpAW
lbw23d43uDDm0jfcX8rJYD/ycY4iGlRqluU+c8Z3crZjQyl3Z7yGzRHY8JHBRHD7DSTeAAvnl0KV
EMrWWpyVfo0JLWPIQ+z7eOg4RP9UWs/YsUJqmnSXfChiiXDELEVBs0Ul2bJStGOTUU2ZMGDcJxiQ
VD1qXR81SVYt4Yav9WCdujEhL7PUgoFymZYdv2lny39MVaX9FvBXEPuIlvGKYiMpP02U693WxvEf
WAKhfjqgcSZLewdB4Ei3L0FkYnGMKlH+XlS05nEZpYQyvPrVKCTNl25M/QJcsXfV/AjXml9xeznQ
ZpDCjKqvaskLtvKsEV3eERQbJ8ubdYIuRlJ34W7MdNxZyhMdI8AQ2nj4lH/vzWstZoq1x2q5oRKU
Sd4pMZS4HiwwIkB0y/1LYGJRo0qP+hP4oF8vkkvVN9+5pXHUz19kZq36+JlcyQHrKtjN3KEVLrB9
xwdXBhasp1YN0+YQDTZdWDc5ewi45TP558SbJYUaroh8mEDfw/9gdLSpOZDYXY43WntxEbJwKOYL
vnm5KO6QkenBexsr3eP3dnYZuxfZpEMPLTgQ1ObZSnN/8/yQ1U/gEXcpNnHD9dNhd+VMJnkYsddl
vbvonjfvXebDPZ0J5ITMYuYuUyWpSRy9+nltkIaz+PKlW2ytwMBq4oqQxSKlxHYjUErxiG1mfpSt
TQIXsWJCnvNmydi4e2w7zXxOky02B1oYJzbkArJFGQjK+APJsrbpijZJGDxcZzkp5AdXgb98cjyi
u+b/yEVIDF/0L9zSDSeP1q/oSlxxXwSNq0bNb9bkOmcK531TQ50b43GlzxNuzVUtCc2tnRtOnE6s
7sB2DBYhGBZdEx43hsXTy5BIY2ljkna9YbuSRtYkB9KjdkRbRH8LBuGXh7fnGMC6q6zCCwbT/taS
KBDxALPdJTEWrTCs+rCv5EAXNDafCRGP1EWeTgc8/0VzVlmObqQ4Kc97ODTNCQteENxYGkhpqAx5
XQIEKiS8zVJzcw9erMoK3WccgoDqps4moIztt+Xtrqh9iqh30gnEqqeryv08dKePgJ7zz+V/e8nz
U3nI37bvIVc/KZssxXCf6jiu3YYMEZnYmcNTZqeTUTvIPZRVk56l4Dj6WwpP4uN0MgHEoy3etgXK
p80TrmyJxQdRRAIZqR4xplKct7+th2fPsIDF1GZCPzdH86wXlB7wPuyGR602uEQm1swMl0iDIW8W
OE7FU+16tXfJg5T+uwx4XJDeeVgx3P6jpQhsrAkcKFHZCZHoL3coKI3Um/U/9mxesMTCrBcJVKiM
TaZBcsPDVE4WzN30mgw3adCgTvt4K3b/ocjvdyKZCZQXhpxUlUXhknCF8icA+vbDqlvfgy44AKj0
FIyrGxO+h17X9Iq0Sl2ocxMRscL8ZPZ2XWwUl9u/w4amsYxOPAwtVea24ypC+pZuItxhKuQserGN
gxrCVYikz9sUcMsHf51C7JQN8ymYlVWa4BrpUxFkECcNSxOsWJathEAZ/TYd6YoAOZEwjMVwbYjO
etAsQnrhWOiGztl5syYTXeRZ1JU0Vyzvx1+R/Asakc70XhaJ2yIMIbAOXdiO560uR0gazcjJyYKJ
XK6MsGOgzypnwlvx1WXabVrcsl7hjBgJ3DJUreeXqSrr6g6NLKnbUpTgayCdbQ7YFycYzcjxdemS
GLuCa7+meseCqM/0ILi7mQawCdswnHuL3PG6GmYeyW9aZOF/XnKFwZsdE4xV1pVNJfBsk9oSoWnC
TGBshoLfvLLk2xIlEAWJK0kfMQ8DF2bUYusD9lQO65zqUUOESQeSjXFsIQjKKkPmunBPCutrud62
yhERMcoGv92h1zgEOz0z1I1MvfyKrarujSBDqC2ufCVrYV2hqjQCUrX57t7n9StB7/MtRqp5dGMu
OWv4xuxkUWYNy/fD0aGHoeG2hw7X9ioTHfEjr0dCWaAzGr/N59D8Vp4ldRsX+RuWqivfmC/ErJ2O
1tRofKQEBbJoTz7EC4WDqi9GU/W8iIY3Imh03KYi4YzaYuIoB+aaVWNj/UWijiM8GR+OJZbUKQzh
n/zilcTXUwCR2zKjUDdcVZmu52BkvONdknGJb6yBGqVKA0U84En7j7fVKOgb9hH/keQQTjN7xCpy
nowfEoKuPtl9yl6xZI7MDSMiruN9Lv6hRPHOYGMhXw95vNVAyqfCKSaAdDfjGZluAL+SNpdysOjM
C2iqcA5dDlvytmxvcGZ81NIKwBBcNzkDN+21+1rsbxtLcWjqfca63K0K693RFVaTp5EtlxfIetHG
RmJwxSlYCl1kZy76WiXLICFJzf64l1FiBLdnnXF+R3VBTryYTwDawClZfVvZ2HSxO20irMGQmiHk
brVMylwpoImfR4IigTKmahTJlvtAh/CVm4ROGLh1LGTyD58cBEUtlnyXv8FAtyNmZDhJqsj5hAg2
6Ss8PxubR0/Cnynh2PtsnxgXgf5wRgD6Np8ZwF7b/UGr49HIaluZBq2WXpTS+NNz98/c9J0ib5Ic
c3ovic5AYKN9DdV2C/bJoBinZW0+PMiNusLVJyEBaqzML09wqzkl9rxgLCRBpzY5eJ5nsVH9aB16
BI2V2TJbqDJzKDONvNcLUQTpUkB6nEWCgmxtd828GKuQcN/WmX7tSReAFNTbfEclaglkn+bDatay
gztgx9xLE4s1ysEw5Ao+Pggm+satNWjq7/InH2jH68JO80ugbMh8XjvIDhQQIW1L6AhYCKp6vDKG
QkEHhqcF4qGg7YaBxcguGNXoS2eHWp3a94Ne7JAXW6+Z8cbAcQ1JZa0g8ThFkkuc7fRhNcYjVId7
cBHPyK/vSRfIyctHw6G26PXZl1Vffgyx2YatKdvR6DLlH0UZSjtZs4y7VLDZkvH6KMrvRVolVHA1
l29sBCXQEXaNzgyV1Nf0VlNvQIgqTmJvIZ7bA2WB0EI7VJkV4So82j9lo/74P7kWKn1d9uKnANDR
V29r5dfebmXYU9Wfktfb6AlGQLUjbPLNjMKKzdkAodxBYa9YgYws3QDV5hfGcLcEnjeuki/AZbEB
7ET4dmFJ7PIBx1Dusp1e77eAnG0dVoHUVS3HpzcIK/ap7yTRm/tkcQ/uj1DtRYSPULBTTPCVzuA9
PCRy1ZwR7tqKn2XJBKppQdPkfJwwR7U2TpMC/+nXz8u+qzOxdvplbUnRUWxgmTa1MlIaZTsVaU6V
yFu9241g8TViRH233zoNECWjEtGMmLfzjhwpooZdcnyPAbwXdTRSXet9JEsFskSR+6ZD6QW5wHiR
OoM88R+3gESGXytBSqoOahaJM6itdrAKoZ/eAH9Mms4qXPVusMXse2Jb8XGSiF7ZQdnRYS8zEEFS
Tx4MZcuDpM2m+NthIPTVdszKe//FfNLNhbfIvBJPawyprM1WoS5UuKqx9gbo0lW8YhbNlsnxHyy2
4UW9hftE3sefl93YUQ9Qx+BSy/geFBy+80j1ubi0muVf1wiulj7Cd81UeWGKOhSuPR0tWBzfU5B9
Ley1vEWFiOYKjMx+3BOLvxOwKOc2iLzna5IJmZR5pme/z3Ngk6+xNMQ9eHIXB1eZ30XTydC16NDM
mJb4IqTNpzYwUPbcIa8M/soSnjDBmFdElIEGzEiGaI4lyJAIwFZCzuChkJvi1UecZk/gvK9lu/AD
67IR86o0SxVMHQV21ZJUAqNHqdN1y9lWerIUG7oo5Gt/Z8Hvr7LZg0xWE+4Ihpvpq0F30H0wew/b
TOxEsyKAhh/UIvFDzKtSvxagURtDLfvkO6MmekkSuH3PRn9ozXnl6o/Luvaibs02jtr31WHmSuZz
CIvuUN/vJVWI/Y9jdvM/dQ+ZAftd5wMVdG8pHKInwNa07QNaxauiA9ICw/Ze7U211zm32lGe120A
M3/AT9KoYekpZZdQka66rdDCkXTvnrRwbnYW3QtG3168LxApBhDLOS5X5EV8d56xPGWRve2EMfYW
dFwGDp955q8rP2+m68xSJTWF+QOHgTGTZ/MqYxN0jn/MZBeZt+agNn+rCvESkgCGPReOCBP2bsUE
x56wMOU4GJd3UjZwPlpfmCxcic+/RogxtSdjXLu7JyXgc4ucOhf00RE4uxQqaxy+2ERBMUI92llT
GqMv5WzWm0lVDt/sGcEuatrRdvThhu8cf7/ZwgofVq/lvxHE8r/Biy/CMFmznyLvX+8U6u7wnKH/
rN1HC+bo68zlHq+t4Pgq7kpHKyQJp/fpjE1lplWfi2SSW/6/HLqnfwKSYF5QnttOFlca09OBDZED
zpuBzQVIZPVCHEkJcTB9b+f/PcbYFnMa5oQY7jLI9PVV+IgBcEhXLUaz0f2ns5ewOcGSQSKtC5f+
kmgDF4nKln6lHggbcXhWomD7njYG69WIImxpjfwRQZtjv3pRg7jCQXURm1VlLVSFQXEqv/90bOH+
08wglZVt+WHVi/TXfnxzTKq+0MGOEKWjdjfFASG+7SZX5r9+Kr2ypk6aBU73HYN2ulUZE4BUXR3X
UGtWMhdvSuFgVqqAnqqFQiONqeQ+EU/360pLag67Bfqu178q+v7GSACq4PJrPpsgzywE8huXIAZ9
JiXisb3RVJK/svM+YcP/Ih2T1FNPw+3zAlaAaQUP3L9/NsgPiLBLSMV9Ti35t7EHmBaNQWevwVpX
nyfX71YCLyuu9EcXJmuQ1j1MJMeaJF0hU/jbVB9l68xEqXq44nccBV27RQWA02D5hbn20taOQYwG
rdawk4CF3lpijr6qaizn4mkgQ3Og0g+tM96l+uBYPVtlUBly6kk5lFIbwkHSQLHATEKSsOF1MK52
Ox5qsPZAvl2iCb7tNyW9tLaNVYaViyYIIuQjG8VPmf5mMTn25Wk34isQVoeMZrCqqbs3BFXoI6yE
2tKWa36siumlGU6hoUhcMxOVuUHyCwPdTI3kqEi/45RwbG2mos8098HDy8LYjA0bmmGmHC29/SUY
XuoUu6lJPww4maoAyE2XcbaI6wsEMIPAasgFhwkvTKfAt5ZEt6Mqy7Qui8OIJbbApKvcm3bfhulZ
pr9iwErSWh4PYJru28mD7aqd0jR06q58P6lHJKM31WYTBDPMzookGYfHQQ48h6scziF9itd40SJW
Dgb57nyaZxxR59q9ZQCV5h7GwqsK7fwWrlocikCu98VEk1FAgqv7ScECkUMB3Aov9fezFsLkyKDR
uB5nHqA61duI3lonssgjZZdr0jWNzr1EfwEA2+iwrhEMfzEfQro8BaABVE2qkFSoTvmzz7c2A+LJ
axn4RyupIIDqwsWLtZ+kxQpl5E2EWeLW/ixeddz13NQYA+Gi+Ndj5GHQEszh/38KhUClhUkbMwcl
LI13vQ+W6qecwzCD+tkMLc8DsSEx66FqEgkBz4oWT4Tqsd8RDZ8wWCv4v1n7t4S20e3Sv/c8Tidz
upcWBhqUd3Ub2HCO6jecFavJ+zugm0JkiiPtLoM/1US1IcCeVTBjFQfLpIHHefqKNtbh1aLiCyRk
bxv00YTAWhsgD5NRTzN+64JcehiQzpg6DI49cbsoG1bT42ZZIEbljvpoTsYTVQcTUoAoiAN4flMH
7CWeUx6MbgAdflgMX5VUEgqlifQ6HiMu4jjX5umkzyswYgPHvXf8d66pVvozDMtufqfuI2/21M1+
F8p6R1K1J7pVN0FpR+pxk2/FMY+Ae81cFGDHdeWzR6sX6fhENatp59a/HgFvwAARS/7QykEbFcV2
d1x1FpPmbD/6y8I/DljMCZA8YCL4MKxwrXJRqTTLXIa0Iacmp7LS7FXSn4kXurpuq2LW3VztTa9J
RFmO57wI1DHOvgOqvRfiZajcViK6rbyo8UZ6Zex0iAu2mXW4/50koRI9fErdnXDpor+6D3DLY8/v
srsc+WpTKxHV9RmmFryy1VofZoZLNyx2kB3L8zeZC1h0+FJRb6JQeZ/ICHMVKm47SVQ9lSma3FGm
70oAIFeQsrtHwZbd2jZ7HKSERE/62aLQtVMueOGPRJn8YsR9yb1oDf/RWT4u/VzTEv8OmaNc4VJ0
2pAXnsg3XmQoIcwfFe09CLLf8OAEde7CM69C1ue0VIhBbe3/0zSLKgyZNhcMVyhVuMURjt/08Vp6
g6DMW1zb/EfJoyY+PVJH9wG3y1dWq5FZ5nLNpGgw2Tl1gzsS1kfkpR+3rawz6xHdfFLBEqIdVqTA
HO4ri817XakHOpqW0spBRaBBqKW7+ujJviieNeoa9uzHVSal0BFqr1aIvYCFfAqmDSZvnUFhFwNm
tlFPJ/9xHfQpLxOVHK2rrAqpWA5xl/NDPGPqtGIfpw9qNFnazMUS5RwF9pTZNC0TNrf3PlR+WLDA
G2FCVZQchkFqtNRY8SCYdzPUPdN/D247qP0RorGOtEYSLxAkQ4pCw//xREyIZ5WPhuK5Ta8zuC8Z
mQ4oTg7t+KoXybUOAXGehbCD59vobWyUOhnPAePNk2B2nRLzlbQfIzHCXxDRP2pR4lx7U2mYIkFW
vUHJrNSQBDCC1G3EOeKjJsBxbTxufaug1rdWzj+azx+7DNPIjOBYlRZiGbgd6jEluFUke8Krwdi9
W6OK38mhGULzftCYX0oOSQa4p25m44x8a3kWygR0Eg/e6f49oV9SjTIfl3r6iyCkXYvfyipkj20N
YhlZHiQ59EHkea46oH0vEFzpJP+3DAaixin53NFAsqEiXsjV9VwpDF/WGLnSNxcK+4t+OiZCurJb
jnkm102xQAwCu80D+cy4Cr6w5SuUPxZ+7HVdCBPVUDMvEM1bl7a3p4X3ldbvIpfEyA8P4VGaKPnd
TCKP8/tfln1Z7iN36/GU6ewAP+JbTe4RYfPz5Y/EZERTUPlt/iMAfFriSxua/izHml7URdp32tGb
/kpKhJHmcklrOnl3wG4npDLMMuMS/jqIRf5cZvxEISIEdigLVF4z619/Ctmov40Dj+7ohd2GAZAW
UZeUTRN3aSnWhMyt0pB7GdZ41lZTg+XbyabJgRmpwn+ziE9LACTDrS+5wRUFfMhDHxwLmp43qzrj
7xhZEOayhHBybJXjpQXpPgWov6dGfda45YbJHUOHb65Bpj67VM2y81VHopDOju8pFnbtF0LnZPtO
jpCqnu2edLYtgHOLEo2jbqVJzQwTiS7+6gnnMY1ImdKxR1ppt8IdhetXGyoPYk5iCSfeVPpUzd6d
HnrJx8MKx3OKlC6+8VqSRg5RGcPiXCjYb8Hiq3PcQMy1ci2kfTGY74icCvrj3hjBK9UjoWGkLAF9
T7cB+CrHGiGDCD/z/mppE6muwg0Jf5DBbmsmxgjzh5B29GdbxiJ3eQp8VWoYG8Y6mRH6GZdEalEK
qQo9y8iTgAt9k3nQNhj9y97go+WhCqKC6QbGwzUflAnGHJIKSWDBv9Y6Os6xUWEzN5tPQ7ISK2fV
GC3IyXDisl8UqAdk4xT9Fe1U7zDSGrrZe6Pqs6LN/zW/jcQ9K93iZwD/ROLRVZWmximn/N3BCj/0
zbYruonYCmyCyzgxP1ex2RZn6QaGsrx8c/DVPoWivI9n9EGBQ6n5Q8cNt8AzMBNoS33UG6b3JVe4
48SAGuNgogUMmrAupgmx+JU+9I6F2rZWHwbolX3AulSbReA4gu9FRQjHbPlH421QhGZqZ3ojKtK0
n7aAFZKhum6Guj42a8207Id6x8EKF0s9WQmvrWnSGIoXlJC/Od4tYSHWajwAs0nZ66bqpRH80I5N
gVmBM0NNY0t4JeQ2NCoB8bE0eoKk2MtqgAxSYgqUVZF/TeEzCNGxJSx3zZfIH4F/+ZoU/VvW1add
7ES+P5zig/QaS0QnYcUCD+EWCcSVnvlV+11M9t9UHGwURNXfiUn1A/Wv+T8S8gTtdp57Apfw9mKp
pyBqAWWn89uI5sB5MMHG6fifLDU9J7QZ0RritrVEJPpvT25jCU0afZNrEbArgGErhn6ePTRwSbFj
ogRdWMAwztIi3bnJSBfzvZKySbTBlky/q64umqONd8LXarR7AvETSbWTE0CN68QtRhCJr8CQGR/K
cFfqFigOQ4TL2M4Vk6cLgK0R7/0QP9gSO2ga+ZkSncRea9P5+U6oaPWMPosLc66AyymRPX6Qiafp
UwePFwMyF+CAOtFS08uVCs/0d37TUqd7qaw8uWcVnxH+UrMMsYc4bQNzZgDOV50bzzm2sUPuA5wk
JVZzluVwb/8yByRG0qzJRjy+2Q3qBu0skHgRY1Ky0PKyHNupq4ZgWfnzlgPsnezGy+LtM16QF5Yy
HOnbe/1Wzn5qunDaELAP6ZOs1uLUlihV3n7FbnhN2s81koAU3TppOWQii4WPNwTJ3oDK05gxKFH5
9uHGaZ85tXn4fXeoPn20s8ySngbW8B+7FD17FXWsw0GWY92vCBiln9m1qtCgL7xLY9iUBAoMVdVm
4vUUzDj/Uf6uEWn6TLVvsCYro2jAKD3nsnfOQCs00e9osodMAqM0+9RhIbNe8nqBiRjQBIzt6d8A
PsOT9iwHjqNpyJFEfAK3IbN02sv9vI08ZflJZtcRXeS2RO9f0TJSdU4rdFk04z411cifHXHUaPRX
95PeZ5lnHb52hgMXwKWyrt/HSQIGgqZmH5172nz6qyN6ui9bF4BHbkowe8Png/QINVkRunvfVwc7
XWmUSpC6GfSMqOu5QU1bDtBoS8wJ0DoP/iWRIZM9KVdEuTuemJNGTlRGZkm5OrOInqybyjRJWxpE
ynSnHZsDEgoOTSPiaKO+I7KZPJQfmsaD/KClO4BcQl6rNH3sLb2a1TvyIKGzmh4ITitsd+HsU9gP
J3k/4mOyDlBYQ2XeyBK+gwo4hoSMU0wcMw5axMA4CtSp00WN37DhY9bw0DQQIaYGToFFemWcaplm
rTyiKSP8rx7EIeNATLIt5ic1j3Cb9ppROBgZoLQ3fY/zNycEBkFuCf1XgsO6nqAXGnc5SM7jY5BC
z4QLw59TRksB42cP9kG8EMgCsiizvf+CCbcBGYhm04LrEVbbwp63C9Jp6a54ovQQm8063AJPgJ3z
pCSNO5yswpq3v+VRFlxGFsg4Mlp36Izu1QZ4MVapyWiDxMWPtF5FoaeIPToHcej7IV6b6k6byqDx
PTKepzGzaMF4D0cLiMC2NbfV7pyGp0vztK1Atl8d53D82c+iwfwnlNc1dXvJRrytKRsvBpiazVwU
QUcToKi5Vzz7BhAvnkGXi3WExeQ8GvOlh5yMghYAfYYwkFHbn0dC9eBr7tLDsWBHMZAKSTHnhfMQ
OiLv9cL4lqd8hqKcyPBMTBpEPQAKZDTiqpeB27fYgTEgk76KkU2vb5+Tr3+JGRtdcgbElhCC4jWE
YBv3NEQFBxn2ovcaOKwbYWXgIoZUlUnwzYsZFaX9M0iyFBiMqgnVy4xihTWnSYO4rp+OBbZkwSLJ
5V98gpMV2TvEgB7h72PJCHMTT3xnQ6VCpWHqKDBSsHI/4cJpRwnUTO6BuMwrbjNqNVUqSAeS6KGK
MqrTDSeKqpgPYiAuEqVFG7Q5mwPzm2tEYzMC1kC9z0UFFKTPjtFSEET6hpbbgntEyOn5oZdAtOdp
uF3MMeZgSBnti5owbk/ZfBHQ8E3+LTOcI8EhePLk3S3Fso5UTZbePDBeS31y0YdcDldzZYztk2PK
Av9bQtCAZ95wEhdjcV+S6Yo7SKisut6GyrZj97D24qGhvnF1UNX/63rubPqUQCDRh3RbxLLLVhtl
tmVJhZZITw48Rz+IhMAnGh7WEqE1sW7J2Xs7AzRfD8Y639zooLsozW85FjWMCSrKW5MoYFgtW95O
22/dpQAEzitydUUjtDL6FN3xMjdi/kmh//4nu+Bx0mXck+DOzcb+SF6aSqrOtAv+58qoiZcIfBHy
fmxCGHXSMemb7v0EINwfwxv0Y/CRituMotyDZl1P6xyK+ii8ApyfC1i1r/37RxGpTC8T5SkAG7vM
ZbR8fnF+SCL8ew7RD4T4kA+/l5U2+zLZFTwp4WOKZ9l6cNweLPBloTDPGmp7RymNvvSKeWvs7r1O
PRZ1co4cUo9U+Jw7dllfenIn998XEwYd/xQ253QnRJHcq2+d4FG4/kw0gAABBg3QxVk3puDem291
3GDERpscqXIE/ZtvYWHhZfoIOopYcZLrwx0uuGEwW5axiz73ur8A7cWdgQJZKbQkdPe7jDT1txTx
4bpuNsiSkouQdEJb5VmNKQly3MYMA1sxYKoE+XhyMCL/NXIFfEzy4AH5PwHExa7j9X0GN2+yfJm6
qC8aab0YgVa21ZcObYGeuptran+YY4LyRYVdZ1Fl3uMYEW6JQaMPdmc2LC9o3BVElGZsgUfeT6K5
YW4X09aU72hEg42BNzFD7rh902E+kDnw93W1n1cEw7kgoRUyP2r6jqTVT00W98hKxPlTiAJ5SVax
RKHrqzFNfXsDvutSVERS15jamjUtrM3G8oQRdOlscQZJEmWWQt/1mldRmF9z/9EEXJrHqnEBQtKY
RJJOPUIc2KUV+igTA7oLWL+vOD3DR5dNcgmcxejejC1qTwl0GyNvf96nilUIe+f9pC7qneWqlPDm
E0+L9M+31vYwzupS++S4tWmPKP1hRkDmTcXNo16cUGPc29UV3JDWL7IGSYvBzrIJ6c/x0Cs/mJvG
nKlzGaGBt3F6UyHc6P3xXDPpSz+n/Z2AUe47NMeQby9XFWLqpxr7oSTYu5oGbGugHw5cF9uAolxj
pOEnsBrIfd7ITbjG0TkGsOQ/6oJeNimE3b+nCXaxETLzW1F1cWYWdJ68rMr1yBrbwON+J7RuCKrL
JQJm9tXKq1yKZWoJovT64wA9kdP0sRII9YlfIsHUaP8In3wBMWhuVQoD+0N9uZRW1xoFqAF8UmTe
1U+6w2P6zLIuR6dEKnTg5tirYh3yPwFeriwoZn9ovex8kexgjT4Civc9RBxRtkL0VQZShNA5kRF4
i9Op1O49RQhNU8TCTNFzyNOQyAvGTodwVihAIyGDJ11ffAqPlk2EexQym53RtUJ+DNc5isIfM3PK
8H/pOSqMQnqvzPKumNbAs1JQ47DIxkskPFYp72ukWSgG/D+gOxe0tHm3ccC2MQ2esCtId+4ZqnRu
vw3waXTtyJF4Au+SExz5bZ3xHBLNtyBw6dG9Awg88ajM2OacloQkSMlot+GYHEYDlAw1Cly0/4qO
jnlT69mHr85HJn2XkzfYPd/ot6teBFo9CIfiZzgUul1bWOmATdUPIihduq7C/shrxvuDQ50yJfVj
ZK7QpvktpCeN986vfAZliErbhCagsKzpYHS9PbqJi5b2ZMgzobHvvXb7i+5WnJDgvTVa+iMnZnFq
A+K3VUBj8GBZG/H8M4RCQmcSCCKLJbecsrpqtpC1oArhM3f/xC8WBNeV6/oxq3/aL1dAoQWmbgxH
/vsk2bBnqNgYjxAjMMHykEN4SVFA6WOyLyagmcubkxc/X1EKN8qd0QnX826+l68pE5sYXvy5rqNt
pdXYopigpzMW8H7/k+9KEDrG4MOsWRf9ZrKjsrtxie2cUvywEbD32Ch0OOdZoubNqE4hqPDnfGA/
H81vcZSGk/QyLxUxkaBtKQnogY3XmK+vHA8E1BJxd50N90/qtZQfrBKjDZvIOV2WCrwWCs/QIX9X
YEhS9Rg3CtyJZrisHy5xdqhgWufGeUOVkLphzGEjfD9Ny4hRyAPqVGbec1+FqDuvBSrc0tfCIYlv
jLduuetecDcAkCKE2xYZ+8LekUWv61MZ8R3tvdpBumcdl6+2InrDJcj5yQuRgwYvwMQfKO8gs83l
g6bT1Tn+lT4Bl1JjH9zOX3YUiqlaS1WZYikNLT6G8Pa6Aizm2MdeYXplDR8SfguzPvljhEQjQ693
2FyxvHQt8Qh9xoOZkPJhXQ1fjrqLNm84ZFsuMpDMr2MHq0dYCJvCe3cAp/QWE/flI3fgQj8Feu4M
BY5r2huPf9qgi7a7Ukjfk4MRJMqG+3OIOeML+xXvWd67eSE99E4zco3HDexJ8PcD9LhaJKdpjFnS
bxQCOdqygFbrT84iJaP76swNrqXLOjoCUMEGHsljVhUqJu98EA6eimzUPuwiaeXIblCGnRoo6gUj
yC6/kI0dK8t+cuwVbXciU57b+s1iZygzA3uBoFf0ufhCW1LY4SmGozIyJQ65h0jrSceBLQN8y02N
uGAYrxbjcR+2w1M9hK2TNDcsVa7Dz4bpKQKf5hSlY6p28vYwVcJbGme+UYQbj5VNTQAuKE2isvLu
oThVIfapNwykELTW+AjEhqcNOgtpmqosn4UBqpmq/8TbVF4hcctKsgc4Kx0fiYZ6hC2h+c3ASbBj
5XT0XBla4FLPOT+VCtjNxOZgaoRdlIN4nyOa95IiyZJnSmkF0L9lYF0E8t+EL3SCBz7pQvOCVwGB
TZscWxR8T7FRX5wDLB7GxkQEMJIgFs49UszTrdRqJJEDRMy9/U8rZ1zrNWVasDwqQeNKJl/H3+tU
5St66LQS0l4iaHjpy2pR0Yrn4gIYRpkbbX43bIpejn+ojvE9nfugwYgie0L0BNYdATMn00W/6EXN
Rkhd8o23WPTXSd7SVX18/JuN6YbOuQ1JFvzPG0UCjozrJsskgbBSpt2IZCmxV+vYWCwfkREwqhWs
lc/Yd8mf4h8uywZnoyJGFkxMZcJ3GWP6W48FProAB3Al33ow/Tm9sExdy25a/7D0nE0lfMJhSDat
lbBWtUk4ZFgxtWKWY8yLCAvgYTNnRmvPJoyJhgyhOBXkYXFlDmasshHsc+wypYHTspT1CS6YPnLY
bRFC7MBSwU8SPN/xIB64RIZivKy1hyIL8cpuH+mDASAOM5DOVXqrwYKZYaJllEdLRT5aAw4bvoaY
EOXgIsTUpLaOmfxSQRXUDni+bJP/bEqKi1+HarSQz7LTqmzNpxxXqLurrlM1tA+j048+Eyj2h8Wx
EojAKpk2S6zEp4wn0e7fyFg6pGX/SBZfbgS/N+Ix5e3HifOOqY9KlfLlGvR43Ew+Jk/4IuXRU6Fv
s1mWk+VYSg3vlIudxgHxVsrWZyRY5w/rx9tHKdKCBC6YrzsZKzQJm5Yaz6ou3Iy0nAH2tLi2dkZc
HBk0Ee38pvxlVu9N22MvyzN3sP/QBeuOLPljACGwZ8UwhuiffrkABZW2K2trdyDEKea7/94L59du
gdgrEtVSk0UTk/zlvwO2G7E1ReMYqFoH7Gg5uiklNKVlOsWKCFg9idLnsaQf0S8/WBoNhGrXGU4o
VC6kRk7qDQzEk+ZL1ISLawbV1cQlIrIaatR5LtbRsk9WIpMw6pysDQULp0QSOwHYoaDOUFo5H1U3
f779sCfgxtMUHyWsxrP1h/MUcAVm7V9zpNxGeu3PzDrmrkrOPRKx8YLVFawo5aVvDNvm3a/bXTT2
TUVjLGwufL9kGFV0F5UA3p0EqCbS74mTI8+G2JA6g77bhU7JHIRwma23P3iW9HdCdQVMNQiakiTp
Khvizgu+nd31NgIDe0h9uXTVxGoScI4B8iDVxV6D5DkhhnBlIFdnIlFJ2fGy/K0lhuWDXvTGSBtz
vPT/REFr3z0QHokbtZZoDt7BlicxrxeB81CcIVRhi9W/IG4ltHPaoHjfboAxfE1Eog6Nk7sW/KIB
x/q5OYTJ5c9eiI8hN8i5fOHf3cPQKqyErsfwMPewgFxOASFf3dc1i80nH+bjcUELAalo3y02abwg
L4hdEKAb9917v6hf1u6ZeAPYS8x1pgVlLNgJgl/otu8ZQipyksg9vXOts67tjf2PLo/3YyYd2yxW
9k1Bmln5UVET71Je6FbQlXLFTPrVW73uj06rDSNo6cA0WSFtIF8jDCqM7rTRc+MFVkeqkk37IgKy
v8edNXbgHYEvn3Wz4ipgev3Hmz+GGvaugaUrBMu+JcOBlLkP9aaNtDP4OplLVBimtQl+xuJGmzTc
q2Y/2vN2wWWM1TvIRYr/RmjVts0D5WNisSZTP2wgAMCPASLD/wGbPe9bHfMiHvrQ8+0apVmFKLOV
hF1YJASWTJf2hNpqWVl4eoLBrZu57iFb8V4Fbzle4FUU58N2PJw3cs2rhIo7l1Bz377cSuzQ3D/o
LXCclvwA7hcAL0X+gdZ2VUF4uyInbsyzn0bel0oDzp0bKXpohB+9Jw6O4Y+QgMXvZxgek3PUMsIH
WQ1bdVpFFvjFAtNXTTjd+CWkyJaeVqhjryVqSYRCp/TcavEGwcSVuutgWir8xguqEVqmSGoXZyrV
7Kbs/zSVrgIG7Edyd3IxHBDIFQaQM3ylez3RcDeLGUDltDm8x5ej9WyBbG7EKR9567MQdbY4AmQk
M7TVMQJF0OPGyXliUMmmzJ4MKMHZPWEOil7uyIbHurzzfJPBkkntJiW8hZBmxyU0PXJAJNGADP6d
Eu6FmS5cuNEdcO/SdAGpKMjdzCyeZQIWkt63iUvQY5W5Icko65CUSZ9M5ysgXHN/1bz9W/mR19zT
aZmxZvcpPAs4ZRuICtsCMxZv6fzRmSqqdqzY1qdn+qkC5psi8ZcHpTkk3p9PD+kswLnJlw19jtFB
dqk4IJ/dCqqvyh6Ek3vg2rs0t7zxnR8Kl3RAsggzZ+A/xmWPEWqyWeXzTdxq2QS+Fz6X3pWjVNCi
FtF4zj/gFB5ZGwtB1/fUabbhbw6B5J5Wsr6P/aZhBYHigAqeLScJKSlLhR2UQCgDrz9SQOoVFEfD
LMsYFX11RH0rN5avknGQRcgdIZE8ATMEuLUj0NHDhHlwd7MPDOEgPcmSksIKs5efd3kRMT2qX/rD
+XQ1xIueSjXI51O1AP3oAICzP0o9Mb9JC+0SNPxxuWFKthC+NUKWNhtQNdYnFk7fAiLR/Tipu6s0
6Ga2gdpxYvluozo9CgprQpCi5+mZ12rjOwXJzqdGtEY5VmGfNdpqHoOEt/MNM1fGzNiSKXJHQebD
qe+6VxBJfOpXXsljJo3fnlDCdc8WwVbSVg1DEGqxz2VQ5xuxmMaMtZzPzxAUxgezTpYCZEzg4ubi
DWj+920NsbgzHtybZeNuCeP6EUyDkgWCmVa2UIHaOm9Vk+y9MP2OZ5cXdyuHfug3XK+NqzbmxoYL
vlH0z4zeigpCzlyR156KFahoIaabxxsI9gDABGUi5EesiE+uwn9bhEHCphdvQio7YpOiwc6op3MS
F1hJtx9xELkuUvzqPMjm+DLM6ITc8mpbuzAe/d1jJfSJ6h2D4eS1wo+rxbHpOXd+TgNyoaUzQ0If
xD/WfUSoSR1+etYTxPFnlCj1Y2eu/P9mQJQdYrMnPYPdfr6dqlQiN1CTZ4xorh7lRqCQEKwGpun2
GgXBgRK+LS9lDp+GDNwzw758w31lHbgU6PGaNcmnMIznZbXmo7HxuKKcWtqcPEOf3Jn5KMTfT4S0
Nm+OO1HFjPkAfiERvKuEq/U5CuFGUkYUXVtdj4ou/91PMHMBebC7cJ4tI3Ocbsn5wsOoODIYCEnW
DDbOerWmiY3Nu2su5B9hrvQ0vFoqKCksyTmHysbrAaJqHpjiy0pq5WRmOqZGq4At935gkYlA19xh
UVi2uMp9FlNh9KWlej26NVQtdP24wN2xD4AZAa+5zfaj4xd1lD7k40PtOubU1yhLdOofhlSgJ+cG
L4L0QaVege7OVZdzQJV0EEhfzNa8iP1Bvi+FfrJ/xBPQQtK04ltGH+qTdTcPKqVxqYnXete65J4L
ncWNqn3QJ2a+2XX2LgKOzQZBSxTGzUtczqkxnMKcGnvhgr3Tvf9w1EUijHx5A2fPOa+x53R0td/b
a86w3Gw98aDR/uxVFJh3Ckme9ndKtV3BbleG/udKg/X9z8IO0iHHKD6rnVjwmwPHwiXWbbIm+OH6
QixXXAReDMYgWoZY6YqLCPDAnF6+py2tXvmLAwUDIHxanjpu1deGxEgWUvOOQgrQf20EYKp5Q89O
KZVMSpBZxhLhyGa8STAy2yLCzeNOweOEr9VOP8BDOAMjwrxYwx6U/BgUmTMyBFZRiCRJdnGizPNC
hqzd17nAYp8R59Tan6WLqM0iCN/gvZCgERZX8f20eACIjUEaxhdwM5nD9aWB+mtdrP0VEaLZFby/
TP7bfrncQvCEq0cYEjXVp1giq5camW9Hg2ut0STapefitjhSJh/DPEqJ0V0uckt1wTWJmn1RfDTo
Qs/v+YsWywzSdg9LetrWU0jLVNhUMWjrsaPZS1xNxY4NN20SmUJ8klpbjeZqGcjZ5yd7zGM19iY9
vem854yw2OsyOHOG/7XMI0QS/66sYJGe2RfkNXc0fT4gv5hM40tUYrv49yatWi0y2cOKMTh47ZyX
tSj/V1bFxpW1prvB1uIf527Ba3zbpV5favrjuRYgnUeuj/FTSF7zZjNnYk3o4gI0psipHjegqaJm
xJiHuLTlvVrWhcjH25+oq6Cg61yu1qMZDyaZ6Z+X+QhA2/CT1W5PuTqmqOULpUsL01nE+g84GAeG
tS9mYvMFfKf1qwS2ytbkkxt2rLsnUjRftJwSZMUfGDJ0tkcD+XpILqt9IDUwSRSzafxiuQI33pRk
8DqSD/hAuEWCW6ji36aGflH7icFw/QMcoCbbbw8WSbX7I/VEk7H3TxqV42cPJVpHyBW3w7N+NTxc
QMwbGowQCoq9xBLckHFnBJ8h2gF5ONTGM6/HnvohujkY9gHbcGHEqoYRKrmDLXvfh/QWVLe4Oe8l
6twl5GsK/mzFWjEoVnBQ5cPSK2DJJtuHa933E3Fg/dhqjDvPVf+I2PC3hrvjhuBshq97paP7q5IF
cs0ypkTUW2ABKZYLlXkkZD0lLRrqJbJvCCPUJKEFYgXt+zJo9+ru2TFllWC7SJKa2VkdKh26CxH0
WGOViQ9yKAKF9FZ0aDFe/yCgB+MJ1maFLYrbymwJJmumX7A/n+f4Y4BvLC92gl17bjafJQu8z1r+
U6BlM4c6/sOD4shWzITzvEukTIRExvfPCpgV4yLg4m2gl1cZXLxLrYr9lxYpopqDOK/YSJc1INKE
8E1Lme/F7ahAspPEkjapqIkDOScm0L+GzwWwxFpXT7Wuijbuj79fl88QRj1KX/eiGW9M5x+sREV8
Cwz80cqRJoW3kw8lF65rqPFKB8iDSZ+AFxJN7N0/AbhjrNxMJxKyBZRND6elm+Nx0/xBb+QeAoEX
8rG+7HbWEZ4thQuglnd7M470DjiGZUTFQ39pKWSz8FPDU2MQ5JBOzOF8+Vwhy/LudQpPv3c/siWj
Jo6VLKY9kvKkEDwRmlrFiEFLc2ZXB80DnNngLS8ZeCCEhkp6LJNahDRUcPLOLL1Ixz+/ek5jTNow
SXM+f2NqsAlN9M1vbINR0uncWy1hTTHxwAuGR3f6kg++N+2Ny7nDltKa7+RcA0nwWT/dWQRR3TEg
kbTYvZTTmEsaPygFlIvIgbfOQQfkXr28uwosZEJIYmRgzrGZFz2ijA5FiN8YESFhcbm8ml/JlQFN
1pMngA769MMPCMLgXPnjK0Byc1HT7Qy9rfTejTkGtUQx3bdzVJ1KNUyqZ9NRUWgtrYlVPfAcxVhi
Wb0eYaq66hv26SIJJLFGaS1Df1Mx70t9CNkIxg8eiHssBkxDwBZfl+vmYJdixhRPLYdKcNIxOUsF
UFcxE0uypBTzZSBPA7oh8iKMXOcMFfr285+MeVQYwEf/D0xd5TV2DGR+XjcfEXVjB+v2GiCJ80Y6
MYx5v45Lazx2w5bAqTVPKlUj4224TEiHul0G6cUVf5+azzDINQEh+Imv3QHN8hwEYpKN0TChzqFl
D0AZj/VJWqLuwVUqJkDcLKf2vFLyAepY/OqU2gpIBEka9y64WoNYYNd2ZWNrg4fEAj6ajVDlG5VA
UjJ1uninRy2s5uSyKUEqk5xJCjfnCIqsvr6sjNy5I8xl/G1mnDG94QR62StWdSe2cHJOp99UUuLO
SYxt4ejSu3PHZVO+tMqJHVKV2FfPk7AmedQXBhAL8a4uh10uHoI/aql+yYijM1W/zwecqtwnPGcc
XaR6XS8vZTr/eAR3sUlieFy7hF68KUnL+oq9bwijQ3hh75ShJIX7I0YxbYEkYBGkImpikAVJlcBd
63t55t6epSw+2pEntkeghN/IvKUjbWTwneeVlZI6yQxKqVP0/vIrw8KYn95KM/oOHjBPBEiNESfZ
7kESjCH8ik1r5fgH0fAkT/3wWelwnVfyYLn0vjHk4rjtpUg4iLxHo1qURtwpdlw5E2cZT8V6D2qz
SZh+XRnht1jkpzGjkZUoHySeDnsuEerDfhP1vifQe5GHBk67j2CpKTX3w2pDR8BaKCYzqJjAniVV
JD+wGn4Z2UsQqTogUiwCA+xHNr1S7iHMReYlisRBEYHTTf4Kd9B/UrbRqitcukiHxUQMseijmJBG
pzdAUKdHx9pCU2CZVoCCqAyqxRoT9vN7/Dl3qmxFRSttzhqGHsMZLK8XQi4/m6JCoduF5BZgSvv1
zDr4HTadZvGjhazJqDvx5RL0qmCGvuR7WbtDxG7FrRE7JwY7xoxy57VsOX/XrhDZ0/PJIptm2XLH
Ll8YUzFoWsZqNx0OiqyJ2A7gTyCAdZ93CTrYAlEwuFfhZEUO9/GhTUaQN+6V18iNkNmXUsHvF98G
twkZbHc18QlETIYsp8kX1A/FmuPIkoMu3cSgkO5Dc00Wa2ugx/1HJfR02lxYu7RTVsHP+tVWfAcs
IRF59G0p/YlQbpqTUHeL2hUfWXxRXxLzQAH1WT6VKS2kExpkFBv3gpnEOdOrB+Z3xXceS7J+ASsg
I3Uia8LmCtobNL05X9uFDlE+12xk8wsyuWSMhyHnWLNPp5QyRysPeD26TI5S7Yp16SusqfDaqT38
NtuykUBNuw0ARr3EsIsw6Zvw2notg/ElKVU7wIwRGPwHB8ghfuFdEyXozN1BAs6reOyzpI0817HX
cA0V1AzB7PbLqB/nGqdDAC21CqESRk4FejnQSW8XqvhszNl8AYo1Ymsqz+dtPdT6nVgw38M8b1xq
0ic5fkhHn3Af+wHROkCELWQlGfBDzDgR26tEHUjwAfo0sjtmMnIis8Gn66C9qaBw2ytLqqk+WES/
LrNBG7Hu2XhhHSeme02ijuMEMoK1NpdYuLBJk/hxWpZRAsoeCKRaR0uNJW5yIZkK0ICDZHP6Cohp
qS4AbMgjXm5Qfafbezz4UtI3bY4TD3X6VM8H3wQ8RcBKcu/gjyh9KFFLDRcKKn/Han/xkwYzMIbz
mYA6o6b2WmDXYCrDtBnJfpLZ2M4LO3kv1yQo2srDZkQ8CPnQFzLO/RyRkd0MK3aVJyMpFDChRHD0
rAHyaxfCREWu8EDTTN2njhiVlAxpcd8/sGG2aUDp9n5Nk/hzZuRzM3KxTfCGLykRvii/YRjHpmWo
9tsz8jkJwTIbSBsHlsz57Pw45SM9FKYrBtA4KIgbFdmWvI0frIjS1sFpWdoSm6ewLanM2eS6D2AI
6O7JgsOz/EcT7g9J2aV2M87GOtesw/x09Sd4Y27CVxwAEd/p1vJSmLSnksg5bJnX0+b3JI4wcUhV
Tqv5dqwovOKM0OWY10SBi3fbcnhB38l6M+FouCXPcQoIkT2Fpmrx2TfBVNB7BBhM3R+ka9fx6hiO
z3TFuGcP20pT7EwMPQQLBleqxKrrPcZ6nusUDeuohi0iAkGfHlAerm6GoC32tpOxFytaItR+LFHQ
qbbEOvl9ChEg3S488Nd0u4PZWbzMD+V8LmktDgpZ2BPQ5vUKIIV8XmUW2nn7mla6RgzkdxLj+bnF
OYkcufh4NuUP2QI299SWWMzISoV/vZI2VakePthR8dDoyopr0vIu1CT9aEqO3iHcJ7tYxIS8SOFz
AF4Z1YrFQWcKstWfYuXpCsVPRgHkQV8WBRCsoslS7h0MqFmdCN6QzYX2zf25V6n9e8ciIV+/gzYA
4JFhfKw/JuQeljiYznzr88F7/6oTikQVPv9NbkNU/LoCp+XJhRcXAwDx4NFrtOo5R/8sterulGj8
p/T07CZiD0iiXFGkdaXlmobfjmegvBf6Yah9I3Mgwdn3zp8Cg8SExE8ZscEQAlZeineOUmz3AeWH
GbAgCTHhayHqSAxJKePGghkx6wwAPZ2e695xpQCFpQgRV8xyCS40pgwi4Fb+iBGVh2CEY0vEsTeS
IehemJML7IFC9+kJbj0yvQDUFi9xhBooDFKI9E1CIaUgUOb7/+A8R95lu6yKBS9FfvcYGFW38bBT
mj0g3boKJN+DRctj1tbOmhLDTJLzjcSRMDSzVwHLfXblnFm9iJgEeRZg2HEmZ2KT0dzgrVd4dayC
j2oiiZWEy7TVsHggKc22qEnt+8U923Xd/z8Ea4O6VlWxF8aSuTS7FN4VK7Jjd4Oyi/OMEfF949hD
MNvs5hnQb+BMlL11RkZQVgI9vEvbESnCfAcLZpW98+sXOKaftAXJDgMIn+6VCXjsT/nv8/iQcdtk
mfqUT+NkpeGxaGcFzBeIc4tEiqx783WpTmkQqTPP7b5y1NKbe3nXEz/9cSGENTiTJnCgO4zFd5IO
8adhCFu1Sy8VeLjLuFXrp+QsJBwPLHr9fXgJ9+FccVJB9x/3KOHo58BZgv1JtU9NKLnzgn7eOn7z
Y8gsDE6UvoJCwO/5tPqcDvA9axfFXRZaqlOGGFaqKuyIiTIYZVPSD402ctZvEaQ22QDVT+Ao7Wao
h8bAtMb/u9ddT9JI4nR23GrsV7n4o5rZn/NrgRfefbByzdtLB4UCz8EQVC5kdD3KzMG8dXoQ79NW
PGn8pC76s1aTT9oOZwbxyoqlcqMisgjur41SaqwcoBhIxSGNk/3v0k1hcqaE36mWo3UdYG8Ambwj
M9x3msVhveu3yplcqr4MBSQ/YJgWEskO6I7F9V9nTljT54sK8Z8v3+ckh/t5Wk2XtBg80C6fl4AA
jZ771KX38knAqEE5Ibl8h1xMbSF+11KDdqk7P/wNbK+u2lMd4A/4lIf8gs/WNrG2qwJQyxIbYBag
IIgDj3Z8g10Mq0loVC5lwBh9VKwMI8v6Qv1wO4T7fQB1bo0Ncb7SgIfiKwoLavaj5zbb8PCxGrh7
mwBxONiNoBJggaCTyWY2vyem8FO8HjRmhpCNXyptSk1YAVpBUNQwP7CWvAd0vyhV7KB/ejsTOM2J
sR+oIlGqonOhHpjy1VnSWfhs/gKhtmO66w62gR9zqd3N3N1316eVkqvh9jgbTR0KJeHvH9ku2Abx
gU3r0lmniCRnlNl1+ETPsecb9hOrlsny2+RpuUpMRlgCM6hlhbZmTr3nrloCub2On/NcduPl8hIk
M4rUA6RAKK2T1Yzmc+LTWehBK1jvjeHqtTt2IxZK4Xx7S/8wPdrzYS8tWqAscmPeK/UtepXqpsVU
133DZ7mVURkyvzLSgEBtQLCmh1hEddDVrhTgLGr+6aAJN27xEkSwSpExfDn0FV+6sTayqPLCdW+O
csyzNyje+hF5V9H0FCIH0Fn8mAtIhbjR3644Ekj5f6YyPTF9veZCMGN/Xu+plfWAEa1GTo4N3/lf
Prf0JzUUGkRhV0VUpkySISr3fkGPfCvIJIDwv706A5pz5D98mX+P03ARSAKN68M3u8/qD7xSxvGj
dQmD9fffJ9wNx6illax5yvNiteWXjzvkGZnOPcptkudCndHOoU8hiURIXGEpPuMTHtXpzP4cWF01
5UrlA89GZboaFnlKug+moz7XCf1BakArhIlHo7XuFWtai/7IIM24cUpmOV4ql2vR+WTHVkFi2myx
obN8rnaphYwNT8u4O/0dV3Zml3EpmrgzihE8kY7VJ/c8ZJpD8MJlGN1/cqUfAZDia8OivhHofKBT
0b8Vgud4TXS2MY9tBAKPJaSBvyk7/Jsfo716MbDSSSemJthqbR0L2+lOpsIhA3e2vPBtdhN6uyrK
HDlgPBnyUFCDlV4SuM9Hf1qyrtXEoT9eFS1oMsven5qXCBf1/Jer564xe+cmRk6fr463ZcrIlwtx
0sg9URN2qxtow1b9sEJPtvSV0XFn7Z4S3qsuO9jrvVgIpFuDLzy6hZnSPBMaP7DDisAuTpC6UmOL
dOipxAeFtSsRtPPo3O45Nd15kWzrzjAi5Y3w/RISb0ytXqm6aRryum6hCoRCquOCy+lq4i6SXgdA
8/TYtEVmaF74Bu6oKbPlRdpoQ67R3f335BSuNrsltnGb4d3Rdqw+WmGTWesU2641+0yC9nC1Gi8+
uEsCHCgwGBMKZseyBWbg+7DwDm/TGJV901GW+AVvza/0l7cEo+R+jeGTYv57sETeQydOSBsfrmL+
mrRYB+uGzyAMDHqMIfx1xL9azv1OppCqruixtRoB6XD2MVbbZvA75cDheYPucfblLbZgSpv0lVxo
XFT09LnhGd5JWVF/5mlg6jTWuLd5/WYCOFHvFmsg7/L/mc9sa7Glh8No4Am3ivfbrJSb9jTX7q8o
j2pFDrvBuqgtVdU3nZHwnyQdHZoZeHc4/YMNLWtxXWlVPwJ5X1DlmmzYt2QSk+qLxRbuZc7hxB8n
g7L8j+RhsjRvstq5gmJMA98muW1P4CfOEm5xu8WK7PtSxZ4vqSuj+hA6kLEAhkkh1k/2XSaAi1Ch
UqwCSN2kFL32HQXMs3A2omLVMPwiZGEiFzv29gZzs7iex43J0rGH26QRGKlIN5k2dQ9WvCVqjGoL
33yr2HVYizMCYVnQcfm0d8WZKiV2YosSnW39GMHmevqpX/zXMkIaP1igc4K7CVGStVi0mDAst55Q
8Sh4Tp2NVHpwDOX6DNoCeLxJB7H2h8VDex9+xlp6TMMlNLLiq1sfpkLsS1zek0DqPyXahdRFF5wC
x++8MxMJKJPyg+Vvw+MfBacmUNxfZFH9MHLbmkzDA3EGMIYRbRpusKcY2eWbViAHIRr8tXeTb7V6
wP1umhi/fGCaAeOx2vk2IL7bVpZKyXTgHrkvBVAuANyHtjECWBFYYPdTRkXa61dxV8e8+2EO4GML
Eixx91gNGYx/gyrZLJVfI6CGAvqwB6lYNrf+2RmH71kqM4gMdRHlTV0EISv1ehcwfULKzUVl4bkl
OPv60iTllVJbgMPveNBjJT4EJRtovWDuj73kOQtbx5L/RgI6k0d7DyixzoC3nh2/WJhAB9J3tpSN
nz8JEfBKmEGh5+7KvMnyCQO8klWhaHEVYWertxA7ZrOhNMFPfPIzKf0do9FoDVKcfRYCAJ9DxOyS
G/hpA8wFHNO38BJb+HrvJz9YxfP/SJb0vkrbfXjefIpd1Twguku2F5LndzuKEVjEIH1mPYbdJVlb
iD9T45Uj3E0Cmx/pAV9GOLzhGM6w7DoMtATdbMGheuz6F260zCVffnwsvv7YAo9SnfUv1ENmUR7M
uLpiWdZ39GaWT3yxB2yew0QWsCnsOPgQUL5NwtWkRNZGD20a7em2+UD7mLmRwXwBAAF5K2CMp/oY
zlv/GdYx6PikidI/VVZslHQxVJA6kM5a+AzZotxftNn/hzTYC5u4Mk4gH1qssInp3Vn+KReK7N0G
A+RBrAT3guaJfbzEB69qr2HCKEU5+6CkQbu4Hb6rJ4EX43Q1ciCy/n4U0qqUsFCIuHo2tyfICSi6
lQCEcNT/nGHf0ee2v4q+z1K1oDMXUh+ZSxHk3LLtJ3iEs7mH6t90rSomtslpgyHqh3/spzC3BMpy
JZxosKuw9UeF1JWeMkXF3KrslvijBd3TqyJEiphRA17XQF/vgAz4f4+65Mp6f/endiHxA+BLXQ1Z
UqpVMVs6RdQCMdv2MJzHUpT4LzxQ+FeihxVJhTB4MABtQQErjJFN5FlIFtXNCDQXV1rJRW1TDhpC
gbVAlK71ehr9ocDaAJaYKdHw8zGzW880AtxVQDr/LB2v6CKOhbsXz6V/9kvdwtNvi/WkhfgaG1uq
mIojQsSImfVAywfVN/JcYjOqVNqedqVtzX+oKWb+ZaFfNl6w53gxnIqvQSRMKNJLtCTSYkoZd2j0
/8s8DZtFL44ZjfRkYUT3UTJ2PRDWcQloJ/NUbMpvgrT5/j3rZ6QyKrNROU9mqS609bH2ZwVreA17
a2k1HgMiO0aHlyeD1nICm49+LV/zoPt7mLfQS0tP/GzKX+ESLUM+we3SuYi9ghY1B0s+7qApyH1h
rFtRitHsly8vXlPYdg4G2tih3kWVCkqLBraHpR/cA72ATwdl2Wt2wCZ7K6IN4e1YGsykHZLkC49D
MIfCIs5mI0PPT3G4QcTEb6n9OljZ/DZmeM7mtLKsbMMwe3iWcNRno4Pe+tB/ZEWHjD7ll/O/v6Dn
IXcl39/t2UNLf1ic8j9WCB4vmGV3haERINerBX68+MddEjQ727FXAc2ASYzGL0T7pC3qMzVb1MEs
i2ulIkIQyC439IjYwkrx6F46+/D81gjoWITRaXDoOMwzdJwR3DsnokGK4HAdl4s9EC+57nAhCUH8
qyvuH0NtXinDm1yTdlLbxnoXVObsnCiDyJ4OkvDNgGA6bxkiMh9kselq1A/CUUoKTfma+e+H4CQI
17Gcvvbix5Z4L0dCZs82izM9IfZ+ATzB+c5kAFvIx9bSQCUFnjxyuW26MSv/MQEQZjU3XPLRhRE7
3MUr3wnuA5m4Wmq2AzgEh9ScHx5Ixg3QlaaLYIDV85HDFcnEChWUejmYN3ojNDntof7Vi8i6eDGT
EyfXc0OMWrYINZ9ljqJgvXGsiciDjOQpW8LB7EYWMBYn1wbdtvn7u4R6VodUptC0hbB6E5F6dRRT
K5CTdY6MKo1NvCmrsgZuMON2HfKYbIFSACFw7kW2uMG252z3uG4A/osOnCqQKr+O9reR7bYKRK3w
GbLuls5xj3qS0UxGyikIPv5rdGHxTZHqWNyYhKHTp6/zUesWhpRh11h3MOKCJlSwG5EfAw6KG20F
WYhKTsj/OC5BCHrSXfQsI4fn2zUPrmBS2Svo7wzCH/VCWncAl5h+D93Xzu5aIvf50vf1kcDr2YLf
KIZyHum0fThl27K0VYa7BzCEjcJY7bqgY/YCjzzW4yIFjJeRsbSzFhSkro/BIhbvddcCpEj7SNnz
auh5AhTE6py9RyZwKllfWempiDkww0cxYiO92bXFqnaBLb8U7oAW1zf35nj7NFParSA9xh5l4G+K
cNFCAXzm8LKagbkwQtXjYQOUr5w7bVyYpjn4gaDaf3Kf+F2bubAXnWqGLIu05XJkWeMY3empJY+p
3CLFndX0hkQ2mXClASBUGvJoB17ISuan8pAA06RCoTye7jz7wo7v/6lkzjbRdgJyLqoB3TlQgaGU
rtKMJuPSL/3/1uzy96FTJ8XEo2beWIZHsgiaYSq0aclibzi5MekJkYitrEefqXMHrzXL9CV1F7bx
ziJ2gGvPCek0xt+iJwh4eFqJ6VsEdow6yVb8Xw9p6fS2+fNU6/8QOdG0JER9Er6zrDxdbLkk02iB
WGrL8dXrVOaSCxGPaFh849vyDZa8d7haC/A9s6xGvDM6GDQ5O23BmMHvL3l0yrR5M+yvRume40Ec
E+TpmTcZGrww/vw9dXbpq5m2m6EmNUOHPiDNGCeD4DPr8Q7ip8kE9tcpuvXD9P+9HCZfcb/kz/3A
6+qJS4VGQUlySzgG0jq8/2ePIQHtCgVamm7tzWOxR4VN0XfQynXGw0kksDMd8iEqVXFN2VSFfdvL
YSkfwU0+d2TTp+GOrA0oJhZtnhKCeZLEao+uM2/12R/oxAhmYyvp6N8THeqVByfFytMLLMn8hhow
k2v7UGhCo3rltmpWSemgP86BmehClSd2158r1dtNHV1DBKnKuO63jaN+Yey3nZHWGkUSO8r5ikzK
Tq3X5IZNohnMq5sf98vyYjGXiHxMcvRuQr62IwbZRAY3xi133ZODEwVtiftXllGwJwRFIANFeVPu
S0XbhMaxybDC5WQfqYZ67aQCtvGAvxVxGBty1E9MJ7gjWWFGfMbKruYeLlwJoWQkKGy+qMXCi2Ed
dO+WDFp2aTponM+1BFawIXlCRq03C1kUspuqRnmefknRAux//WRGOFbNC8COgd5kCrzcVtSxjtAx
Nw4lLWn9KCeGlXPpCJ3b8iwaJNv2DiO4KTfWej7O/Lvkq+SjDVNGhVZJGOlcuGeklkEMy/h+mZwX
kIEujGAoUT4TSkl/GRCt/QQ7fogiLmk4z1O/H3lVrsvTPfEp9EtemQZt16VlYWtOjHfgODjQFUoU
oBmEdpUnjoomC6h2ziMZuzjg0QKzxQnueNu8tiE8IhSwYfRcagYUx5cOn3R7HRbc2s4Kbb4sBbZl
fBg6Y8DacinAclPG6YHlojmaFO9hGlp56GXjeRTF//bBiYvzFDXUezTsq0wcdUbcxmzM1EBMYanQ
tmBQ4eVZbdSCF+g2XHBFnfpHHI2tZc2RNfOuBF/jvgKcfnXKk4x5vXRNUfcKkLTjlfT4ND2nypob
5Pfc94m3HPYMcwiZQhZotIADA8CjiRpd4WnwHcmMJPFfx3S485QVSIY4QiuhDeU1omlWmVdvF0If
cvTKTGXwHIXAnEU1F5+jzoHxR+RGijYf3ZUwyUgkR5VLlHkJsHPCTMWskIlbrZq1FIYQlVwOIYUe
WOsBNqL8LkaK/EwWiry0Uu81B5QxSA5spkelpscnnHlkcGEGnV79cb1zNp8vzNFQN7R+xF4n56o3
stcO+E6XokUMNcIv1RtOVJg7jwx8IPDtvoNnhzYTsZEU7TZEIaOWi+kuCRhGlVK4dPfbf2hREgDG
2WU0Q4xuRAL6CLOVn6sZud24eDg1hD0BxBRCBfzng+M1UWTsQv57iUoP3SBhuzXUK3f3sfGZ1IC/
NlndEoO6zhHB/8mt3JHoZVOHPmzVvJXOk1yR4Sare1FGCsyzSzOOUOb74hwEK2K6Cdg9RnIItmB6
7hlBZlJLNxxqVv6RafWF7bwt55NnT9qj9Y9gj+ff/15PctuiG+0UNmpaLicKpD1HMVks8R3La575
ZbK/sZvA93mQevkOKQJlQy54j6F/i0MnPtI3NavuJ0Dc0HI5qmR4Y1dWqovsaua95StXMBHCq1Ti
UHV5Enh/w8g67PyTIvO/AeHgnxKKPYdOwqxlDSs8Zw4xf0ENUsCctTApckZI6E8wD9lJjbiYw7au
ATYNnVKWXIjjLweQ7LYBV0ldLqJkima0kQO2nc0w/SwpdjPLl9JNCBXESltE6uhQijny1ApBVwPx
1wLGLsrT38vy36n0qYm8cbEjk2HH5K8PfPme4QThKojf8DMavwpJNk/d+NdT5orTW83t0g4jTMrt
a6wqIWF5S5Yk6H08/wVHV+/QBopllfVjH1/jHrlpUt29S2EtP/NOWscXduNhyyj2yPJp3x19Me7F
eBqtwMinsx1EsDSrD5fCuKjjipmH5mjdJ5oUg8n+IRX9gt/Xi1+nJJbCYrvvyMQxmF9ayX4bRpfl
Iojqo+2SgGlyzHf3SZfjc/3UDpCqCIPDpmTNlyu4fW2w/X5RKBDxu27M3z2thXldqI5kePxmoI5M
gC8NFzh6+RRa8e2UBLzd8VXdExxfSfz8Qmv+e1o8PCPmcOzT0X2+fOYAXsX+/1E2XFIquxlLefUl
a2ICgqNSJKaYKWVoSuVmEyLXimFQEMQE7YT9lIo/jJ4QkUt6uEc/i8xMHzfkBBDxRNORpIoMELu7
IDZL/Qr7a96ON05MwQJymQOvT4/BJSw8Yy5IoMlsJoAbZzXwOHfSUjymw7awlVvD4N1qiPU9WocC
NPaNhIGQjTVcJ2StDwNXCsDhCxb9gRynV6zT4ORL5a+rUUFmv1M4cBbv64IdLkvMv4rKVyb/gpCS
d47XHiYzwnMf9zTThIyy2plptKw/DtbykCI90jL15mqZks2HJNBw3hIULeUXGXaACn7GQ6fnVRWW
TIUnfhA0r7nnlARx/Pqe183HQgfSBJOwWPuf0B84i36EpKst5rmD/3BtZoDyOPuCsr5UeY1f/6qr
OIffp6D4HauCdxHFqnIgaLcPwwqTBYR2pewor/+7nYk9DN5/Kd1klfbJLwTviRYY5PzxQxGqdCKs
mK+VeIlZGIP4ItIrA4QaJOv5vwHHnBGOmeGc7TbCSG62S8iS9uQKpCwBaPugCu15vfpbZF1K+zLJ
7asBUKXWbed22HGlHtj3WVFGuP2EimuLjcsZwCJJaCfSyOavDkZ2CBqxQKxkqmhbo0jf2qeQ0DS9
1wHoctnTe1DTMOd2MXkrP86Gi9ESE3Y3sNYBJhU8tALkxbr99gNFMwkiCA8IxHXOVhslRPw3SUVu
O75rLq3Pt7R3Ee/MhNhEJCzDZRCJYx/6WU825n13m5cRELLKL/FHpI5BsPV8757W3iOya1acofjT
NT1hDjW8PXnyQD/sNOiT3J5JL/cZ3EYzmaRz5bPlMqiHXRFe+4r2kl8jgFC9XlgWiWtrjjNDmF/I
6chsEL3T7ScB1CEoxNCz7nYeYRWvcaEK8y4ukoBOCrwwn9Ekbm1rCSNjjkVK1XacKt7qGu7ccXOM
mhygWejXaOXRpCotiJQQwFqRNepXMYM0auvcAjNCKSTJ36Y1FAC5l08c0oRt6csY+XMqac/WQ2BQ
V05fk+CorGEDqDZqtj6Ut+TAZnUoEiqFFOWqiOYwdsw3bSVLHG8bp1EX2ThnXbuRtwe5SygxVooi
msVP3+UzMK73QcYIfBAVKG2bkZ9zR9UXhn1o6aLLPdBLMHM1OM2GXD/MZTCaqwuumtwiFrtQDeq1
xgtzYZXO1KNqPeiSSr4MWK1pMe8u+PfnvKxJzXIZSOovb3zmYVjbDYbdKlsv8dZdbXqkY1/dYcii
Z7qx7/94bHbzkRTspOZK4KcJTD1SoNkv2tHYjBD9ZcGEb8FilM1m+G9RQaAQmkbRqNzvqOEWS9ox
+S1ABBSCvPKsVHRuSLr3raMWFosrZmgk83wyzPwdPiusAGHhTWgUWCRePZOWRt8yZr2buSv4aqgU
N7bsYT9P6BWEXNe9WEV3gynxpj71BoZHiyj54vcp5gdHGhUDVKcE2HReorWF0WfIyydJeFXMSdQF
0vbenVP3suGjlJ4bkh3QraEPFMsDko/Ntu2EAGPfdkCw7SkdZsPhl/yyE5mGRGUcZ8A9hAMW6Iwd
ysrvkt8/GAH3RLJ4sDmu/Ran4Bh4YylM09dIZ4BD8FGlvf0d9ccBj/R6IUMAlemSFitqXhAzKF2u
dlY7tMtXoUutCzsbV140a6wWeb2SCPMMcIDh4JAqtoI57Ggb5SK3TgJGPcoJITsRFVJa/GWRjKeA
DPeAMsbEjxbsHKyPUpxm/63hDxUgsX4I37biUo6dgSy1Ry+VXjzC/w/NCxQCn6xld/euvf0Bv1zD
81Wu5xDvBzPXBbYaPHS56LNa7yrb659eEb767a+PfDMqpaaHZmtrTvVNZ5qK+UcdD6Hf0Axd2A1W
GGX4YOeWPdREGBQXx1AjSziE5gohyYiRcwLxU24UbHa9RY+7I9ovSxshZhFHuhLGZlK1W/GA8Vem
qBFeefM3iUUflGmQmvKP+W6AvBaI9KXvTwkRNIgpL5S6DQJWlNc0mpVEmkR/R+UbRNgUwYi2jMQb
4aqx7GEumkblU0GPP+g7ucbYTouPFLk73dr3oKoLoR5me3ibM+vYfhchoZatCzKTtskthF4g8RFl
hZHXqO/89HhdV1jx+YMCQs499Fok75CobrF0nOFyOANGgMb6fbTzv43oy/A8mU1Zvi52OkT69ijS
P2DHsxbjQZcxSFtXzoIZd1K24eSP9mDxc01iHrLuVPgC5TpLZ9pD2MQ6yZ7te88XgLsUC6l7epdA
aaA5jNooiHiSu0rMH6qDfVYqcE5p3uUSYugU4IN/TsbStj9Fcg8rpcwNMeZTNcqF/cCeOLHmAzRh
PVaZ7LLQh+kgce8nQjG6opIbBH3gIIu0/vaJmECG8PoBjctg/k4EEUe9O4E8S9E/mAlmkehTPxrZ
YgKkg5Pj4AClr2qiYGWOtnneOnBLugHRKihO+TN6w4u0xLM/0wZqE/LQd/sYPKD7/m077soUcmCV
FNbEcQKH0xL7tdaJAhCRNd65/DPl+Y6hBzELSaWT78C1wf54Jteue+we0BYHf5ghoiL/Fv4k+iCA
EggQaQZsL4EdjT0AFQ8Og3Nkf3T11bkblcyKPzMRuVCLn0hd6w5sRbW28dYGHliwKPK7bykUCIvv
v+EzG02DBz1ewrmEs8Ud4v7v+bf7oyItdX5aoJSNRI3bXidxxWvasYYjKVv7JVVHZphwpUTWUtjz
UmFlcF23fkI8I0GlhJ6k16sIPEKchRpKGadCksbRcBWXR9EPbQloNpkl/+pdZiKh4N7/myT0Z/YL
YLcd0Jbze6pl71jxLhdQxqfUuPUJv+bwHzt2GAEM/5G39V1vTVPMy0OAqaRE/vNJRCz8/GnL3HUV
Lc3rIpkY1XvDyEYK22ScmST/SAFO1fXUG7HwZ2miam+YkJy1G8Fdn+EeXaWolsRl7V4F3xd0YpBm
5wMrl3a9dI97aoM3rILdN4uRIPJsLr+JTAd3a5gC/AIT5cSnV6BE3KdDy/ErwBiDJqsmw/nSwdUE
ExhLkvX+tup77DJyYp1WM10d8K6EYXJfOOiCzr0Dve9k6WD3tMTzN+KLW99CEx2WMFu0bHApScC6
C2DXYHLfY/RJOZdpFyHDkjWhbYMIeHyd5WaEm7jF3iN90OMZGhoU8giwXBAqmZkAdz+cX0lCDsNn
cH4j8Bx5oom8u6uUtPYh19Sbo05BaK5ChuwSyzjXgXFjq/XVVgFnQc0pWo4NIuYZc2+ZQWIpLY/Q
AR6nEAvCZ0OZ0j0YIE2J7eE7GQRz3DgxFohLwC0wL61H/C/E4hVHIpCFqPMdIeEro2jXdyEfSWiU
RxJRxOddP1piM1AuqoLT1tV1ek1ucYbVGLLEf6nV6w/l05IlEFrXtB4fGxq1t9jV3NE0nNTSfdSZ
gMlAmhbdQ2i+N2yNUdkdfzeZfV1bwaJTnW+w0Qc1yM8ulPilcGtMGJm8CjeB5kFBeoj3tMN+LEMC
cwphXImP5GtOuagSCL6bfRFe1Cos1P2HEdZrvnrS2KuxSZvNMXL4N9c7KplmIav+7TywHP6qInWO
wYY7JAKEsPlfmgLRxTDUogN344DePtaJ1AQH9hm+swqv1wDadR5+PyGxpVpeGal2Jqhq7GGC/11i
MU0LMCCkMKfly8iKF+JQj5ARuL8KiIox2m2pXyKHbj/k78cgUDySNRnSr6eR66evVBG0pDdI3Qm3
yku+YI5eci6Kb6ZQcM2ns1G9Qlmxy6+3adNpl7KsuB3DjcMt1NjKNptpSDYEW5hua6GlwIqd60NO
vQDPLCA9ae3IYvGEN/w9N/VfTQvwbpEyNnssUVOAPbLV0hm2eZpZ/OZ4FVoVnssbHejKRidmPQdK
wrnDNZIVTr0F6lQCDmGNKuOqoegHTO5qwy2i+qlQoJtKSL5n+eLTNoQuZTLLFJfVfNLb43mLlcjj
ZSSiczfl4g8jMdKRiWSvzegU6Eyj6WuYsLkkiWw78fyLbEWldWRAxexhVOdxZ1UucIUl6emlgdLM
OxByC4saLUvsm0/bph8WzoRtZ0a4Tz1KmQba4fhrZSDN6g5wRbSrm4eFLjFvPoBSu34YnFzyCndf
p0hXXuV3izHpZCY084tEFtOHOHON8j2PJfakC1GFbbqewFRpX2eFLM5/GlKX8IgSAWlI/qOqA5pA
roaSsvxd0R0+yQYyyTjAYV4BPXbWSmj7PPwNAlGGF2fJoSvWHreNbJ+hGJTjuo/YsvjxG73qwOWE
n0mR1ZhlXLAT3VQOVA+xCB5Vyo9sYIZtWUaVyVErjvyWu4l6lsOp50N+TXWIEK4kv2jkac6YdHpw
PzWmJA/bDqc/kmrcLA+U3ako/JMHyoaGNqC+/J39Zs/N7GahbtV5p5bLbYrOwKfA2bMhTue8JNU5
3xmZXmcQUYJPr9utFB59BinmGx9by4ymm7Pe9V5T578kabm12JsdM1UFcXRiXxvju7Qs6BwY+e1U
VLem7WaOqJfaHvukSWUjmpsQIjFBlpAhuEOv/mn4I56j9KuGKBDY3fgyWrkOmWfDYmN+kaRmECzG
xMpmkl5pg6cA+NKb2FRYbFlrcgG4Pr0EjAUV415ljy/bMH+hHjuw1m7EPIe/PvvW2TVYWEkWjihN
31MzWjboQiuc7xJbQzgQd/9qurFL49INUl9AlHpwt5LCxKGWpzidDQBkjIg374SGPUv7gLFI+LR6
wIp3oSFg65WuTSlPwpK6HMAExRsna3LdeWb824HjpyCbMCVQZqCoJ94ZFl71SPppw9+rfYB9WN1H
+1HE2464LxU1yyDjnXvMpTmjxdxDc160F7x0Qqiagcu3qBAv1ZidKqaiCbDxbFhU5aOB2qfW8esF
j0VbTTA/2QSUYti/zyHpMyJEdZ2B5suBXxYI7jLguIVHLssRt6WQOIq/bSnselQv+Dc3GNbDwUUN
jtESZ+mjJGY6vwHUqlIS98JdCg5K8fF1xcq1Btw4WLB91Ns5BDiRpevL93kSok4gGdx6sD/GkDYr
8KJSclU5u9AdtmXlUiOxsvUKHtD8Quj+0JnthOcskWbWGalDJ50i+m1q4EIcgUJ4MThtUMaux8zU
r2U5gc7r0ucBSFyHzskYtiewJA5ZB0D2DDLqEjlHcZu5/CbcCiwSh0quHDvHDEplpA26KKQClD8Q
wDQbK74DBWnHO9zI0yQEEeaxLWcHROcSYwe+eXzTrlkQUhFXRp3rt5jFGh75xU9Cyw9vO1AC85WB
Y5AYpwaNwj5Iln/v8lY7y/42tagywyr8iHSdhXh1bJJ/ZrX+VGxQcD4MEBj3sNOdAPkk9LeUg4V0
q7SCvLkZwU4+ydPsQbEZjwaJa2yrtSHL2agB6hFA5+An2JMMcB+T+H0QrOAr7YRxFhugLX77O1kT
queYgYxMWBtKLg8Lk3LjT8D2877jVe1n+iPJGBCFKSOA7EHKd1LX4ZtnwliczQRanPldWxVTQUs6
e2cyvTFCUPU/enuUd1jEj4HEZ+wpYDyYKbua2dYf06NhZdrmhhnQdJFRA1S7vstCjgaJdyzmvbyf
xoMz+iWL5wgMlujiVodRn+cny5GONv5MLBlPpN7pVevpb1hdTh4z2BsiLw+ZsW55y70CasNDmxyj
ycK1vU1F14VTiR1Wo/tXodipQjiGJCGJGS0ktDXfTyWxksdhO50HTASVpMDhleqYKerFdg7/H+hd
Xa3+aMBU6jZiQVEZlAJiPtmj5nccg/Y63RnktHINjvLZZH1ktwtnHuEddcDLa80/+lC6kvK7i7pr
3DmP2LituGkrtyDrtXHuddt6p0YvYbdhYSGj2wFJX4p5cIZseNn2BHvXZzfSO6I5TdmIcLVe0Jac
fNDrRakyHCoQHxScwh4M3BIdEJJB4Igi70ELVbDjjazKFvsSsbibMsAtrPGXuRXzCs6Mgnvqgi5q
16U01kE3XlqOKhlgTcNvnQ4ZTzA45cQDhCCxO5rgSJaKryBuSnukbPYLtykU5XFmoYs/8DaGHFcA
X1+a1upVPppp709ItH635BRnIt6rBqcWYLBakHlagK+wPoa3VILAntP+NXi8mMntH9/vmNUrhYic
niF01MoPlc85KT2KVmhiEghqd8xhXu3Q5OFDzSJc9+W0uWdKsTSaqn9EGyCuaEala1aVLR20dfkh
qdfL2fUNgQ7FU3GyRCXHb5a0KfEH+CMO+Lpu1qCAljgBhKlUBJu/cK5U5K6li2YV/lFwwX/y3VqS
p2NqaL9oljE5NbzPzyNNy2dr6RzqJh9lkxKytp4VACif7ryJ1c6KctmWbaVrZ5EnqKf1kUKfTgx8
Pj33Yd+A1hc/IJj3Gddw3yrIOVYW/pi22gJPNsw4eRDbrqnHe6mFB2IzjOrM9eccGr3NrHma3dBW
RCCrlP26CEnChbuUQWSA9M6astc0ghblExHLRvA/UWpkfR69AvY7smpF7FG8kJ7LkKrJoiGje+1+
cdZOeN8MmnaclWsB6QHM12cIYJxqdzoPOelR/0A9w7ocvfvd9ctWDHMJEnLgJUdPjACpLRSIa2tP
Ct9CdEwhF24jKdtWuwJ8of52eH0n3HFPQ3bs4o0IdOIRSXYCk0HFk3D/jE0ATabRf/tSEnrikzUN
UAtoFoqBaAdgYSOueUf3pANtqfBh90xCFWvIyhx2TNv+ct67iyUr1NYhZdO2EhFuxUTkStgoC6W6
//FwUt3eKwKcla7MjVvp+C0iLq1z29c/lpxXMQpY5nT6FMyFW9ap3GcYlS1+jZYV3RRK0pF3aoT6
pQmI+xsX47w8FdIaL2t7lzfYQ4aKupHNA80RguzMinb6n4jMFN2T/MndKoHeh0Ytc/WNOX0QV7/a
x/QT3CuZVcDcNZwhGR9RSgyfcYmWVihtNSheLdzh3nDaQ4htzZJxArT/z9Zg+vMwhT6PuKKsuml7
kJFbRe5rVUiKt8V9SusGRNaNzbgRCqPDGAseR9eSQsZQ75GH4yJX/O5GUaNR8iZBqhEC7Z4u5h3s
VaYKCBpWSLw92GTyhMVj07XCjiqW1oM4ZWvQUGcXDeBYqxFBRUIHTUCrcZPLTkc6LcWQiPLvoE2Y
YLrt1OS2jdsG76Hgp+3rhefFHHUeVUhOdWQE2Eba2vjYUjrPkuSMyI1iVLmN31sp/BxuYSJ8q1h8
r/7ay/rkioGPC/Qon1CIbInjN/78yEfiHJRtIqDy+bVGpT7ortmJu0j81gwTdAL82yUUScaxQLyY
HlceCMKdGvtbVzGV+JCP7mUM/CnUQYE9sTH+brLdmldb8bxZJ6DEeAc8/wBkstxozJIQe+sqM5HQ
AnysyrE152XD+NrUqebhcvOqUfI5WqcwekqwM9z0RFcZ2GRe3bvub0DdlbsTRuTtzi9pyyGWGqiy
bS43E2EHySu7Ork8qTYPTuwp0fFBBfO7TNecRnNtqWVni9CWnahTydaytDRT0bxcGyTA843jJueC
tFDmYO1WHz8XO3Iwi4Brry2Bhzo4i39kOY6XpPRtcpzcaXHQt7fNCbKDA6QcUWcIKlG2EMnNShJ9
58TmWlfTVks3gCeOXiztxRf8/l6KKEupElYLYDcxU0eRTKbqHLq/Ql9eIIIi0m4KLcmuXVplUu5p
pKSDr7BaLB0MiEFavRyGj3UsEsb8mjxI6tGDc4KRPNyU3dZN+BVKVzy9YIIrCtANMZNfW5Hi8Rmn
zlcmuOyk//t7xKpjc/Ss152ge4tvd2xOkyOTgsUkNxrslca4rlvH9SJOdiZt8MdnfNKlH/QH0jk1
SSzqGLL6z51sxvJpG2aqEYsQeSJO7PE1NFKjBTnZAyE6ExwGvW7UV7ljW4nMLJe9Fb2m+k0dj+vz
j/x1CIJhJ9q7eZBdDlY/EzH9ntsTx2siXNPPlZI1LilGtviBH+4crzCmwEqyicqDIynCwPrN6meT
/kRLk2fQc5lKFo4XDEMZOIfpXpcX3nHiUxqWNZtqqfGIHuPXuKwT9lpBo90nPehZsSVwz/eKepov
b/KLVLolr+yETXPOgMEkTw/9N4OUE0g/s1EVugIYnngzduJyPQ++7/wp5vYVhCMbg9v3CNfRCDZ3
EHnRQ7sEiKHgR4Lbffv/GeIsMditDaVUwh8fozR2QUgOh2+jNUozuvy66rT3KuOBJt1BVu/g6osp
aLvUvx94/oif5kfquLGBVJCel1hdXS8jC9ejACqejwuN3c1elu4opH2K1EIFlQfyDEASCjkjHIXJ
HZXeEK2SVQ/gayTQmgK7/Y01ZqOgdGo14K99bKJRHrTs8LFzWyMoAlvLB30cJ1wDLQzfb9hp2Us4
JnJnZN+6C/xJQu1H86eDBtCq/0nN1ry2vSDu5Gxp72z2w1cGHslaM5zhGSLCbXNX4O7X21TCthnD
oUer/7sFOQdSRuYIQLIWlmzGBlJgKGwjTK1feXWV2tJNbNd7+fSCcNnhHwfdFyiWFtXIQUBC3eni
pnPAop3WD02ShDM8GxcJHRfjBHpgX3iOuPczwvyirMAB+ukNpxZh/fXTIidvlJMnWsSj7EfU0ee1
n2Kc46EGco9qeCe+XgllUuJMlrzHx1IfGJrSCMzBueNakWFA6Upu2PAXRiL8YK/rs4VRMAneTDtp
0lppi4WxAIwYPnu9adLpWWlUYhViaVfA81C1Y8IaZa0IpOfbIbHhwSMDDpfrscUYsIX01sWO512U
LMYMrAcC7k68WzuQAVsndh0EdRHHKkgGEnkxugnM9HrbpqBPJD+0iQ/GZfLhqneGUszxna9xuhxV
K2zLAG2LXCRmIn0Z+PDk9XXOilUWsxLVhrow7RELtqCwef809LNpeU0gumsqm9IP55TD835XikY+
1MDPV6r/C+z5ORvH89FY0p5T5cEDk0W4yMXxgJ5RW6RJRvuUoKj9qAlNYFnGqO601Vkcukee+WqN
g2hYlHcnIkustmqmLhfAq6R2oLInkDsa7ZAAv8Yuv8uIxkfrjAhal3MSb/Fq6RQFSRGDBgVSRqss
JcP2fedy4Ojsbq2e20I9ur5gmRTRa54k05CyTbhOrn89sWf4LZrKgUGwotAMCMnZrRfgUNcyI+UF
Fz9FELHcfInZGnHZ51lAbqn45y/7wujm1mZCCRY6F76twyZdkAWGEomI1BnHqhjgebg9LqDMJpCs
beRZDdr2OuTlCAExtNCBLhk87CCNXBplx5zm0MH9zUGGj/mWH/Ky7RjEStDMwedDA2Fonc8/Wc3Y
PlT4GWaWRy4FYw2/ORTInDCKG+eJP3fvs6wK2vmZQp6/kXWNhb+UXxLlxRu1/33Eiqmp4CkkKiVm
HV0tye0oRa5wqcttsH0TTmdMGEvoaRhzq2mIcBsend6dXyqu3UT6AJQAT4OYBwPfdZ6/5yo/K9Ng
62AitdidnNbBgo0PHBLklHKJEayaqctC0r7z+N5A/a8XJNnG+vVPW8BA8mXVIDNsn+2Mt7IfCI4s
5zeU832SS9IDs3wdh6B+WQZD7mlZhuamKshEhQB5GINiw0WUD7Mg4UtnSfNtxu4rXx3QQMTrPG2N
UTuJ/unqVHAB1Qo2LJYcNl5ZWp7T81paYuGRGpkriPe7hPLvNtgxTjjsVRFhT+Rx+FD7K6dNIGR+
oOZ/mLuolWi5o2OstK1siERyypkob54UN2qLihBePQQl4nAaQZvbPmPAyctlxYH/m9t+ao+mif5b
5VG6gHIL9kMfgYjKmEQIkFeFggzgYJqt6pIVQplNKF2o//K+ALebx7AHOKhXwIxCOu0xvJvwD3sO
oYqHw8bv/Nk9Gp3h2ZiElJQg2p9BV7AxPRfFN0NTkCuLZRa4w3iNBwB7j8TXBIEUYhil0BTAwgJo
XTdPSUK40t8GnLx5ulegNt/gw7QzKdmLG57MDzpISaZq4Chj+zGL+BfpOhv4G5P5deIh+iRLHbQl
TMuMkAX0sn+HV9AjvV2kdcGDXqj0/00DdtKzUKLYZXjbbWTLIgIkbhYkYSeZ7wIHN9tY9tSi3Use
DPZ9L6OA/JE1FiiRh/pv8fErBUoI2evgYWoOAHdM4UQnkOrUmV8wz3tK5W3H8vBXbsSzs57Bu5L3
TcwcL8I0ULZr3ZatlpVpY5RPEgvJgjCIBxIAKtsyRMioxJ9NMINHWi3aDD9kv5JYMkpWQFkDktW9
fd8IwRJEl7wfB4kOmrVEsZ+ytgUKyd0gYTgKfLIAdPzHPEEB+OsUUweFQEL5yvy3atvO6QYEZtu+
LmAv9V97aJlfbXtDeVZKEXH6amoshmtOtBJjrBhfWiO3rY2DLKuLQ3f020Mi/ONkrNbX6IR9VdXz
HnxiX7hk5U50CWFgRVb4HUfeuHMrgTEvwGD1JntWOFZo+W7n0BAKXELAHBXQ/54qzPmZ7FoJnC0V
Ur4Ndf+eQu6OfJt4jkj3Y0fjlh9mWeRm7IVuzWhFoLbaghjm9jToRbj7/HlZooJsU1RGcYnOFqws
pwzfIdfa5BKVSysQDFWK6VAoCBmiYv5DwcyaZC4gP8YHf3vT8Ckf6Ci5Ljg5mKToVfkxT1XJQ+kR
OfdXBUdQ6P2Vy6J4qlrqyj9rydoRqYD4Q5huAeSLJOJN1L64PG9/USJZCpbYPPgzL/2NJl5Uw3nh
HiYx4KOiPAic3lYzpsusDmWdoAjOtDfX/6kJ0wUPZXCslXnubP74BF87C50K7IPRP/6bB8FEsOZ5
qtRkkKheUyuZTtjzELfbA6N9CjFufbiwOjvqUzDy58sh4w01tWfnmAA6LqMBl8fPuOnejUvtFdRV
T6LJAL2LtfUyzN7bxzlc/VtxXQKMxW3wMaC6fHmNAlfTPmD8tKBxJkr3798cNNSwxWg2tNhjDpkC
y4vOmypkfcp/Pyr+BtD2TvmmBdksz0vIV27ZMr4xIG5Nzi5KAp40w4AoDq7TZ2MSbUHfNTJTnZEH
dXJ9aJwx9QKr7p3bLiNc1/WRnOj0yB3CwCXZgmfw+JSfBb+qZM5P/8qhXopRulmulbm12QlzhlCw
WbgA3PGqip9iGLs9gY9ZvT9brnCbm2nURTjTWrxmmEYYwuPaa4VbxZmJ7Xs4iELQYifFyk+5lBZ5
W+CnNu8Q0Ed/PtVIQnmyQ/eZBl+bn0NFnUtJZhgdSz2KeA3GtrcG3gG6LzI3jyAfam7Jpoteaa7i
tUdSpihZZzpogKah5PaU+60Ch7Ha6c088oF0+/zQcKi73nmuaVvxbIKJnl2N0nmlV6ZFKYsCo0Nb
GY5gU30s3RGIf2jraSStY1wex/RGiQt04IqoBa/PJVbMqpYk2nz0V13RsuFy9C4Cd9AQw68WVYxN
Y2/N9ZoPUXVCaKC2qrgRRXluFn4lInx9lKvLvOx4fqo+RPcpyEVDbxRdSRCp6tRXGQJarlm1Eeml
3CpzXcmAuc/4aP6Aphn8vbNEdK8FG9AVS6TESQiY+RvBLgHp58SVe7kL5ugdpHZD0mC20LIXjGba
kzpW+lzkmdO7ybSQVRVR/PcfZgy6RtW709oVZBerA+SQXXx0O6YJyOTQWD7DF5n5gzH8H8UbFkKM
qKH9Q0zFN89zMAe6wZUFNxTaAk8CWub82yI4SaT0RY557GWpeAsOajh57NTjqzHcKiWDje8VbYPo
JVg06piTlhqLvjsqEE8CSNnPvOslbpKoj3KhIdZaQwDMfCgo2ih2wAohpjKHVn6yi32YauxR7lps
TmisO7W+UE3mM9na5wkQICT8hqnvwdyrkEo/4K1C+PpYmFMxw/sfNijT/4SVoUGFPWieKqmMsvea
XYCgmfaCmTTshImi44cymB2htiOJOJFH6UuVZDDg2snBVCECgGExdeSXZZdwLnhalCJEJFYb0nLE
VgdUElbLC8jp8FE3aIsOdlhTBJ2AZRNjr01SF/rfrgCxNTVXKM6vBHQmFJ2aInwgS6XhkrjScXKI
WmOAqjw20mCzxdb0GAZ9Nv2vbT2YIrLM+3aKURXkD0NCMs0ZkPKMTqi9NXNLIJctNfwZFGLyip4s
4rq79oSlYs9otbgK2YxXltMOeeSx0FcM8PuQ6E7dFYVMjKSUvefJ9bHAtFnrjjQ6t+WEt5jemJKW
Nj4ROvb6/XmHEJwYYZ5bmdsg55i6YyikuC5MADe39GwdoLNbJXpFaMAXGQBxdgjgJHSuVVMVsGHp
p6uA+Ea+FKQMYTdnbhyXzz2Zlw4wQxvpBL/focOSHEF2w+/gomMh0QneBvlzd8Cu8ms35DXaoWSY
WinQeyjQOG8w5qvVFvcPQ8CqcJSTz9UFMqnjwrATCCbNbfarlSeVr4UA0BCKkgVZVz8gDLIzbo6o
oVewrr/HjqjYzSPRYA+JIxi6WcBjZtPEC7s/joeeNHFnfHjfrPxBO0ACctSpMF/1Zoa0JfVQ8PLi
kO+zRhbUk7b2YkOv1k0Z79nUmM2mubrOgNZvZfLK+fo08qjNs2ZiYeh2jJKKgSRM2rwHfZ3nNMey
ihtcgukvgm678iGQ18nP8K5AyQ+puPvFoJ0CE4q1yjfh/1NoPvtyzuQpdLVT5Ln6jHaZAK1K0zBr
4fzBjAzVfOLRrOANJ6y/kMNbbEeCu1LN9T/Bs9myBZicOgTKweuXg1gQug9z/5VyOuCGintEE/Hm
cM/NwBI+K2NgIA/NX17k7o49bgLq2JQgKijlqCplfZwZk2JOGb1bgIikE+bbKSXE1wLE4RobaMVq
1VAzB/klG2UyqMJuZS3Lr1YDwLaGFKoYUu8iuHhx4Sx6DTKgEVtgJrDgUzYKXIvkkBogVIt2yR8/
lxCYypvDEPaODEIW3vVQKq0C0DzPKiuQ74bT/oJcY9hbVmzchJkXKaiEqrNWvAoyu0e8v5rE6TLp
dNQNGb49qmzo4i1Ood7sVOG7hRIPXjwzUtBoJutw7+WGYTAiTG4/i9sdoK1ObcH8e8EdZDG3Qzcd
W4ucPLpMidL7KJ3E272YMXHsohgpsttfjHkXAFCGHVaxa2MtlFw8RlryfzVDADPa0cN5bzQBEIIu
gxBqBo6ceFsrQioAgsAfUw5AGEvQn9E1UWs4CMV63nvrZxqQ50BjqC87/wsB2cG9Sdn42yjCQL57
ZvVTXXtKMFSFLwRzuhdSrBAhfDWWWtTaGU71qy0XX5ZdmptFUcjvVxNEity+sjlhbqTbVylynZFB
pzWpJPVPFLppstC/tp0mKoO/uZIAdJ0uE+88d06IH1UXxHl6ZbRieiAm7cL1Rp4INFRR7RUY1uqP
hs5J/7AEGisYuq/No8AZR9efpoqlAwflH6PKsxW/kKyJhqJlUwpnKBfaQqpLFIBHluiCoZEMc+yD
PwGtJREXnvJSkGcdBmhaiLIUStuFkA5Z4dmr/w43iquWN443lrb8um0FcgqOZ95U9JPUZK3JMqUJ
vM2bUKygVJUtWunAX2ODe3PvwGqzaNWDBXw+B8WO7xxsD6HQ0wcFO4qBpGdBAONqdPu919soMyCn
JQxrGXFHPRCJw2n/514Mh0rit3N0sMvCqtMUiVYEizjao7i4xRnC+UUOZED9h7QMMCLfcf4skFaF
6hjwFeWu+2uL6bjomufeYWEEAJsYr4evbn8avh/DUV1J+VRvql56O2Ola7+Tsidi/VXXlimIC9hF
xHVmMiyNfTBsDzZR9bXwyREZgoUcjTpYv8cYXLlQ9Y+AF/jgqd5cMrOi69++rEqlQ3tFD8FYvKyR
hDxafLPVfmGNMFJchcTRyli/yA0g3j8ov8WuHaSrJbzAngxR7+Y/FJIbcbOE/pmen2B07ok4Fsoz
Dq8RvAacPbCmcSXV+2q+4RxpufyGH3/28hUTp/7N9LDgdvpVSqw79WiUVoNXMZcexHwxD0IhwUmS
88nIDWbNMhy32nUgHl5jsBjmpQMV+0jVwCHwKk4TPAJ0t99jvpGHTDATof1bS/plIgE3D0usuxH4
BRPZh1KPzInx5nkXoWrdzO+S98RFCyZ7IdgviiycAcmAK6akksPMiLEEqV23OjCyn6wSyncqPNAL
urJ1DN8fFgJJPZk/X1XAKMc5AJNGAHAI7C/AV8XoUBI0Kxj6heVDF1uY9h95/K1G6fGK5hcrfka5
Vf7QmwoHbcr7U5CTDqGRfAvgjOrlu5jcFZrdVBVEO1JdgjSSvBHLBLM+9o7j1k9pX3YcG4ueIpY6
MVf9OdcWP+oDcxaRmYIOx6sDQcdEBh5OqikLcVgQk8SsDyKRheUGtjNhMaiEhTnnQe+3t8AzZDjF
phhIcyt0zLr5lMGBCm5wkaLqcnyqR/S7sDP1pQ/d8uJbx4iTNt/yXCUYT2M01s0oT+ZrbfNOrSGA
iiIcnTz8JDCfzRzFwCmgRwZpXNR4IVuTfOaWjfbcdeiUw5sSwEJiz+D+nbBCuqyVHrABw/RjVFDX
ouqVo12klhiJieq7ersUCOBV6lw+rgD4oNEMQ1J6VMVlbTVroWuaizm6q44LXs0S4UT82q82jKaN
hWAivjuejWIiLfIoemyGdm4bbOSKMZfEXI/SUfANYWYRkGYqgK4x4qdaj29k9nzT8/0Sp/N0Gsch
ubQUPtA+Bq4WuXDbNr+CnJje1cZ4LRL6hI+B3L1RrW0quFdCYBH72DFRfWu4XF1VB+OE4tGk/rnc
pYhp7kh6EhhgIed4WjnhuFeumUh2qQeiIjKV8GcZDTPFdl2/3egrMngS322q0bx9XIPxPRR3iBKm
PjDdobb5lbUy1IDpDKn8NRqihs8pKraP0oUhoI7NC11Q2gdZEq6w/cug+BoeUPWBod56Ofr5zwu5
lSQCHM/enj34y6QG9Uut1dfxq/N2KTrbp1rdw8qrX/OEoRB2a953qaj8EXb1i2tuLHIM5vg3/OsQ
4YUb1k+yGiqMiV+frLIPs3L3GLE0FxnyH8r5quTb0TBCic+hw9QGG9UHCHp8ZfTQ52ACmbUf2qcM
ztgoB2mN3Ql0HHUzS2HhP0YSaG2MqI9VpzH+lP8DL986J3/UCZ4dhutu7xnn2wgrj5fQmN8wIRzf
jwJrJbUIGVqOyg/atkWsjhQ/753oUmTBJXZtl/Ymw8L31u58SpkCghgROZ47wGL4aJyxjrFpbcjs
zEW2w9RKbs/y2wg3+AthxmSWlh4pRblSmPp+qD/DozRlSAyp8c5Rw3D7LWYFbIFhcNXROAdWFbPL
hhx31lGEjM/VjItUVS4RT4lFIbw1hZaquNERGGcrDfpZ56qlsT7RcgKNvWVBa+K8a3kirBVA39lt
CMo7cC9R9cgCGrmDO03dDnoqnk8jJL00V85/4NJpOsOGt9i3UQj3FDpOTYfbYy8UUcA7d1YqkBAz
UthRoncoiUEi8VjOWGCuaqzMX87Obpo5B4jvqh+z42Fg6RvAkNWsLv1C4yBE9nsQ8dpk7u3I/ERh
XRDJymMh9GreaJJs4WmkpMobnaKnaPi2tZDJvExr+Uo5Akgr/ELzE39M1EzIej23/wcKPrmN675t
Ddlq0WL0jT6CMvIe2c6TbF9XXaegH71L/vdcWgktrulg48MI67XBcdaSToXVWSgfilNkH2elP7xh
UZmHzWeHOcIUNDkVrwGdaih2kxma0yxo+DoyXDzJ3ZcUGNWqWfWN+cZ6D/tLR52zj1FFbatOhHRh
n6NrTwALlj/a24Z5ENUvcKp6nVs8EGcycUM3x8eC2ykljva4xKGnBLQHXEqqxfA/0hdbIFovMatD
wujDpOXKAmKDDqnFVm1Vq9M3nRj/Ih48/oN3yzliJZhoBw9k5Ae5h2a+NEGD2egX/mASq/x7iYs2
waO/BNuFdwqzBnwJn8Bz+4kRkA/TaqQBXBxCisInxM4LCb0ZaqdgQrWPghg1wLrqqixQPNB6OdQA
JpHZ6TQx1dtpgxXQYc2/e+1+0Cj2afX5RhzGvFuRd337QASrg81Mgw5tk2siV/WidMl8s1Vn/t1m
bCVDPtJQyIRSSJmNuoUt252BKin+wRUZ1k3oVT4dEzscbIHtc0Nyk63GJpCHiU7WbEsgf8NNj9Uv
GH82tWU0fHBJttFNW4aLmyZlHjRWco1A44oy7JuVNdnWs2YFwd5aEm8F7dHcmxz757vsj8BKM1wx
tIB06AACQcs4/BjgxUY45Zj6+qIhc/hGCFj1U3u0BoryKzE2WKb5qsJ1gHjCgQ8WrwCD7FHjjyip
czyXVpylqAXqXJzZYkPBBOITd/Qf52cP/GDovUtVS3k10w1n0wWtwJjiNlXB4owuhn6y+pPexLAD
EHlTMupnSUygDi7yVB+fc1Lf3jF0d3hn7br6bvgP/c5pN9SMBwfZE/zQJvNNvVrjYyffZPBpWR0X
Z3kWI/rcNVZ5pPHh2vJLfzLdVKGuQMggYrSpC3X41jvICmSJRMSGYLIx5x3tj2Tz9s5GJq1W67cW
Wg02hrkIoipwJLqx2PpzgGgEFp/VgjUXt/Y7jvtPI2L+Eb+uBCmhWmgsKzb6xBJk5p0NHVlXiKrq
M9I23OpLMRCh9b1+1hG1FGCx9hPSOh0InPhUA/HVd1lUb6piZuIa2gTw+yvdNi/Tz8i+FiZMN1OJ
rgKK9A+DqztwrERooBPo4dH7AbjJJoFsNotQuityEoGhiFFDqWF/klcoUGWKq9UE/8afhGk+gDSH
v9jx9VbL53w4sLTBy1A2DTEuyymv0WK8Q+wNFVInbS+Rudb8cyz7i8ginJ+GmAa0x4YdB8Ojy4Gx
iuZiNJRDYP35NwaETjNZeNLewzvW8ui8z7IA4e3RuX1UvzN8CNny3EbLaOj8G8QDWllPPiyTzupo
FvfYao3E6kpJqBUtzS78gu7Hjb0VJ8ongK8uoIIiSxQKRT7H9bf6iyWHGoB4wPJLBuYObwZxZ1qJ
bqokOiRhM6FHg6CWnGo++dUa0Nqfj6rA5nD6k2GEvELHXcNOLQOSSnXSbt7yjsixtkpe0ZKd65dH
nW7sfx8HF8tc74vdYoRsRdIhXRhaTVJykgEf8axizZmhkvD86Snj0O2A5N9z8YANfiVL0KbeWC20
aeSzGfiv0hV6b2F3T9buVgUblHLKyIuXpBGOmrvBm0o29K1xJifeZs485sqYO4QoPRjMKYOSD30k
p0Pgco0UfW0KXCYD/FvdlKQZrYAAzGbst8WArhxOjZRuwsnawDgcafYaBO5oY6vUE2SywVn32cwI
tDMrOXBSDAp8qTMZEuWhKp1CP15he5yZANh05RQhvOHXx1aq5YVc8t5NhkW+zD9LJnt/A2Yp1LUD
RqwUxogUqHqqtQ8SdeRkbuhySeggcnCCrFjiNhSFB1A1BcMsJF/8u7TJV9HWYmT3qNTJZw+hl9/v
+nchZ1/7XdgUE4v2miREUPL4JfoLBo6/B4BzeMZj1QINPg7QcCZarcTru4OQmLeyGmivWPRFKDz2
yyH1UzzDkpRtsxeuf+/ProxJV/0Gw9E8mUlscs12LuopSSr9pIrxivLeAD8giJJM1DFcs9/E0ogE
DkDCKaez9aBu1k1qJ4mYuS8aqRFQgN2Y25ZmxdByXrqZ2zwYyxsMkr/5m1PhS+nKdZ54nqTiGh4j
jB4ir79A39XZg0raY7m8lJWZyGmp4s2u6+OvkwYDVQg8vIWpEBT55c3PDbHOQQQJeT/WY25wLUrO
dQrOAr1WoGGe+MJBqvIGAeas7nK/Up//e+B7WBMl0hZ6PHeCxPejPKQ31y6yPgVGJhzqZ0PnYa7A
//aeo180kohup/03JME6gxYmAm/XK+va9xT7p7dJ3mFbhVB/eFlhTnB6xz9fKLJKGbh3Z0mHldBF
rV/vsXA6sORiAdyMObt5xBqz7eBeZ6j+XarGeqK7XV+dxR4VR13+BjlKmsI/yJMYHONABq16AbMw
bFXsAVryi6XsspCdXdVrV/s6odvyT9YzSnIXyJpIWW7yEguifarrQBCAVqlsljCrkw72U3S1St26
WfO7eNTe690YDOukXV6fPk6Qhe2iHH7cmDlyUxgqD2vTV7B6sA/XN92GpCXlGWCFZpXfcSvAOmik
3sqXqwd+gbAJ0cQ9t4Art7hucUiMYggyGpyc6tBMZNiRSTZB0sDULW2hCWssrACdKIUvru1EUqey
yw2QBJZL4+dyNHT5OY2KkHSvQ82M8SuRS78mbtPF7TyCyN2X7TQOqEaUvQ7uf2sAm5EURwjG3Zy2
dYtvWrjIcMwXAg9sWNu2LqniVMwKA0Mug7BQZFjJEGaVNAlGnpT8cgN+AjpeLKscVuR6rkqf+1Qs
Qhgm/s68xE/OldGF+yhR1i6uZ1457h6u802L8vZ+YEQGtleQmya/bbkD/Rcq/UBSIciaAzLmFGTQ
a40HdvZwJLZOb7cRSGgz1EBlF3+6u4TWwR2VBUER4DaQpg22QnBSionUavxZXSU1gftp1unTQZwI
8tX5yUeYsfoJFC02uY59GGbDV8NTcHQhWiZOtOGJU0pOzeAywUuGI63UKADh5+8d1NpavgyZxgQ4
AXi4vg+OUlQv/sk2W59HzueKZupvdx3I5adWJcjiIlR4kRs1mOT49Gk9aJCx7Ons5j+Y5abmqoo9
9excbKATQQfwHajMaK0do3YEU9caUZLS3V5aIrptfffYWayJ8GtAoYyz/oFkixR+J1AhGKy+d8Wi
OalvC3FVNcaR/x2qTeS+lpK2y+HUPOngCoFOCwDYp3WLKkoHqJTiAx1VfBxA9LHr6Z9+02Nqngqj
zeMoDk9tU6TCXovB8SR0GAILarJ+H4d9o+wykhNxqStVaUWgulPJxpQJHeFymOPqSn9OiDGtWUrV
cZJuJChYng0r1gyEDqJQerWzg+h5rdWCURsH2cEMtZ13CGE1W13fva64QZVg41bbjMh/uP690Oib
GsVJdEnVOhoLHZ5Kp6kb9lD9q04menI6iAIjAPtDaPzOqohwG2XSJoVYP7komOXXAGDlilyVTNV9
03DQYAm92SREv3Djyqfx0aVqix6GCVKDB/dyo836NIrCJNga0rG7oKIMwpzpkJhTAQw/G0GG0wWm
nCKoK2kXTju+VazU27aS52jbJbagnZ6fnJ6VKBrEBJHd9ywwarVKqiSyn5mnd/Xn6zuaGT5s+oUV
NBdiEGO1NHOKVp9wEdoXGG2QNwLO+SW7zPGZx9a865Klm9L7ji5AUdnnP06nzsZBs0m8v9m+wRYl
v7rcPjY8IWc6PggWidKtWAS4YwcTS9yPo9fW56tgePsKj4mTWEXBNU6LUBJMGeWXhlh/0YX9kQ5f
kM8kTy3PRvTRu4CJL9oVzgDXeq8l2M/rTJ0xDf1L7yHy2AwX9ac1o/bCOxKQ+OPJ5jhfSVLPxDvX
nInyl9CHXsDBhLBf0ja/4ZXfWqDXdzUL6FZ/ASEuhFZGEkqsMvGrGgao8Cl5diNFr2781BzeBS++
it76de7c96M+EQP+k68Rs4MDGo+T7s/6cWPjOpurMnYQZg3VsxJiAQL7EgJQ8t0QvbQGp6U1OiaG
byqNlgJvWMpSTL9cAjmSCOIsaZ93h+adnp2jmWLsgEG0dyTQibCo+gMCBxk6B7sXvFqoiE5KuEJG
OK+dg47LIiRIV6tLU+8dik1FPILTMbUh6sexue+EhCvbkO6Sfg+bzTYypWBy4X0mRBr+XevFCbiS
Pv3H7neRLyvQ9dBEmh4lZSm9qolN14ks9SFfbvOZ9MsDV6r990HbT/C6x4sf8369GfnwhEHD2XE/
oXq4rSRJRbzxFmJEhMHBb1PhszqoOat5gWUThxwh8Lq9Jk3u7D8l5WW+m9Q2YdIfgS9zh7pEmOLh
Q0my3L+z45iRf4VV3gtnKr52qJ88vkHpuHi6GyxjneNDWh9epZRToqv2wcVXLcq8AaRjDZvUfAl2
KP5NTav2AyHNlWc1GtbrnP/1i4L6NDe/lecpRCFKh1xsLwRoW8FNMQGtZAZtbphc8r41dZNEI4b8
nBovv3So7TVsRhlCVxvwNIl80ihQD6TCRh4hMlFxhKuvGVW2a8FjmbbdYSR1DpniZ+D4Oybe9Ybr
mjx6qICeM/AFJJm5R0JyMWkO3V94edXkGHKlYF1AYMhgzR73a7XHi4Ws2dXpg4ITxE9xVoeuQuiI
nZ1egzf5Lg1PVkMDD7hfs6uFXx+zGlOXaSZhWHl8VZa7+kLsJ2iuODPyW8jxGz/6u3tOwd9hhvI4
96XIFzNd4zClWFJd/8ay4R1wnTiOuzBECXZVzPq4imXTCAnqmDayKgKugdQ0WLzTutuhHO2b9dBw
m6cEzDhVZ9yFobsgL2SyI51vcw5T2x8KxJfLFycxwqjsh+Hlr/qJK3rE/l+xjvplZQ+AgGHbmENn
zGI7L03KyCXzu3UOODP56ZJjlT1An7EWL3qhaWKENb074H8hzOJra6zhBBYu1xfSfKEJbyFyvGIO
7eDavq8tYuCwwMRdm4n/lAbn8DWHpAFUAP8IayRgQyxVL8lPLDXj8hGkPO30HfVb5RCKlW9mkFqm
SFBC4nkdMpNlWybIfGgMZHMs1VjTnAkHXFu2t+UosokQMEEHY2i10VvtWmYsrnsmi3w7/W7olV0d
UewdS0My5ET/tkehDEG1VJ6JWRvdcfg69ZuZdwgW49RRGuXdSs0SJvcm7Y/2ryz9UkJrFC0pL8Yz
w1SLS4iFgfjkq3KRSIhiQHHtEjt+IZFKh/dg1N/xU/3R4ES1O0oRfQ3cR8ryYcN+tiKOPbHN4+0R
WlmE0GPPxh9b37L2NHTYAMUVg2JE0O6K7k0l4Qw7+6m7sFOtmqOnUpUFR5nNO2gx4D1/7XfeZTnP
a5/wNLJcqjaeJnemmiixr9dqbd/GefufP5isBTJghe9spbb6ymJW4djWn3vva841fxw7lzR4RnCA
fZey+nEuPLQlUBC0TM20n8xdUnhyxcYmmvYA/jzPJfGGFaYvlruqF7y8IFfWRqFVJKrIlsQEkRrl
o4e/OCVz0Uj5Szc6hwShre9gbrcXaXVsSGYDQaNP77Vl44algTKsxar0nobP1WY6PzNPaAPUuw8P
iFmhcGyr/pgyYUg8khND9S3dzJfuKgeS57ppN60WLuyeb4lsss0k9ReBunjiwARjM+6cqnlysv1V
YxZ8YI2wFqLiUnolombORvfPVvFZWaCdhJ4sbLYN22Y+hMAnulIE1SzLvBKbAykQiEGSFI8F9hPu
ZXV/YD2PzGT7ATBAC38EPIHbcrIS8maf6GcL7+PpkO1HeS+zVwTNICZROAMiSO3r7p+Cp0X3CtKC
WkP21+GwPPz0Z6dgCj/E4TUf1rUlk+OqiOOLMraRlT6idHGJrRkc7QFLoVlEewSC318+foH/XF3K
Y7sW5HobA7M/5UnE6h/Q6W9hHCU2+S7+mP4yFu5Sum8jm+nAeDG6IB6zRZOZXu8PFn+XYVQZ8m7c
oCEnVKKAdpwpHPnva+JFeC5hPTzT4ls/DLbB5EX+tPLZYpefgWbGf6Cz0y1oH/rAFDrJw5nwYNqi
eGZ8Qu3JBQEHxdtQTOJ+gB11IWUjwc0CkIy7uhtSyK8Fbj+GQmNsk6Ju2Bs1ZLQGILZPgRgIj270
PHWi7Y/Fzbh+lxVw1xEFkBrXDB/1yPrcbVH37AIhaf14kfFSZDvaRoe3mgo7HqJjeV+nGcqeN3H2
Ud75WseyHfC+Q88Lhq7oRU432ZsOrh7i+8tOTT6OEqp4X/Jvj0ENGAvhbo/oCvHZ+BiQHa2ws3nU
dzMgEDk1aghVC9VvIiMSVC9FQ7RUIv3h16DIvctVerfYBaUKE/X2Q47q6mXUDTDdrFGV0euimJiW
9ueGfI7AzSetP36ueO1ruQu5er0oGXjZNWC3OdJ6AgcZrd9a8k6/GmeKwgkXry1yMc64akR1Ko95
3iaUuxBsahE4UFePAsAU1nArpUu73hyJSEqu28GiSasaI33R87+rvyBDBE3CeHMuE30RBZeEMrH9
ix22dSTgnkdeR01/785y8QTkoSLL00lYh/PBqDPUFNzeQhAk5hJE+NVSjxhCKAJmxNUmMqVmdHFd
4VIJmy708NTuXp/KyozE2qZ3I+I/cygYUf2PgS0RXciDwWdeffByPLWa6eESKnVCBOv6g16+340u
rLBqFh65SJc3DrW+cLNCFevHtHYVLzati/nmzR1xZE5OZGP8L8qRhoEeZcJlqo+Zkacj+upuqNEx
tH5o0JRPYQ7igFO/dMez7Hgt0lxWt/9OeTEebFe8Bq/j3JH4aM8D/oIp4l7RY2jOadJlkDImmXXd
a3xS+pkyUVNmOgwW+1jKmbBe5y2jaAKIhKk/5oDU2JFiUyXPE5Wqa6b4yT+ICk7P9+K3CqcmQjdO
2M4n1ZQdZWbgQFr1fS/+CN49qDvUoBlftAm7uF2Y7ClVGDBZdDGZAflQTA8SX6l1fjiDrDaXkPFX
OaC+KUAgvrQ22wJjxmDosBgLFo05RZVIrz7NOdtl38phTBj70REtZ/leNmdhPWxjq0II5wDNvWSc
nZqMjqVI+iRnOltKdb/XO9L+zjllh41xoUPxpHOoUrnj67a8u5eaLRX3+VVkw496+eyMkWP7heP5
3eV6HAcIrxdpR67qU2vjXm8btXJJw9HpRP7JbAyQUCukHavUyh7MkbQZx+oGMx9nzMkciNoSPZKg
FOz19flpUwz9cFB/Jg4D9kdBBIJQYxw5Z5yyEM0rMxIixQzlsplJM51aYb2Wz/ZRMswpWSSfAqp3
xY18cVl0zSlxmJd0RSMmaZdTiZ8jKeo8qf4M8xjU9iE8UTp4C7v0SxxCuXcVNbPoWXzTm0vIR0Ql
CVQciJhSKvzcgjIND3NtdkLsxwy4qdQ0e3wNWwdeQkpdgQqFheaFWOoFCSm84EQskEHMTClZhi6u
UrlyEWN6fcLLpeokzbeDKQ258dnJz85mt7DjCSfnKMViYQAng0rEbYn2iZme2Z6KuCWk2YzLveXi
6jwbwc+LhF99dXLQCRXYSmrA0BZaw2S8s5i9KQTTjxQh87RW+qjrvaAPDTyZE66Q9zMOCDQQUyrS
x6A1bI/icWaLLQaGNpbAQpeRF/R6drCGNvFQ8Ehs6FCT/9j+dmbQASEVUhO4GOrZ3HCCUNcxy4tJ
vC9BTRSTrU/CF0yTLHiMtqYZ8COFRImKM3/was2R8Xp+LmcFu1zhf7vKEYpq2w1YxLe2FM3PRqbW
q55d7IK3DTgHZYFPa2S0bB2v9GfWg7Rd7YQ/SeFZXRrIwfDcEzlGIHc0AewcwDnke+16E34AkQv/
REOGvu0rnm96QH9aCaSA55S0/hJqFVkXG/lgJI5T2xekpLfOXpMqcj/F5OLfOt58Rgv/x3faOZco
u4/QT7cST7uKI5fYoQYXi1CJmGy0CeFVAbte1zPw83P+14muDP/o6+jnHF01guLzxE0y81shCv6s
q4gpCRWcZYz6DBlBLTL8VdX/M5h82SbOd+kaIMEvo+roViLLzdojRDEe0HM4QiZpQmIs/SD/QSUM
IXYAdE/j7LlXXK0f12QBIqI7I1r37i2cMC3X4FfaaM2rQrqWCuPFf04jLOr3JxLGGqYGiMqNsflG
1D3CIIwUtAcRm2B1fnFUxzfJgBWrjNqCdBxDu3TP2Qtv+6p346W9Y2Uc8znTJGg/A8TGZ3UQ0LFJ
Wj/bcReQtWJR7Mr+wwK6sK85PEHSG8dXFls2wVjeWqz/YgrNemtxmb4cRc9fS5I2SVPE8uUwpZ6G
o7PTF+KXKPgZMdpgx1gugcOv/6QtjoHOzplZfXMOC5717tIlb9UQa0p0AB+Y2Zj2F2EBfomtGcqw
7lLkVcix+BYP1i0VkLnnXAXppLr9AqMu4ZNrku+o9LTuyVYMCdFnTPoXzl5GF0eSx4Pq/Sb3iUhs
NLUYwEIKDY6UmamjFvpzv8Pm5rt+jTH4WdGBDKls+0BC01g0iqpUky5ZrqzVaWJlCQ3/zdiM4dM9
+a6o29XaDoMdu0IrijNVsCHiFJcjO7axXvmJFRC9Dk8ScZ/1R5cKoomekwDotbLy3fx207jh6+62
Lp2JSq0UPM3hewYFtPmf0yIksBjCWrR7jWSuL8oeZSjSCXn2wnISPRg2Qp2TlmeufySrbcXYiF2b
WlU39ECewuj0R+uEAO/ZzwmrjuVRzA0gC51HOaup/wQoXEP2bZTDUAGk6fbAp9LY0tX16kQ3n1md
L9Sdpr8oWbw6V7f7te0Mb1/xvqBxKQf+q3pk2slgtykMZrpYe9kJ/Ne9VSaljwxGC+yIIBaR4IbK
XfEe9GdL5P7ydpDFF0eizi7m1f2InxwrbeQMXrLP4XMHIyIiPigzyd+hMNy4R3yfj7mx+siolbrb
u/CBB9SWtIaNtrNOf2GjqW3pU+OoHylfor3qgb8YjYpUViViA6xsrO6K4/oL7YweaPnmhZo0/Woj
P0Qor+iPMsVSw2fd3FkBYzPYtoC1YnOt97PR7kxezb1d7BwvTDGW/pNvA4/WtjIE6bObRMcfh95B
U7exQy7BTm1nEEISqyUXN4uDp0pDio/9bxwuooEFq8rhPMIQyM9ocaw9//ZbuY10khwzOt32Df9C
DSi0vpzbFZmw4l496VrEMBnhc8zZgJh8VPp8J+HW9FqB7o7OHYOLQ5IsPF60BvJXTVvy0HW95y/1
n7M4BYoeGw8sakEUCll6NcbBc4FsY6BX16Gu4G1VkdrxxSJDUPhg0AZehuf4yBx6L47TK6lipYc0
fgSqCZbSz8Gm4mu7ba2MCs2BxaiIyzCRpLPHe/dmtSzQeAJNB6xYcaxzR3SHu9CsBaaK9M97JQF1
cYffEmXbl8bxiV9fJl47oHsxfby48ooXKq+HjG1+aF/+gzCazpEw3zeygA2/wFD+wFndRiweeqBZ
Ly152Wti0X4VnqhS5v4b4vMpxXzSKP7xBNwH14Kcx6kaex8CJkryPgfg3/3TDWpZDTdkVfeFdg4P
CctPudxdpUxwG3A9+IGk7xqg6KKywejkYqswlG7agt/OqJlcB6veY47cLWZNYltl4rYcX/Xuyy4Y
NmGZTCIq8eyJLWmoDk7ncGDrSWX4tPNgnHiRoSsHJ+n/hFOcnc6jUtCejTpXfC4OyoFOqdoyz97o
Mj7HHeELyrmgzpU4wxp9UB+FQIxtpNrD570E323TKTTZBkaVWNGuCIr8lnsIdf2okUTU9JFhmg9Y
LJKGOkg5AE0XHJb6D3yuftxtjbEaOa6Glcd7zuHzhSCfRIUOI4OopgxG1W9toqZMhTKE3RSbCspU
xwAN+zFQe6mxStTIwmU2mf2RtvmNOxt2g4iMODki41NRCj+TZeNicFhtEhjkJ9n9YE51mf/4Mk6i
+6wPC6oyI4q7WxWzs7TjIgaCy8qgNKkXi1xnG+DJ4gx1AyCHxQb7dP89kvG1qAqSRS1eKm03DAhm
SPu1sUDnjvEaeJ4DYhF3lQWHd72IzBQSIChpMIZmc9KwcrH2SsWpXUj9FUlc+gAurFb4ZCgEccA0
/Bv3bLAgJij/7OeFZ3ZcdXuw/tUzDs/JAxrl/GfrtndIzxxUWqqpdM5yo00VAD0Ntz5BSj959lsu
Un34iqkjzIH88xgiDPkzKK3C5aCVeFwudNhUqwKwCI2d0igsLSK4tyhD5B0TUfAAyBgoyeWuHYzL
/WNb2OWODR7wQc7TGs8SywK4gdPyzk9HPNdDQQbgn728YCokcghqzQQJCc+rlUEy2E4qQjXYgIgD
dkfkh431vs9K5w3tqLZuumhGKYsITbENTeW58Pkw2PhkVYEooiGmc3ZtiNdOr6KtQgrhV06YUf9a
scnrTnKyVrkHnZwEbrA7s5kwR/Iyd6Q0A+vHKNTgJlu3jjdq4IdTAjC1TBOzFf9yh6qqLzRGgvpp
5T8OrAKQpQx3h5T7cIHag+oWXFdDd+jhsiFXapHr28hmuFO9vl6qR0Hxjf9KLic4I4a3kmoownCx
vOurDzljosm6p7Cd5dwefqNZ65fgbUmg3WkbjJ5Qt3/sNfzSQzu8zSeqDKXQHa/7XT/etVcToPwS
jqQlEBPXwpWMFzqRfany+52+0vCGCTyR7ldovrkjL9toda68CThpT76O9cvWvUk/GahEontwiX5c
Uon6ZcvcTHNkoolcquNfhPeTqE5am3hfY+6zdatVEjAeH7NNrEgAZpLkzoOB4g91Wtrp/iR3Q5dI
WUn7bnSSz3CWWc9d137P3NW3ACnowM9D1earAMtnVfPXTbj5H8Q9Hraw2heuLQakGecWnZoKkLDM
l14IAELQ4RijPQCQn/wZJ4+BNkJ6Neym5gKVrcIr2up89Z9drsg9rDgfHfG5HHNng9XwOqZOO/oJ
bF4+lq1iEwuSFjmj7BBaDUGOxeJ+CwQvDyslYv2FLx0CRqO71qcM+4U/R5Q3Q5pSBo8HwW+Fk5+z
kOVzZ1FtrB7WquajvZXkW0i/r9fjlmrcAZhEfWUp2L5ch4UWaM/33su+W6LTMQktHvFNu77c2gwc
sJdVRCVSxFbsFZR1sCqfmjbkaKDnX2sSTXObHL2AMvjkJGLgV7g4n3+HNnfi5tzr6tp3Bxiqh+F7
ZN7QaaFkNBA8l042yRa52A60Ar+JqE/AjsyQZ7unA6vju+jI/JWOY+34BJgrZPG9Eo5RXal/tbk0
1F2bImFugtStdBt141EtMmoPKHWtXXSeITzHBGXch/UW8b6ADbKkILikd0Yc8Nvushgusf/djtZJ
TFZuSlRsI7e9J/botfruDD/HuptjKGuYxVf53AWAnmegfgdIvgt4MjPK6LAvlpWh7O86+y3AmnqJ
TxJLw7hqZiya1WhMNonXgE6MSEW1Zj6hN3E+32X0i1Swi8jxBSRUWWeFUl9QHU9gCh8l+OSf60hR
W0cAIZtwqJx221iQCfK7LVlI3Xq9tP0zxi/UY/X4iqLV1wK8t7TqMI/lJq1XrCp8hi6wVMhmRfjX
tNrB8nSf94iWHjZzfcrk8wEe1AFzbQbY+pyuGcB2EFrRoCK/zXVse8SBknPQpZ26MzQIYMYFf7tE
mbKMIVV5tAjijgRVcCEHtE3Pz9bYCxCsikEfnX7mSNH4zs0hbUjxgxKFIpL71l+TuX8jZh3aBX/P
ZWJJFp8ZGc+eXj4aN3CK41NbA+1AIMwEDQKdSukCd+G2zNwcLJGbyBUiwIDNpOQIwAA5/rL5dZWN
rNgJK1zahQFEcqRC7Fa4fgSi6ELIOCLXZF1XdM1cQ4ZNDRqdQ1UNRXCqgzBCRNDi5N+VbSA4uF/2
Q1ytYnp5fYqQ6v2LEC6UZ4n7ktS0zYFI6gPV5bWz9LNvRHfrhPKOHvjt+0ax/ORf04lHyGBP23E1
w1BwNHxlowIY9EPklcPKKRwIflDnbtSa4WQ3xL13JfL4RVk9nSvQpgmSZiJJ0zfjiUCni/PNHy+L
5LtcaQjbDJ1MkB8KmPExI11Ky4w0pqj3AA2pg/EUKtc7l8L7eb9kk6eaHQvyNRUHDUunTMJZ11I3
yeIgoh/D5UcR8hK4os80RYeOcyHoMhQZmWSOmpEGdvmaeWuGWzHEO/FNqkOhywvBdrJJKX9+wutv
CkbHX6fGKrKyjAwB1SKrsg1PCtFwkqnXTWBjxKmq81jEo1FDYMagUGV08kIzuTRkgzjEHtIzueia
1LovGMisgZMBHdWnEbB8+3vfiAx+zk5MxQJgY2pjQVQKMg2f0PnHWoqUwN08XC+8Nw3tmSIYu433
/KmNnfowCGal4nolm+S/QpOkiXFWeYfxP+kEzgHbfmg7VLw5unu1pNUUN+totqLcSETWOcc8aix/
i1S7rqdVL27QM9CM2feIJGqbjWbPCDdmUtE22etEDPITLPdmtMjdYxchyxI/rVql47t2k2l2RAcz
4+RmCKKtdXmw24pptWx8kVAHw+M/X4n1S+SsV3qTqdpoL3sG3AgG3dwc2rZQ6mQuZ//hoS11Dwbi
9Y6GQNaj3yJ7M8pp7n4cTPW/9zPry+Qj3Q6AeimeHiIpwSq3g0pxqeXITxTjZZN49qClFFjELRId
JmFBVFoJHDaw/Ls2J3G0+5VM2Zk74VBXnHs50tvBn1gB1QQTup1/pbrjE5FCJKfopmvf3ooDa1sq
xp1HGCSczs1vB/pj31bXsrYEbRC+Zn+6WyMhA5h6eTNVO6UY/0yM+H0YIMoZe9nd2ay1dgQsW4Ba
R0p7DrrfPaAvLsqQLoQN92H3Fu6IFFXkeoCtucPwew6ixKk9ngXtpitk/4wAYlzZNX8hp+cMZegT
gre5k1CcaGhWf4JVpXau/cOXwsTJLB41jVYuPQ5Q/reDPUd5A5oejBj76g0z73s7koKXeLaL5eVP
d41rNqX8p+wKXYqj/h3DGKN2PZuccxmWuv7CrrHJWFkawC7OO8QL9KPEcSVWtx3F8hCPjK3koe0W
JepfD2NZ/jlOhStOXckPK1PaM4YPMEiITP66TRwC5msL5iIR43H6xOc94rG/QTus+9vUVKGlpPy/
wCj38RzMZWVqBN9PwBQKK4luXtXn5H0WLC72lgG6IejPL9i+QeJrT4qbxsaqU+QS0VqCyACaw6md
PIat/AOgxTPOxI7F54efkB9NSUbySLUsq42IA8ik2T4HADsLm6rxGNyIed5ymD4A6ckChW8CYaEf
VKQ13Jjrj+Hs9YFV6wtW1qMlJ01giXSkgLauOYZueTUeHaORyvT2DXWrHGolmb2sl9OQ5W5+SJn9
Xm4KKvQJSOTny+fVSMjLGdOKYVNtHDzzgjri8yV+bwGejhYwb2F9jivm17h/7yfI7nqFwjcdBtJq
6e2IFN6j3utBTcqndSMaEzM8lWrb48BBG97k2t9I9QQt6bSuod0VdgPM5QN0PQPvDtGrBsw8YSjS
TZZnGUQrNeSmX9NHCMNioZZVHPBTkRdbf55owflAkxIsueQSwuuzgBe64dQvPP90zNMQSqHD+xtF
P2EZ8ITn6pwFpoEQQLki5Pe1G334vTYR7cfUALb/l1Om+gCtzZ8OLOiOeA71TGS0wYeWqKsPlpj3
PsY41SaIb2Ij3YaT4qtWwZYnL2x+ftc71AkOHH2PZbXLHxxJbMQ2yMkTR6zywv5HVZONQiWjNLTS
Jm4KHGrV/yFYu4a9xiewXnXdSO67cMkJYMcs2x84NkWquoIqviuXclGyVfbYTwAYjPQm5Cpk/eoA
1AnNtP4FizFux/MoQzL7Iu+UKq0iwuAiB90/PHsTg2H9rVA0OKpqOHo1f4olrmgAZzyIH7YTqsr3
FLT06n6JMxa4uRS6+rNx2+UshYyhKdptCnNqg1R5q1I5lOWrjemPYn+wnQKrSBPK6OgzI+W5EQ5g
NYOO3V+iLBRxC1Ozj/YRl1Q6hjhqVPz1wFYrbDH0wXcitF6hI+lBdjxExq3CUZGdhlbN/LXCIn1J
hgiKwtawyYFH1pdcIwDASqbt96+SIWIWwmZFg8nlVij26l3E57o4BibD7Rt5KBIa9+eRT7zW0aMY
EA0x+wGTjiyeqf/iFbnQq7oFz8Qa2oBmjqdNCM2GlIRMuTk8xjhkrQIP023vYk4rEy4SW+iiV4Xl
oQJF9+KgtaBEmG6mTUTuRUVAyBVXO6Wn0oh6vzjSAfZ7zyY7+RqS+ABJyEcjs4r9YSRCxQOamHuW
eCmySireReQ0ZXTuVYvRjgNdapRkZ6+A7M/xbHmMGSvW338uTeLT3MLDu3wCT1pasBhc+bJ4XQT3
KaPfj8tMUs2V/gnzkKu9Kk9yfemUY6IPxD2UxmQzIkVVFOOjndRQtmdN+joc3cB+McDO8vR53Nlu
UJnRvG08xPP9jEfitzEeYuKQo01Vpn6rMdmlwo9UDehwcQl4Q84GSJpaK8cRn/mnixzw4K9hzEBw
4F0dTmoh+HWl3LJ/zf9CGuTbaqyzoCHrQR8pPtqCLt1rHsjTzuy6lPg1d7U90e8gUmflFbt2YtmB
0ldwh20zzsGGXNgUfJN0+qJKTR7kpUCVlbPKACgsWS2/rys+yKzIEhHzrE5Y4gfWqnBDhBUyChOp
hzPkUabV5xHfH7bthlB7LQ4Ky9KfvJpxwZbXYFHlknOVHm9tTmllvz87MS79j1IesjjZHcpkmW/E
qUOvOtg2D39dQmrtgP3l90R7d8NrtIgmqpXtEL50DPywdymREBXdelxKbV7k0EN4ws19Pqi0CdUi
P65yEOEo6OmQREf3cYy0/ExBf/VxPv7IRmnzBYYSZtAbXMcUdpjoMspw71WStx9mb5ab5B/7pYcr
YF0Hz7deIv9AXI+NQKr7ueAmW0MdwKhVT9RS7boudLsTUNdN55FLOG5M6SOuR3EOx/Yj70WIDM3Q
ySleN/dNUa7XQ8HZv+ly8lJhA40qn1NlhoLEE76G6Fix1oPWU2zJttoOhdEk/gQtmAebKTOwoeZD
55gr9nIPFtWsevb222/pANLdVQtK6Tvb/jJJqDox1TZsI3REhEyV2C/LnJyDa6Mw7iu3L79c7AcK
3nrynPuDnEVg936SXQli6st/QFnQG8WHcfd217OB5XPYHW1/0JCTyfk3pFLZjzN751H5XE7z/rew
HULgQ44nbPgVpPR3f8pXTc3NzMaOX2heNKUKFP4JEwJrDBMzjK5Q7ShJ0XYrNKNg1CK37fdJ9Smx
rH960c6ZdVF0s+qYlVkz2do5CQ8adWYwztWchzKfJw4aTHw1N/yvFsTCxVP46okqvzTD4S1FkzBA
ic+vMCUWW/y+5k0C1oSujkOvAFpzrJ17KkJI/HvEwqjAFstX0/yYW0o8byz/jNpvsfUOzbhwiz58
hIwWFtv9EqWGKVr1M5KwNZl8XY6BRN6Luk7S8r5aKc6kjxUaoCRrTsPhxpzO6c7RyBArxxp+qb7I
O0qbNUcA2QRgd8y00ADXPKGLEIca6aJ2fzGsAymzYX6+iSPQLkVVX6voX80MTnLTCBjcTzz4HxuQ
/LuqkdNJZfqaSYLdlyBLGRiNk3vFzSskE+n5ut/g+w0yJFqbj6V8XOBVPvoAIZTF48qudxq+YDiC
BVHa+9l1IiuHZ/jZ/ai5RzAUO0b+Flu6hn00qUxPFCmOhUbGPfrRnwEm0yY7LH91pH3ePHFrLENm
Y2PiubeYRWsC69r9OSQ+oL2LQnBpOUmJH/pn88eMarNrj1p//UUXVxbm/GZWvNudcJw1VLfP3g+g
JC9QhD+EmhYpFAWVHRbf5RHjowC35Bl8bOK5tG8W0SOiTbMFQy/LwiCNdRAZUzr1mZhXo2uT5D+J
5pAoO9rmBcN/Sa4pji8IUc2ntLChxGfu5iwbfY96adXz3fLQj5Vkit7DaeuDPJCboJ7qhoe2HvcK
yXE19weIQJSD54Hkz4b9Wg2XrIJJsd0n27HQrQyZrGIjkZAzs25RtKHAbATrpKJzRvXPrnM01GoJ
tWwaJKzUDuspqdyS0WlNOVnCD9E93WFxg2Y5ORTgmEumPChaKuAoIbSDf3MDeEbA8ofV9lnoAAOI
1ZfJj8Gb9RjZfQRZEOx8lz9myOcjQesQTpdtTVwnfso/lck8IXt3STGCj4o1YUDWzGpDLEQ+N53J
gNP80v+vzeKApMB6IBy5RRMek75/JSE83MXLVwczZZkdvUqGs0qY16hq86ntXHmjJTtyhRc1/ZTe
ITFA5nRjvEBFqN7WYz1MiqR2p2Y37HxxDHpeVaz38WRadGKgRskHdltNCe+e7Pod3D5aWB/3LFBZ
sKlxDBRsyvq81CdurZmpAU15G6k0bn49fT0882/CPYih9gE/8jkVv/kNv39mvLM+LtOghPhJJygj
AcyxrgUY9/uGRh5645KcDbuwaX58rHQtgJrC8YtY1kFMY8mvMJPzmXep24cGX55nOaOQLYstAxkM
i1S4UwA4dMaXocnRqbCFqTsjYvjGTJo/i09CMvxEiwFaisxzoIlnrY53BAsVnzgfWl8g9a8XQa6G
OSei6wgDv883spB4/Deb2KNwcstr6vWy3lapOGlfKjK46dL+MuFIwV9H0eDKhGfqwa0+bt+WLZXU
SA9bJhEtdgehz/qxmy94M22EtWbpd+cHwrgQlncPgZdARnfILteEuQA+HCZCqz0Xe0Ss2Dsla+6C
tI/CFZVDbPlnl+UwW4rHeMk3fJk01vh/yOBjjZFeNODnN9cApJEvoP2KNkIUn3IlbKiEoYxzEDNG
yr/AOTLUBg4bWNCD2yY0O3OXfHwsaqwwQq+r80CYRZMk46kTR42Qg932GDodKt8gU2YII4E5M8Ba
1O8hboEE1gjByTmfhPUasHq7cbg7ZHLGCDoM7KMkwJyk+n6ZCA5LOAvmGtKcJ8fnF/w+9/NjoGlN
wzrXrkzTUvnXwyl1uL7+PefDewgHAsEd5pU7HqhcRrsRVXKJw0YJzcB4IwjWQ12WhiRB9XysAG4f
ZUmOJzb9KVMpmhkcP+dq0utA78TQVhUgkVL8bovsnzXaVZUSRxhPWLKzJJIa0CbIWMdDZuoq7BLC
6mHFJHEF52VqmbI1CHVj3SzxerrS/IAlNFURvUt/MJQDhOfKds2qMrcpOhmBTMzouDwMbX375KeB
a/GGUhgKpqsWzWDfbjPNt7cWGj78GzKWx4e9K3tJ+12pU4MV00GkYUdp3palukR5bueZL6AnWTEs
ri1EtsCMjxMZfDp/ctL30+vvNeVShDo2Zw+OPJE+uUvy6DgaGuQJ1GaOjhmsjJfvYTlFibmvnVlX
k7x4hxo9F/45ZkzlcSkUlLU1il2IftAssrdXEu/DKeMTCfpTGfj4zIj8T0/9hs05UPfB4qj4aW82
YNpjj6KVUCyGXYThPkrzVyO/bYq78u2TD9uUHWMFx7vBOw0cVGLAzuAGQk87khJPT8rWlYrvCjrK
AzGfkec7vdICiFyrv/OVCHH8sREF3FCEY/WaHhqe9TBIPUwTiifWjYoK8lWdgRKjHym8JSIa99wa
ajpVoXvipnTkfByHnxn/qzNCmjlM7OM1VRdbAENEeB88pjclTJlvu46Yv7moAkFwUE6YKbkHYso3
X+O7RrtEDWrT1J50Va5mpByERmUNkqLwvtHtWFZph4bOsKlh6h0TFxfSILhLZ5q3K5eMJWD/xHRn
xn16krwWscF++StPBB0iR8gPWOsLqoRCUNtI0+N06uI6EBKuz2ubbnVFABjHA2Kuc3gN5TK2mQWm
7TqroFtjEjnrFf1nHk3ghJUJZ18dI+4gz+UXzoKVsu5m+yD6V0/lV/vkCxhEF7X6QfADF33X7GDV
4RXVZVN4qoh/eu9FgAwLBeBwuAtY0jN/z7Ef3zTwemVRC3XWWpRrZMmmVQKjH8NkEhg0ApW9IgmL
AgZWw/LfcOsXh+iDqKNcoiKqez6lr1Fu9Uy7OWl2LbZ6ZgVLmPawfIai2jk/V/rIEwYajvacIneH
dmhwuCPdsxONgEaIyjKWJe2rdGfFqyrMeNACGWtt4ZEqUzWvAT9lrZVoGXOgtXAaqHsH33rhIDzc
aWJ6NHqRnItWcItIxlbar/GtyKM/EcqQDRS88uOf13nkQ3CHMWuJdDU8LYYJqfS4FdAv2fRnebxc
ILsJqnPauGUQhkIw593+5uhiZD6y+WXztGyk6ylgpE4CyRYbi1PuwCdWPWBFLB6Qdqw64qTve7ow
BSW+d63Egt0OPN7ODM8cxAFFjQ43nanxsEChCRkDiYRWfZrvPOP3H6fUQNIDRtxLmaKb0X6Li7Iu
qDH8gbfAmZ3lpbwgQab9ozWPQCPcXdWwUxAGDQTcOYOrq8UbTMkMTuhMsOAlno5py77bF2hTc7MY
/iXrwGTLO+JoBPu85mCD4OGikpPGhiJZ+o4jMkU4khhWYWFpto5S1/xxcCg4g33F4AzjYQVbcXDQ
vKhWi0uYrzamehvjhNu40CKHJk45WAkLL3NU9U08BeFJDazw623bo69cxNCYcEgQFNNrwtgP86Zc
e7DbZinHtaeFUdv6DH51BZxKM7KZh+dV9cwf0V2xShO7PWJGR2N5bjdX6nKsksrAs31xsuRyxMAv
fvo4U+d6fvGCwv9ZI7PsxFeA0kV6PMruz5pd7nG5v9jyAnTutUDG0/IIaHeqAEmv/EiQxTirU+SO
trx+7rdsN4A41+SlMC5GZUSiPAxqAVcyiwMSOF59CqqimG6p8x+W28Vf5DTrYV6FYf2R3sl7wvEB
4S6jsyysVbCFmXfk4yQMG5WY+Nr9vzzQOIB8EvU8S+kLujm1U0snaWcnBd69xCoH9CQCSHkqAh64
uognxC8nWyGO/4XqOLzfsIjEu5B7qokitsEnBvLR8qVPdC8JJvXX41w1QjQVQEJh5XjXd1jGUIOK
RXB/1UZnJMGCV+Y33cT6HkizFh0qU7rvpXLRg120iI0Y8FTjdIuVyp+3vAPRr0CwdFp3SPCJqT+R
uYjgU6Qbx3+L7qYHsIp/qtg7BclkiVhvN971LXl049NBicTADsxK7RjWA03FSSRmuKu4ml5LbJoL
mwa/C8cx8YExL/bGnn/UreVNVbMspu3w/wodsfHSr8V5XhI3Nn0VOhoTvhyDwPnxNj9BJwOsGi/3
CdG9fDPl08h36nCYKMK634Ocnb6QUQ67FjT61cPyJ4HkTt0bWV7AFDwIR/pAZ0WttX+craqCPr1K
toYbp1BYy2Ugcg8oeXa/ampiFQO5n3i6wC4WX5WWTrrA5jRho2qtTlRC09XpqLFeccHQV65fyFb/
wOTzqf8zQHH7JDxtFUeIF7JycKDVlm/cmPeFFeLqtspbg0ikmMUSNtNnHfUx4dqZZtIKiUA7A+b2
yOBPZ6EbtZHDvF4AqmYu/qjcp9rFJmZfOhdp2NrhkA6NsXSlHejMOH6R8t5TZ5qOKek/O/TDHDRO
vXH43vz3pcLVkLfln5fmclw6QN8s1RlFu5zEh2oursN9DISzEbnweUb3c+UvC4lP8FFTkjTtWnO+
sDx3SP1XVx2+OkJWDI8azAiuQpWfMcN7fItlbGX1G3mMlFt1vv8AYHZkV6fEYMuXs/D3DQO9VjX6
jjR/H9n1mmuoBCbU2Q1BvnnTVgjOILeCXgpPeUZr76Ng+oU4KeIaL/UPS8rPHnfVkpu4VuaDdOBs
PFy208dEeOt1GsTmUE628EXmHOlp8pvN3/AQhdG6BSZEnrkZ9et5vaeEhh6GMufNQ3ea1g7p2AR/
snydZIliljOwOUalau6eLBNdZaX2oaUqEEaoc6Sqk+p0GoOcWTapuQMsBurDLjrc1DEU4eRWEGhR
X2S8pBDVv63LT5gXdvuuj2MW9vau6bcTzaXi9rdm4ZYY7mxz8ZmTIidIBUxz61Ns5/+gUKJs97Su
Nnks3vDsfXZvugw3m5N5x9UI3C75te6ppZzwbtUU+TjfMroLYCcoTU5aSSWRV5u9lNcLcpLQmwji
2AODsv1JRMGdKLz72MNIRuPJ9OReOU9wrPsJxN0Hd1AiG37GlbQbzz22XBM+ellJ/lCC2KD2Rphz
FgShT7xYQmQhqogPBz4UN+7DK9QtwPTBSLYzFG8xdrLM7fG6c5ovSL8WCQ6pUuYYcoyN7h1sTMta
QLKH0Df+qs0HnjySz7W//7jNMRjL4JEuv4ZLu6D1SWXX9KhP9C6aswJkIOmiy9Ar/YfJqHwF2vcj
4vSxCATWiLoz4wvHwiSIWsfLrhAmCbiJjCBozmR6XfO4mU7OMMOlilhvk62tLnAZvZGhzqOtIu+0
6PNRFZj57hsxEiN3L5HBDicLMA+TLeABzkRn13Rs3tzXafnOcznwvehYQp1W88o9QtM6m+vKft9+
6OpiejZZw45mXFjuO2PXxUIqjSolyUSxTXFY0u7PJ0mPybOzc3lAPjNyaVDmeilSVtOGXUEVuMyG
DaezBkmgvL5fp7JTAwTEk0Ho/bn9Z7R0DejFD/2EO15Ts4ONeqqL1+f5G6zmK6/jPEXeNWVdjxuv
XosxI+iZf8Fa2mcf/cq9VWJcB9YpZ4l6jbCKbsQM3bQ+Y4XNwByuQlMV1YLzGj6x741SGev/yAp0
/6z/3ZWcPrsEqxhqCyMK0jPjhwd0HwPqGWxJwWX8s/9I0hJYp50FqCd2O4klxE7X1T/T7vFcOIjC
u9S4mdTzZUkFSCPD/cz7HdMuI2D3IL5dc4HnP1ub7NIYT+xhJ7O3EKtwQJaADdlz1UbUhpvMGcat
dHjBiZDCQ0jAUdm4EUClZ3gMw2XnYZMqfrOqOkHVqIqQj+2IeH8I3FrKCUx4hCu+/3zW8CdYuwvn
PhWXLFJbNZK/+6IAoj0wKwtKbuI1pKUvqGOSpch8aDf+g09loemQOjMjWnqT5Z351RxTR6TLrhwA
pBduw7Ea8hxKbItqxd1v56AlBrQGRi9+aqLOEQAi1IbLknDgzUKLjcc2ExsLrI0HBWouSn4ZoQbK
1Z7X/HfOWYCbQMfWYa4qKbbKXMXbxiFhmEF8r6XjCdbvd+s4fXkxpjIt48bCMFWcJ4vQ+se4CGRk
rxrOLe2NZkyqDfHzp731yMCWbotNMmN+OmpWa8BIOBu2O2Y8QThWxJWrGdG31VF61boaL9B4j1DC
2MEKWjAfH32NTzefRJAqwOCcESSqRbOV1m/kBtc6g3G60ikU1PdD+kjx4zqdKChDc0d7V9a1yxKR
H9U2y31QhdrK1BWhOnu9jRMt7s031LVwmtVoZ+OliOOeoIY3E3M4ZkD1kYqh/PwSrKlEqkb9Vdph
dumaYRJ81XbdrWfFvdjm2HNWXHX4OEXOsg9UKWFr3yzLCpHDLsZZRjgsR7HXTNPwXTfvJCbg0Fy5
u8nxkdz+3QNvdQliQzH2UoGl9ueefNY2xLq0MaLWIQPRf7RqV13aSa2NJRCPCJ7BNendWbsOcpom
84pAwAgAIifdNGkeGTI1XQPsDyw6xU5O8AfwR90UC8EMeYg6BfqCDzErsVs8XPMqL+grwdf2mEkS
mAk7S7QaBmlgQ7hJI/DZFgVkqIIqTOMU7UHp3qrRxaN0ibKaa0fcYqJ646vHoSLVxi+cp5skp1v6
aP+gfmdk42ZhbjCDv75ACx7P6sjN99ljJHfxQtDgxzZhUoglH48pvISrkdDCtjsjdYb2DUGtCLL1
xLIPo0Z2F2NzjiQPJAFNaheGaCFcJYOR1j2XlyP32eSVEMNOJBW9zfVzKbx9UP+7g6sD/6nF2ZlS
1yjEvQjUQEVWJI0n7PjqHddh0F23OGvoZ9BILNYayQ69p1zrCFALosZYvrd+qy13/Z5tjXd2ygwN
tcmeOyY73/UB1NCYUpZ3gcT8lI/4liCyP3KrjtOB9HqrakgXne1Tv91YLvGkRBX80xwz3qILfazT
sV3siwFm9GzjHGdVRkNt5ICmdWSXhu9TRO0EN86Lf+AmsGdRjwzTP6VKbt8q4Ib3a4xiIO866FYA
2CIzxyHNl3JyouhBfHWi7Xuo+6QNZsYSA2a1qUtpZnS2AWwv6X+VWCzz0MLzm2shksxh6aQ1Y0Pl
r4BKyKHg9ko5fgNMaZsH0z3NgpiGO830zgw4PMh+Rq5q7cvSdbtKE1ZQHY0t6uHHLxtB8Otns1hd
d5i1MyUXCL34OqnjGhxaoZatdKhYbzg29ESE8U8QmnQdeOq1HF3eRJpxKoDKiot4OI68xcMEL73A
JP/SDmFueL/aD1UPx1NhuwrxQ9vlJyfGYIXSwUtMHQTLxvX2sxlU4SY+wNLO5jE7J9tV1s2D01k0
ckjE3xY+zKZUDCFHl2djCUvIswRFrpYj68PQ2F0KykDrzTdQs1RxpdKg9tgNiy6UO0Kd/M+pWytl
OEcl2dhp/Tsm/AyNQdouHmcWpE1DSbq8KO8mCOKp8xgG8qBr46VzNascZj2aBLo1M1A7ahCzbyXi
1vAlVtTC7utjVIc1mg80rFlVYJmYLn/yImeWtZn4AJOXv5pnOxWPepJ9Xj9nvSCSBigYWuj5Un+l
EsaukwYeYIR0a+Q1IdqxGHngnkIxte/xx1I2i4OVUgDGpPQjj655Qd3dqll5HPShIOyLHXAjMWdY
n2+OYHYYmmhVUMm8cLEWh+BwRkUFdKwvFVzDS2QKBHVxXGL3iT849DFbcJKn3xoCZIG91IuSdLIg
3p4BESLrNEFB94nABj1ZcWch/Y9bd6XStftD/0T3KMc+FXYjykY8jZVdu7zumyyJH7GV3rQwkrM5
a1QXSmm0NXJt6YULTkwkE+F5i7oacgMcTQZiHKADgrpF7aGpizNzPKjtEqvGvtv8VcIvnHGlqWkh
HXtBpA4rXUFjUcq2tuMZ3NAq37EO1C/0eq/WJqGJzV+S85rWQdNVwyCDNAPr/eH3BzYQfyZScrZM
9O0hV3GqQWPalgcYB8tHeWBLvVn2HB3P3RjWyC9DuBJoxCXDZw0TETbFMMhiQUWTgbHRD/RV/7Od
HGE5Asxol+Xrtx90D6og5SxMXPVZWF54pplx6uGKntCXYrXDVDDSaRnM54S0FT/anzzXuWQMPYp4
69arI5bWYNEjCWHp02LYIfpt78isuE3B/5gKPK6ylVcS8iK0eMeGBilMCV1W08mc0o3Q60iuo7l8
+Johrk1AA3JlTU1qFaUPZQDova5vADG2Sa1IYZn2Mk0uXMBmucjGKmEFtX1Z/L0kvwXSID1TLSxb
cqud/Y+llpuAmLLlvEnWWbbKqU8cE3HwVR+2WckLbr8F4rMXgVotgr0yRWHUjCZDyUIn9QcEELJX
3ZM7ywydB5lVetcPzdZhjXixDLWp65F9UdPlcX9l7/74ZiOV3mR4JnKF9XynZsrPOmx0vDlsv/ye
kdg+/y/bFRRpTOSwTeBDlafWYTuFf7dh/8tNemZEl+j7GCAEdm8R9DnjBNGV03fgDcisginPFq4H
i90Wrt0fM+kWyKRLDG/HapyZ0XDO5ym7Nk7BSrDYGAvTyXiWv/dhYAsjC/5MshL1u0WRZY0OLm0z
6V9dZpW7tfJ2/gABbNGj9deYnv54d2uLreUYXcm6dWKWRsgbPGbOJHBBUlUCOtc2wfbCHmW8xQGA
bHEjPFiR5hjs21lBKNBR5RmuphF2f/B3ONBVfW3VtB4LDcjpu6Li6EJYsHXeZDvZyywN87rc5W6w
gmjM9siSV12YVaX7M8Ay+lNEntNWeCEaY8zsfFGOaZKGpPw2ooh82DlwRJgyQSXDCibCBwVyHZfO
XjpgFRJCFpqwSpwQNC+UUVoFTWvNb2w2oFBb0zJqSEBCEs7eyFkkOEdt2PD9yttxk9S6wGA/cAJM
FVDaK1NGJXa2h/a9e4GUyiI81WYUEsW7YWYweMF2qCyvvXwa0nbEwOWvqPVjy/hW00T4DAy7c0lW
1QID60OYppCJc2B+AgvKNJlsVNO4+tCnqGT5FH5eUmpMJu52e+INKOrH4Uhu4O53H4a4Jn6d2e0a
GbGFlHBJNkFLLxY1W7r0VDcXY8RDTt9pbFJhzQm/71GdlfNmuaqf7Rm94Dk6hhgOIuv5y6uGSkJc
N9nCqFAUl//X97r0Jyu+JOfiTkWIRRFwGJmYHD768cCt7GXcKDzXiMwh3IKYiQj6NSUyBseBjxP2
c9yNhgDu5Wf/D+MvQqeVSOJZSKjYNfHkZucx989ZARfCIgJ2y/rM5jT46rBgEBajP5+ZYqcMdA6A
3iJrjTxrXMVEXkw5J6I6UWnB8O9gud/Q47b3UdCtzzn91sUSnukZbbWpiv0CLu6Mew+12qAYO56x
2jbEaLrw0cdcPiyhD+yRMOY1hu5P+zD3Gixj3+B5mYMpm2xkPwwerZrkcapslz3VbMlfYDHdVABx
5QRoq3YrxmpL6CnzuwOD1UhGJFYJQpZ5aTjDaVJr4ON1D+2UPowAkXULg2DN3KwQlLG55j8ZEHD0
qEXT6McRgexY2jYhge9uXEMVWhK6pni++YGTwevX69ua7XC0fnK5B7/NqQcHWAnHNNCaA8NmslM3
67fZaZlHSeT8xafAtK81y+xABm+s7ygwyaNwX3rErBG6vyjEhGAd3WQ+S93lg8HLtjp7yvnSKjOK
C78N2gtUXSGUCp+q5xsS8yMTapEWD4uXAdlHh3dy7R5GUfFeN4LM+nup+yT9fPP9dmJ38I6vW/Ia
Py33BbNhTGXwnAB5URvlAp2Z+GqQvpyQTlZZD1QFG96tWV/0HgqfmfI1O6FnuyePStgGiWlzk0+D
s61cLfxKcEIZMgooINsyhqap4hrNZ3BoyM0WsdEB3It7JnustO7gmSa5yUYPLmSbX+TUYl/yR4Ms
DsIkpGirf09g4blgkNl44w8uai6CpW3mkg9vOjNev/b8LfVNxpi7LYNzhM5Gt/Qe2lWdtEqnow0w
FV/lFcYN3fcbK+d8mA5zBmnSOrXSi0Nmby4yzelHMIate7UJ0tmb3rnHelw7XMfgigbVsosjOG8A
luOAhL8XR2Counpp/PaXnkBhai0VHTmYSrc8X6Yxgz61zA20QZik837zrq1VvDMWjO8XnVuAzhV+
IGf3rl0X3ykElMI9QatZYOmp0lY0c448hmHt6xc7anYa9+JpHmT+1T9/vB6amw1KZfPxy6Thudj2
G9zsP8bCop7+6Ul6juz2aYMBhOlXg5gvWVWFflba8bo1pVGGbNhWh8oUSAbS/vNTBQzkUNtalX+L
JpQ+L9imxkwB3rHO7U0xIvGB1HZwRN2UGSuUFF42l62U1UhxHW8fdSL7/MBxzXClNaSkhW9NVRf9
g7es0uDbGHqV2MpoJ0Tznn2vI2VLpMQO2GFP/A3UQWv0LIpmAMTUcEf6hSXFE+sgKu8q0XAFnm3D
H4w6qJtRXs5RBR6upFm7FUqDB2DpgJdDw18+REB64XxabvguBJNcbhjXte5QW8SHsxsPBge4qyg7
wZx7XXyBk3f8hsIi6ktJl/kbg7yK9hv+NmzOQJo1RPi7eXREDtAyLcC9m/4+cPgSje3h0y/4FX9n
berZ6dUNvcWsVF+XJuaYRolgYcVqVn0Li3ChIfNAiOyT5RRjT9OgUy+pVS0cBN9oasPTAtVKpbv+
yMuVq8tId940u03ICvImA8uCRxGACvRvJwaUXUYGuU1b+dse/W47+lhsAzPTl4JCmpqljIqZQ2pm
bnSZMfhu78uAmRjlDRFjfxYGyWKzqTvkzzyYkF19CQScey/6vYnhay6XdIAi3St34WYZzt8ypKfR
vXdh2qdL2scqlBrzBvlqscG8leUqGGXNzWRhKBBIpZ61sBaz5gkGt9NbAvtd+p06GoUAiZ3y856B
qJfe0HbLLZtY1o4GqHk/yZbl9Tl912fAJ75wUf/Y4BVqGTbKwBKTxKvTHcUHy490z2Gk04mLTszf
alOIl+VX6ovnafpL2Vyc39mqU5/FIWO1K417zpUhvXUeA5HKupXaCHFBStG3/nPba3HeTmHQWeSj
sRvCARhNuqxnWZPn25TkJm3mZqvJ0+zn+ZivArrMOXypDTEEYK3dJyehyVlTdkCEdf+3iG1vzJpN
C13YoMWjLjalxCRqvf4lioVfms/nO7Fg0GIK9DQvOkQPDtRAMLL0KRet0+jgEf7g5+k6itBpUd9R
b7Thl0y6UIBUVM9hLyETrx1u7tY9F+/GMFJuAQv+UCtQTDBS68ZwCxi++tkqjYOhVty6PrBkZkCU
G+LDOFvxyM4AvYV8Hp35vCWO3YD1KSH0oJOegyS54ZnlHtmhvvkU4dVzPZycAAG0bExoOXjwPyHr
b457vqFDBe9O4/khC9ZcSXtg1KnSEovsO/YvvGdwhrqOmzJ6seL/q2brkkrT78zFXptntlQwoLaH
CAXlii9xLQPz0VgUjOGB7ReUqFBHVDrDvpj3vasuSRmrMbUUxCL0qgZ1yGO+VS9l6jjei/sutgb/
RAuDU9OWvPnRX47PfM+NXBp/6kB3hK3Db+1iKN6NWceUqWrPRwjWu3XxoNNf5rqx9SvoXMJg9faB
c6fCXUghozXlZfTs7LOxxtbi0pJiIgAH5TchdBMZ3kSd1VQlQyBsoDtpUHaGLGgHCMiiZRQgXYqt
5qAzL1ublnLUGiW3i44I+uAADGNThxK2P+SWExrjFeAJxv/cCG7jWf9El0j3cjMrTRNWXIRQzhf3
PRe2SbkNVOAVQ+1O9HmctiuFPpsZScfm6q1BtZS68YqjDxuIKiKBWPU6UrgDv5ljJLs4So1WcqVa
U7bBx9pts9SaBBFRi/HZas4PBL3BGb9x8rYN0crAu9XOEm2nX2j4Ro1zXRkko6hvUE+fprGQR/LL
0ha0b+5DwUGJSHe0mIMfbEsL7dt1PyxGKHhH0aGuutEWvMvVVbESGFw7D8UTPseK5ecCM5zvNslQ
8PmM62EEdn9H6u2vwllp1bu1KydIAjTVnmUQIUZRSpMqLP91RyD2SlG0lt1rgvZAd+D7kHP1/7HX
OoVNhRbBTaUgQ0srInHHY3w1K0kaKWhVPsXugK3TyazgKbJT06sB2CjTHHQRCiTDG2vI1IgSGYys
FcWvySqITtjI4yTAHfZapQEGqNZjaIvBpO7oVufw4peCv3IZ0wZdoyv+AF3jjpOr6Hn/sk9Q/xUr
wG/JZHs3NG30zL8ulTxe++hIgnTtMxYGWIcna6+85KqsW7V79m094S6GrfgP8dIXVlaDl5AYl8YY
5OV5lKx/mDIYfzMsry0ufJae+4NhnefUUlDMq5JxEUynovVesJ+a5vWoSmgtujwb7cGeFZSyyISx
9kIhGgZeqkmS9IYafKAaj4JMkvP8bTfMdDyffE2GetLIeufzpjOx9K1xFqg+Y7f8RXhLrNZ7SOGD
BMLOxGk0rfjGpRcYHnCxjqpEwNBJglc9r7Js+utS/XS3BHjokzZFKE74zK6m8IKjv50pcjEh44TR
FXlhiii1C9vpYHruZhwxlqDINfNhLgOyQH+e70TR5A6+cXtWO/ETSVLLJriv7vWMndgV6eOb7wwx
1gMjcWLp0j149CrCCSG2gKVO34ciX8EBbXr2UBYqL1E5G4tbPCvECfFOb2ci0QscWSRyMNkhDE41
cK3UFwCllTu0MIcnyKES0RhI2TE6q+LtaunuIjIF+iDTj0ZLKXPy9Dd7ulkIV4piyxEzuvI4/OBl
VOU1vs44nktv0pze179KGZOJWwBMaaVBPC3rxgPECgtdcIvSDe8w1S/xtcREuAyS0CJlO+r+lqej
J7GNjY3Uuzy8Tzk2mhZhzghx8KA4UOtoxmnhE1UmL/cSgoaCFqdCxNu4DlmBUsn4cX7LoDO+rZLg
fr6nVDeA1ExdDoC+f0J5W+6NTe31+DwKb0SctrLDZVw91v1l4bPiYehdpL8EFfjPXD4LWUazAspY
IrDTPoZTivTxIz4FOdRkTbCAEXsGGYwPNBDj9OEj9bFpqIt7pEiDxD5ps5ZaA4BoBNajtIAAcav7
p4kr8h9QrjcFnkYpElYFDfI9E4whH9PqRWq9gAXY4q447qE+RFrvi4zM4Gtvb5ixpDZEU6BMQAbm
cSIa1cU+Il7VBSS3K50vZo9YYy101zQc5Lp7x8Kuvq2L+QC3mcyaSmpLW9AYdECo1X0isomg8NOA
R6JLCMfzcK8QvKCrDRNxnTmQMy+5NrkhVMX1o/sTldL4KZNvoeyiejbtV20i+xn9CTxn1pbpqSgm
iC7lvt8mo8rMGNfR4849ucJbd+MlQW8dFfDtA1FcgksWFfRxqNjZK4hdkGqn5OLghJlncXB2zanw
uujAulb78M1Sj2c3aVygO+s2Jk+KMl74oWF/SZN6yW7lAgnCIOEeFSXpxAH0Lw0S94OTg+A9hpsl
e//SSIbNKc/yPo7u9p5nWRDrkzWKAFCIowl7Xgj7izGI178/ko7acPJLJK9SpaTBEcgLJoUdbRVT
46SL1/SPXkPwWsUespH/5KRA3uSLZJlVIPRHe3MtxmmcOjY4sWou/i0byGKT92iBG7W3+jBoxiNY
WqsT1O8eH+DrMD7Igt1qLNxsP0Qaf+l1he1O/ge8unzZM3caH0ObTMAiVboLM429p9U2CDNumVN3
BuSgTctD/j4C8vy0aeYtkBRcb87IN0+iS6y7MKYKSTvpIxFJ/eWYUI9FxlKnxKyhvww3paoqnRZW
tF2Yt2c9VC62CDih8ksJM9AiPWMDbmwCcecJwFRuWWruQ8y/AWvCukdo9MwR2cWENFB0nBwNhaqU
7yqsm1bzZikz82okHe3XfBzEmIFWotwKRflJglR3CNviziM2R6Wn28lXvN7/RBDlTQkwIIiQV6wZ
4bQnn20j4RxgQsfyOCNZsQkYdTj6RtrDr/R9kwBeiMWDHP/v4gj7RhnhzzqmjuPs7jTIBYkzjfri
BSx0cnhALrSH7s1I+y0YtL8u4pgrlDvK9gK0VkYGbfDCDLQRuYJuUWwzeGnHkE2dpj4XhrfIAnHF
nPCPciFvths51lKIeYHofwT7XncXRcIs09I/acv0ekJFY9B9uwee9kCKiYNOykWGZx6xWjG/1qjZ
XRGDVfRRULhc3l4/CYW0MtyIyWzadolF5yaJwYsLb9pwsr7YoBohyFNmzOR0HO4r/98skO+zu1jQ
GIJzTx/UigMztSKou8Lm2kBtlLFgc57YB/34du3SwAIsmxP5g7lOwiyTU9jBdUKxQU83QapUdi+G
gGzBAdGxEp0A20D9qFN65SZNcd3wFgV31U6qwXN0diqKF91Mj0AANID0r462gYHuf8B1qJ6j5MO8
A2ZyFdm6rTVkgtOaX3U9sM4PbnPfZVcQlpw2gLjN0pTAE9eUUtbKRDd30RkMYmr+kT9BQUCHtKu4
fL12bdR5igJrV+aOpmMWVUE1rhiYytwDOSiEuqzHoV3i1otb5Y+DvsDlbS2IbzqhC2B2VQT0yY4T
rXVdtaDGVEQwhFVjJdxzdkrMVJ0wlVF1k50PbE+juBVkjqwFAhrKQNSn2iQGmkz3aT0MFwlYaXxe
YJIOBktyWVrCgsty4evcZsg5L13VIKuBEBv00D0kZMEPCqGTUQ7/eOd276irJApBJH7cEtfyNhs0
2Qr7+0y/vn0HfUbfl5uqjimyAvdJM8W+MB51Xa+Xoh+4uHyFHA9Z6kb6APpA303omZ8EKDHAbcoD
Wzq//KlTTV9BKORFZNS5UcxV758yPoL/7pPnPnRKybZo0bCQ57voI1WWSmUlLFbodZI4JvKw8Aje
SsjwB107otdzcCyjJkDWA+O12MsBPs0itfHR+S+Qju6U7CWe1XgcpnNWC0F9edhPiBHp/ZQoxU6X
bO12ygq4Xzl3kBKDrYcmZ2HRgd3WwbOCtvIe1OL9YxBeA+6YVYsEfeVdaUPjD3L8IG1EyhzSHOmT
avhO6JaaGYCz58o8f2tHLN/8TlaqEYo0UJAuUH/M7Bcz9ZX7qxh/t6DO2i0cqoTw48fUb3i9qxha
B+oocmSMH+9IHZbRtAo/TIBWSfooaG+a3kbFjuzJAKJxQPGDfvcz6JgYbU1gcW10FMgY6mkzKIEW
KuhQbc5hsda8a92/84lnDKkw1W8fJssX33uvhOkrEs+VJlgB39b6AQ3u57hugdblt5MMvKHcAwRJ
G8GjLFeQzme71WQFUgGxG3Z16EwcURhczGPtyKOeObL+vx6T6QRzebw9oigmdgIJzJSrNwyKklN1
t+I5MWiyqY6EDQ16VKUVRzGUM8XdOZBPu3badR/c9COJFFSQkT32oSvy/VjG+xGP2KyaL9/aoNRE
1G0ngn/ZF0JMjDzPaYbdj0cTW5UvQTQJW7+qHvsaVzls4eHoJK6G3gqrS8rQhi/xPrjqrGEYmbsA
zUlkj1KQkNZgp+bEO3fZRoG2DD2BsTMOB88KgkiVhCskIa6+saV7F5zgM6yrXwvwrWKE2gHl+0OL
spsUEiCx9NTY/BA0NFcFdWlxkRXChAEw3xbSLfYzGceUsXW3OTZ0REP0h12vIk6taeQgh7sKLOy0
pny6ec9rZ64JW5iuw6W4HY8IwDQBIFKyWYap/EtiETUbS0Z5d+ErwAC9Q+48vkPyaBNQwqB6O2v6
p++SQp6njjWtA/LEfwg0Ck7egdGA2XJltKQUal6oC+pkIsrFTIY60Lk1IAIRpQvRcABmqeGTPtU1
27jesT2GwTNjz7Xq1AhCT5LOjWGiLTv9UlA1DmU2Qx3Le/A4SGaTUr/jok0ieMrU4BOMYPnNoeF8
pQBgsOQVEXXWbw8j177io5wmnuOjQAWYmG3E0v3ivuHZyJ6BwL21YmbnjzW75o+xxYeMV62EKjj4
6tiLNIjHQRCoPzy0bWxTypSRxrP+s1oyXpPEOjp3nehkG7VEcsYirJaCNnE5ztzXuFfGnuNeuhZr
5A4r4mcH5boVS/W/F4Nj0ucdXgYzT6FXu5SFmdS29d2GvUAZJnpmFn54/1mUHRNSZgU/L0pDYsOK
Q/y0Qw0kdKMgCHegdMAArCM98SHxR88GCYzai5ONXGGRw5Ph33sWryR1RMW1hMLWuKWAEJB6dhw1
9R2vyK27Z1Lq7/2jjN6axT/fop0R3U2yU/OfaaJ/bbfMyHp85/6B4R7Z/Pbx+5y/kwJxWhbiZ7ZC
//RLRwSDC75sKu0JdeO4MlG7I/vpKA2GOhVOUjU4/WOOgKahpWaiUrLAq+R85dB2gSUxEd0hlpMc
Vp5RBH+4z+SHtQVUn8RFWAiAjad8LiD9AQNL+RTYMF9+eCvAppmZkAuzYEHLmCpIc1jpMSKrT6mm
07JtOdgf3jKUAAri1U5g/r9RDf/nOjmrRW421j7MDybvB9s57fCETNOYxaiBUTqgtHfCDUSk8vkL
RIMYunv9l0rDUPffEs+L+TZ7ynTO8zpU6DL/5ROgtJOxGUtTpvacxlpMZKiSFxMIADpgQONCfK5G
s8YAAlTLAb7Tucw5/kTpmL7K7PK52nD8ISCBq6Kl0/SzzwyMYvxXWfljO/6vW83yGyT743kd9p8A
+ym+UmFOUI/5L7qe5db/PuGycVo74C27fqtOmFW7a757zVTpLH2SaNw/DfrTPIxvnJayfwI7Spu9
QxyoSNKf2QpeG9FCuMLv7kw2EQHERnO/KoIRQbxQ6lLI4mm2s+FlNr+oopL5yFcVauvbJEP2dDEw
s9xiPW+Zc2ieWc+pudISMQ5GkNxw4fJs1q9kLT7FALiZbVf4gelpvJHt5pg7TtI1SWOydkuWsN8e
tozlWHvlj+FrE4Zqf0VLv2fueEzkVaoEejaDx8dSOwDYFDsm6cs5w85Tnz18KCkzCFrVKxlPRDcO
gUj6KX5G6jHxWWZj+DLucxDHN9ultFd5s6O5dB0dfW5dWp1XYX8NELKqmWJdcBIDUd3UFQmRZVtY
z9A7kiLU2z2RXdITOrY/F137ECtC3NiDRRVNIFthWpGMX3Gs/FOtIw+69Ca4NEzYoz+87tE7q0/L
6JsZTPWLyjVDuoZf2HP6UUMDZ5j7GUzPkeo0sDtdYh5G/zJRNwtb+xHWLgecnxN3AykdreNMPLkd
h5N0sFiy22FokTfhMluFnpRHklBErqe6AvLoW3YeryRYwDIoN0/LP0kNSCTX0voVW5rO5V4AilJz
6+oOCr1J7+N38/H+h0rL9xLQwUXnUG225Htectf5NIva7Lvv6CYJto5lnVCXgZQkm1Yi6IONgeRW
iY1e21sUCf2BSOv+admN2e7flcDoQ2laNzM6eqJtBm/mJCcs8z8NHVSkcGdGHmAHuDYaW2QRkKnw
EOk+waDj7IfkdsG0iv0L8yy92TsWnucLeLOE+b6vvapC8QqHlfIofqb6yeDRMXyJhNVFMhy/YkG0
jbzcvnbmoqy3xM6pavimgKGkiBcqsGocL4z71jxzVBT0auKm2PAm+hv/kYdiUQHQhAStC85lX5nA
hh7M7DBXSSiQaPcHJGWTREswR7NGNS8h73xVWjLQUAvYw8da0JR86sAfwsIDKEp1RAQjUPKFuqJ0
ZHTJ6Qtgbu9Xpbdm/BqwyemXeg8B7pJzzL45t+dYI7FuY2Ye7VOXv+D7qEJqSDHpFawMPZMC8BZQ
VBN/k66ZqB3YM50BO1TmOZOWyrdgfg8y+YFUMsAoD0R2FyCnt3fi3TftlIr1xDYZGmA4xezmwbtw
emA8NyGyRpCUTGulzaz6gDnIvNUJBSon+7NQVF7L90EPKpjtzMoCPsZ1GC1VwSfqmyb9Jr8p8+KM
a6AoIYxALkLGAowVXu1cNXaWoSqq7IqKbZ9+Pu3Rxx57mFWo2F2kCF25Ex6lPH+UTxcP7ZPZQ2AV
HkVtrwB765eXBKGRAjjgBn8mi+wPkMVatMZxNVJCp8NMzC8eAQKtiJE6o8JVSeL52+r0W8/mvRyF
CnHZ3HIrVgejUQcSfZCwSFkEt8wsW+OLuXYxAjqTOVEc43jkhY7AQo36HrWu3+FujThWfOPYX7nn
wrRt7DO3k3VBmzLZMCaJ5MQd2S+XUnvvUE8VULI1znDxH+4AIMyxsQjmKodDXLX52DFQ2Q1n5UVt
SxLFVuNrIcL/cSmRmxnJ7UJ4vRky7GrOfuQoTPiSHyqJoTPA/46u2wKzSPGzQBZ01dabmattEeEa
K2NW/cy0ZixCWIY0hQdlqvLMWu7J7oX/HKAyt1nLGukPu345F8QJLjqhmEJp8qFcDi2G66YPMgGZ
OdZNOdVnqq9eP3s1q28YLnm6IBiE2xwfvC0Uo8O92PH3b8tbpIyngszT0VmDiPZp8USTSaaVQh5G
YSC8RS9pwv9vSlZwGfixmxvn5bAmL+m4MbeybYTnynZab21h9pp6t1RuASImmhIx5gaVy054vTtQ
VC+1Y8ovLuZBYif9cei+nfFdCMBRj26QDzRisx8XZu4uq19DT9YSR/Zvn1uiCck/dKa1u+lTwgIu
jbxQ1nhKRPCOHGgpamSDPXoq1hR71fZQ3ULCwjquZlzbg70GD4Kl9G39ZI2UZkk9UFky3OtBff6L
Avx+4UrbC1yPfkrL3QLwFlzzpD+2ftSiq3QRkcj91lXSNBowMxcuKV+9GdqB5a8YGES96TXYh1Br
VzcdqhNRQN8cJE2V3qD9YHohKJRur6kbPoyYDvBVtHIWk1rRqqhBAeQhM2hdIN8SMB9ald8o2WQX
PZaPVZcsDQziOCZjkr1Dm4sY6aW7Ga3yjcNoIHkKa13R5vXGZ1ExM+VibVgbiO392wkMQ+i7XJDO
sKp5iI0gJ8qViiqaE19t4Q7IdPQtpwbQjh6ya1gzwqtiVQoHZjT2miqh1/fWS5ESmMFQcttmL2Y2
jI2ROBNzoq7b3+wHhJQRbdqXcCbqQVSMHn5ZNswN4vJMPbP2pmpqO5W3PoPKjf3lHg9SGc93COTx
TmC8vXUy1wg6vdQkOEZzH+uNlCmIQEJ5LahC5ea1die+7VXkTV4iUcl5Xy2EioAwlpxFxI1V6pCl
fir3KcmdNcDDDGaRscsr/UGWDG6X1UcrKXGeV2y9rb6LwSBwvQLpmn8Q9/xVlTkBl+Sl8sjUnt0T
5iWurE9r84l0Cide4tNlWmhMYpmOhkFbV/teoFZ+vHcI0yO/xfYEfNfnHBKjWJaMegyAGu1hFe4v
p9we8xKsEd8YPLBvFjAjUuxklGU5846Xq+SQcKfi2a7JmK5RZsdA+7dujQhZZIXFCaMFIJ1e0ZT9
InveaPna18vmQJ3u4Wb0cb4Ioc+hqOmnMEgRroMCBNjqetbcBQBC4d1ek0zyDQT9HnSb5PXMxOGW
DY86pfPnyjKWFJJr2sc4dUfWmXQxhzfkt93SWrQEyxPC5OZhUuieRK0ykXH+UiGwInEOfn1eVxyJ
Y1nCL+47b/ivDy/RGe/2490YjQn/EJmO/X21GGjwAj4QPcyRhIcbBPL1qE6YsmAKnZIkNc/A0U6b
gWwYBvPjgVlh2/n2KmZNXkkBFBRk1Kh5zwIfLD1YgYRstZLJVl45kAJsEoEUZdJCxH3vTPrrwFhE
2UJ8oqL76wip6oOiS8sRSaOgq5PWnoWAzAXL4OPAdUsOI2ZUslH4NyWM9hEyPoA/yM+lVm0wmUkf
aPCzgQHAJctG7ejXjf3teqvAhJVwB/iLhhjTFGhLwXQXqPGJLkbo/ud41Fa11ZPoPDnQ+QPGyoHC
1gHZuFsJdD2XW2BPpq8G1qWpY3kLeB2r7hIlRkMuv/VOr8FKrQCgkRFHXi92J0oozUQnk6VDUEiL
GV5ZgD6lTdEcxzhz+RBMRYV6dmzoaD0yHmBs793Jzebe9nnwzp/3AqD0eJlWh41knBd1uFm8UwP+
7mMcBiIwr0I2Sjn1gxJXE/rwd/M1+J8K+V2DVK0r0d7j6gPyZ8YKMgzF+abVNiWSzjGfBdUEW/7X
fHzH6t34mEZV5s87oF8W5cgTieVowXPMGtp+8CYWqCfZ1RZ+uBDGXZ+NeOxC872ZmCzjXtJZdtez
qCwlYD5TzcpXVOiyfcij2WQBCTc3eO7t3f1PnQ7wsQ6A2V7ckkCLilJXNJgoWzE5KsG2qfsbvOqh
5hSiPSqbM3w1kiczmrQfO69hUdTDHmLZ90jB3cj3d1ssQqoa1YtPEMVl6zSPqwBm/vhsfxg5tYBN
jkduRkbwx1TBGnEHSPNCiH08Lrf7y3pTg9QCBqx7i1ynlS7tBAlAm053+S0YtW/vuqGvpcG6kcwj
r/Z8UhzHgMYsG1VuL1DqjAg5Qt56P0hCzk7yd3GM27pS5BVmQQl309BCA3Bim+hoxA2eFUNioPxo
2dxf8PIAJgFBopHjcyqwzKRqv/P6X52c5X111JOM3HdVMUa+9oX26QV/7IpgGsAmAyl+9bO3S2uH
E5qXAOBTRrQ2g+N7oo2hO+6uB16biNCTwnOCIw+vTI5aFZqC93KG970jZ6bmPnbJb27Ilct/QNdr
cwAU2Ar1yUcLu1ITN5c/AymoKxovnVQ6qCG4SscqicZYqViIQTmgXqE0nZLUffiBFoinh+EzYvq5
ln1f9jNCQPHveQEUhuZ55IG2VDYUFJL2kH1alEdbmx2u04Y4Kc2UaiomerEftjK9znquazSvezLq
jNNqItJo8f4M6hhI7muza1YvaxzsqkxvCnpmIOCzY45Fpukz10Mav4qHDsUHvX547zMAba8kQSZi
g5f+AAoHAF0XRlQcFyIENDBtXQWkQr5fc3VMRVxZnkLPXDYge5QTorIe/Pb3Axlarku4GYRu5wqH
bfdGT1H9LxsQ94UMwjLSlux5RaFy00dzR02eBMRpDwCsfv8W33/B9YwqNKopEzUnlWxu6l0DZ29a
o/CBgyVcwsVSlZYK1SPgBXe4ejQtb2iRRN0q2YdKjVqq1UFkKXdUHVVUtoEXTEvq+lv9DXyPAlH7
NWR6eorkW1qkgDKHwyLV3bpvadnm33HuaQqrGpNixjQe7foSSiMSQ0ByjjFTcvF37fmPz6G4y8j1
dF6qz0IGSRUIZCBHt9cL/ZCnYg4HjdJYhb8oJgEBz0+SUC62v0S2ZLHr3kwCs2IhiTrvG7jOcBKg
gRpDtxFNIne+6FCfIFiKwo1hqkMqe87ztuhzdTjIHWNUOGi7vxbjVX3UBR6kL0cjSgQLPXqYn9QE
cO60jrkOEOjIXXApJHUT08GTHmALwSs6JahbhchUYCopnYTbWbQHxqGI19smsuZiwXTEgwOSaQtd
rBXcXJPjfslqv1S79mNdKAohoL8QL/QSHPVKhbvMwSGvD3KX/+lVJCC1ZtkdWpG6TTMU1jMVG0g1
fvfCJwwixsgU0wpwBWBBBROgeiHRcUoeWoLSMjEGeQuE8Z0yk5ZWOhMZoX4FuXMajhYYP4Yj/QMS
EShDNggyUcGCLHOGycrZinXjrlv48TYxtSkqwAzgVImc/FFIEMReXPav/KDNPUIrg7DOQiJHYVlg
2H/pKV+3NjG0hj9q4OYt0bP0NZc+qSj4McM9Mom0YccFFwHEw2Cdoz0KusYnmNDzDsCgYvJAZMeu
2AhcYp/7D8oRlkrWesmIbS/+WNTbpY0jr0+L2ifS3DUa8nxhjZpF8QibUSc7U0EHePMRe9KCdpnL
DULlWph5BBmdhIfsuMHDt+1JljYJDMHtbkMEIZLG8NBlrY4GM8DEVoyA8GISE6XasQp0/pSZXy2d
5Qn5yIWsG7hJxzETLiCKGdkClYZOUz8g5RJppksTy05jKXZboRluEWP3LtvlJ47BYxN7VBkgp4WA
eI7T0ICxyKZEZ6K1H/Mkw9OBpDS5NB3G4eZHfBI4+6olvrPZ2TQnOgQsV6fWFEl5mafYW7tF9lab
3/ygIZDRehxSFK2MGUfxTljao/QUrQm2ucTQU9yUqzuscz0ereQET8ruj/rKy8TnS8nnl6mecmrR
ZxhQWGsAPI4OyW6+u71eDS9c50e2n/hgb+0bcs5thV6RQfZBl56F9045G8ZwZfcZgrmgOCJgB7mA
4XxjKimXuYpUHKMPyM2Ylp53b04Rs4myc4hVS1WCvlnIILOE1eyZxWcbWsgv7lSv+/aOmYrC9/B+
/XVUzjjblhx4ehADftXvkth+teZJzx8b9TeS1seHFIom3mvGr88Dcbm6O8T+fegZOYwreKiSxRqr
dq6GdahvQMB6xccZQhXZmrYxKSJSYBwMQBZ2UCaupHCSOwtWUp6e7/ydaeAOi79pTFtxHspJ1ZNV
JLfJsv6nNmyd+kUQpLQ89o4dH9AkNAM5qYaHI1NkqcfSZ7beQCrjmgjQq1YNggKY5+w8Jx6FwkTJ
PLjdbzu6/thE4Ryoc2bHYHOjNuEs2JQrhX2BKYQd6sMcyOUeEF4SiMUaYgZmtFGk4eG9GNij+6Yz
/HK+xsuF50OrfoTiGZmLw8LGl0vICxQvfyiiQM6KPA3FPlHlLKEDlZp4OOeK0xKZxPxascJHKtef
Wymfz3z01elNtD3ej2zZK8pwwNWBdWbuvoq0FeN7JDFAQFjVT0hs0sLuFeLfosges/0dE3ZPERbD
I4Kg5BJpnLnMX8BMwDSVbs9e/1lgj7yLUhY8UncTPBtVeJMYGtEgJSEYUQ7LH6fWkvvE6rBfg4eR
TpwEV1Y1w85y+/Ih57a4bea+VjtQ/LpxwrJBaAidew6OkyXKnLPGo1YHf/bhy9p2f6t3PgOvhZJ9
Jn9wbhIxYmI34MqwX48BaEkqop6IOZkxzOml369FbeyX4ydPjQrfmSwvF5uzvKynvbE9GG7kx/CP
RfPgJf35MRukveUU6SNmtqeFM5NFG+5OlivyrqxRQs93yg59rP5EC4ivFHqud1sEopk3Z3lBQYlQ
LWFN5INhk5yrFcd4mUzRXm/7tWkXQx9UVl5rvUQy1JuB0LWGQ2PTmjBUiaiEiFTZlUYHsGfFpDTD
nsXoKy2G23S5Pn1UDD81jiauPkD8vDqmbu5PvzRBOYEGucEyBwgEtY1kbYCzCJpZNRQF5fA67tOH
SKxBBF9qk85T2jXq/+izQ1MfXfsfxmev84fJC5rUbBrmMyMN6pToE9qrLGp+1irYYKphHEY1XanO
cNPnlztMK46h8bcbyQPbmlxsdIL8QZIsbMMJeeMctQfTJ3w9iULpptTQKeonmUWSv6KAr+8iegmD
MWj3voixIqv/Zv+Gfajs8fjguN7zH1mIvkVCHKV1O8zJhfWSxEOSR6MFtaYqqqKbFBIXxt1GbaSy
YeKmg5kxhKGnnS7lxEhtcyOWQlddj9HR/ZYXhwUEd4HV7SWVzUZy/cVaPg/gKhV34kIW93/Aj7Oe
rhZLeMcCMewA/nnDyHF9R0guyVmUIA7frcbui9OIf7CzSqU85w8BLEExzuDhQBXWz3/gv4g1pRiv
cHoyZa2NaSWqioP2eBlrz+ylQ7Btp9P6WmuUobp9kUYs7Ibzgq6HMcXtjuFZqhL7BI87y93e0M7e
x7qXC/km8DJiMZ6hXOestJXUnZseSdYMdlSt29o+sdde2nhRWqcmuZIdFl0QmXWHYGXHqKdrGlFf
EGnX9tdoc+EwXAwmOQp+m5PpK9QV+fNR5fjlt6jO2gWaigxvBHFnuF7LPkSf1B8j8pTsLnJQepkq
m6z1nX0+ymHyEI80x9TXqDZNMT9LZRPISeIVSgZk0Rt/UczCxHcpXfv+OPl4soJGIO1Evu1SlzQy
Y+7AE/xvaApxsBBoZ4FQGgshYbts7nXTFpV5fjoqvOVodohjyab7G83+xx0ud/yx7n+g85BxG6V1
TarNHj7qPGI5XMyBR+Nvcx98c/zyF3GlRqDNVV8JLf6PQdJo/KGLBC6UXGw3qL4tq9FHs3nw2D3D
scZkRhExXlRJxpm4X8oKP/chifpAG3ipNjM79VDxfHohijvG0Uz4XO+r/hPK5fPQm/7m8TjBKBgb
qyvEGUB3joQnatUXJ9EzmHq7rVjJHi+2JW96kMxQAwxLK0O8l0h3XhUqQe6h6SRg9Mbz2VTTVApr
KZ/pArTD1pDnRyDodLlF4XfTeLEEKHbEGdsEo1SFkOWdKlSi0+qUgZTB2t7gH51PCI3BygceRZbs
x4irIGPSxpzRjphtOtsVFHFAZqVjyejL3rhAgp/RKrXRT4h5J0JiErY6f8qcah7+ecEp5VZB3a7+
QDY7GF8EDrqZoKyuuSboeE1PCzTMZfuYUBpboQZrlUgJdV+ZFIL6QT0bVvA8Y032z8H6EUqNVvQQ
yRn/erg2/d3DTizf2FbBg8vkf6mwx11s0oS91/kWGLgcqMhCC18hL6M+3noav+BtyyC2RpJ5YJtU
XKh32pJZESgVoIJUy3XWn1JlakH4K1PCOTdgN1P0P3vr/PhqguMoPXDlwdUlTaYrN/434zdlPeuU
HDy37UprXEKNOBRXVdKzhBAl7At+evuQL4mcMVXPgebaMYsWJAv/UOTfs/hbL6cJSa+GeCYDXRUo
MTxexN7F3yoBGw8zdNf/EZgl49lvuA1FDqCnsD+/ZT99AC/XWRrfjlvHWfpcF/8XU9Jmo+rgJSDO
d32XitVbtQQI2bE10cnnxxmJuTFkNKDcW6wLnpgDpTmoftfZB0Cl3GS0VBG8Gy9zxE4wwneiwkHH
Wy1qctKcl3vlBAG+Rjw8Mq+c0v/0xDKTEjeJylLHVgAS/SdchlyQJEwnkIez2Yr1gzXO7mDy3QcI
CQchlrDQlgZCGbCA/5KpRrjNTHnRKwP8yXeVuME25LqMIJMnXuum1n5VX+OkjKKYvyh1msDbOWXH
SobHiIfokGyawidd9xAk++6EX1+5qNyFtGPNgPNGdVaBYA4molGMKNxAN6Rk+jMlPVePrmZqJLl0
AQgStO5BQ63yFo04CPOO0N297zjMECsqRK89iqS6deXtRaJ4a4B98nET9M0uUQPNPIn+BEit4vny
Cd6cBiuqZiXe4X3AYXZS5tQ9g2TTwisr+si8OmXqq0aPcD8ZBUuWoKHqGY0cdv+4TtXzfdHY6LqR
/RPi2fDElDgO68Z4ORyX+8MHIJiwc9AOpZRMcN+RIyGt3UPEScsz/8Fk8FJCmSPO7mcy/q8MtBYr
XvpTtrr5AYuUICUu+hLK/Rn1Jkoc1k4XgD71mAmpbUIz5p4I5R0RBvhbHulJYZVOu50GLqHZoFNI
pwLOeanQOTMEcoMq0shFdvNxDoXiGSDdcbLIqjGAS2jo1Tmb6bsDj5vMSWLNU09kAmuZzXNbwvj5
CkPtHvuyu7GTufDp6xwVQbQBCCAYminlBmH+2rXOxE5qJloTyWbhb4GmU+cXPKwaaz2VWyHj1OEX
6ejnGdglS6QDWsr/EY1E/CXwnxncYIpELhMYuIpJY4A6rCxd7SiQdoJQAqawvj2w0GDriSUHWokk
kim5rIzPUX03vJ7Jld+Zxig5rfFF3o6rqdhcsHIUw7FTDuFh+d/nqJI3eV70A+/vmQbfTXMcwFUl
v6UdSnyCXqrSxxHxYSL+dTdTYpDwXX79ELvzTZZ+t28JhWgjWSG4E4WDUbv4Zgt6gymxZWkcuKyl
E+mlSMGIdv+Dy/NR0yZty3wT1brfoFllTMU38Cr3fSqsYW+s9GMoc0OCgzxDaXPvMEpuQEhUuRoq
PeqMDbCr3jtmfVdtzGTh5OQq6FatJ1WHDYujtvL+zhhlRZuY7LLBgNur8txCxv8SfS4A54WfL6Ox
R1NJtS7JDK48QiGWfkvqtbXpCYR0fhyg6hWVVwqaQ2SJc2qKwcBRXJzV75GK8fBZhTOGjyTrvhR7
ZtKkv2M7rPPDAexEU8PwQZQpi89LPnTzlYeXVE2hq9M2VZNpgNdiDTDdc1DGjNtxi4FFhnAsegLx
r0ue9zfN7c9r8hrjaUyMbc3dAL/1Ug+uc9G6MQybruVAhdlcqT+N9h8gJrCnyD4+Wc2P7fMX35cx
hFlFpPOR6Tqr0ldB3VQQp7ehlDGDJqoAMORywSAMI6RLvSu3BIo6wuk+r9J/0pGu4nGiYUPN+/GH
+jjR1ZkDsWZ1iyx8kuHVdaLX4DYJ45wsoIk0YNvh7kxHTLZ2fhEcb6Ru5CHEP5QJKLiEfU5g7fni
Yj6/HF1JMnNBWKI5YCGayyng0v7Mxn5nCsJxwB6rsMDpwyru/yP3RXZuzj+BTeRET0Pqz2U3y+/q
HjEcAq98SggVqCkY0dGXccafealOW41I+Bkn94EyIlT4kXoUpQ8CtRujYXABYIomjz+9p5e+OHGr
q216CFdp9WzhQCLAYqsxTFPJwlDVcN2ULCMMCj4fodByd/bXPeme0JnFxjqpATIgkARxRF7Se5Rz
Tt0KP7ZpY0W1SXZN/QX/X71sL0frEbE148Tx3jmTL+vzccqno1XNL6Zp8iI0ALUQ+p5B567s8q+i
JpdrWVZ24JBQVpFg0RcvEz9gR380DHKXT7fSLKueYIoiZNJo7vK3HgWigLHLHsXg0fOhJSDYYFXk
ApW/ehDYfO4qQ4n2Iztx5F7HuiVpNFrWrw9ENuySRpJ0Il8QtM4VCN71Z8Me1zQNj0Ytb4UvquaZ
6PVPhVZrvQPq+uPSZxMd6fJkkzL+O85/ybxfIMw0wgrp26yEnG722iXyYNmb1nhuawRzlpIp8n1H
8RPv1qYZDQNXCE2LzXD5pQBMK/sItWPcMveqhGKErEMnpCrjaiJOmX2q7WWivYezMpSARNuH4RCQ
qWtevTzmTnTdDWNPx8GJD27ND5uGHliK3nZMbVU6V0txr+t0qo1W3UG2yGTkaRX+pMb/MzSP5GsY
mYkF0RjgF4JrHxvhsnEi1lvmLCKA1H2ZL4vi5Y3ngpwNSlaLNDw8MUJNQapc1q2k4CrjZiOev6jc
mTUSKe4AC7bOzED+iXBjHtmhxAusA6YVxBiMMFTQxYmIC8ahNQO5ir2k5bnsS83Znlw84brFqZCr
/G0gKN3zYJd/gYiZDh02IX4tiTzXWazeO0EUwg8hb57hdg5m/fPP/O9UHYPsAnaev0XhX+8AG8Z7
Xdtkx8r0E79xuE+hYRjNXPgL08uwFUbgo647uspaOBPJQIOK72BWP28VnjLGhqjCBzR89s+R4CD7
+CS5keMgWphVh/8EdQApcPmMsphya7vWdjvnInlyJCkf3U5oNuWm55JnSgTCmvxZSwScE1RqfYPP
RXyX6f1Kvgbor0RN/zjrEE2RaGNDlCBIxsIpkxUEhl4w9HYFYe8LkEtrYUV5eqBEIeulK2mm4cVd
SQH/RcUkVNpC2uETRyu5loXF7ITaKFVKOCOYuJZhZ7XnIFtv0GxdgGZ0MXp2Yz4BYYtozuMIH2pi
W43jqoNYYYq8x9r2WmH+ayhL2F2J1Wj/jw4ew+X8J0G3zVXfYmQ4avzDZBSusCnKErULtOEvCzI2
Rnd61dXgQ5Vj7B4XzWxQ6O0xB8y9LeMKbr78tIocDhVCvuX/lU8Y+LLpwLxkdbk6oJkTLYw1nE52
sZK0tNrJgs8GGkTGLnPPn7NWxyz3SXUSABI/2zco3VHNiZxnRiJs5tONSLr4U0hRnErkKhQhCVSW
yyIYrZayVvFOpUSmpmBtVsIhgd/EQJd2DqnYKbXBrOuiGykZJsTF/hmMeS9rpCqOApb9f4HeEJ+E
RDlxfcHxfYJK/5vjLi7VAKtGy+5mKPKGtX2zIopH95MNh4T3mUKlVGsdnwW18uS7YCcybQMUlQWn
mIZJo/+f/2Nw2OjR4T5+Q+meHA8dg0NoJ3dmjrKUIKHiquLZrQ4jccmUM+xlCwo2SYurNNhnAVhZ
E2WJ1PwET9CtC/f5sMoDh+hClZhKmHdC+uNbu6U0n5e9G05SYmo/gwp4dBJ1u9RhaLC86dCMtHkg
2fadrIsw2gsert6ybyA5f/z81USHFDDHVjIpjMBRaWLT7s2SEMOoK5P9EBXAQuiEcVUPfYZnV0WT
/5X75qSOuZeqwbO+NAzSV1bFMUqi+M2uWC6naWkrXUbZVnOiZRqsonJDdx5f4/UOPxRVi6ntBbwd
kobGUku7W4JHfHW5hOG4qe6GtN6xTPF3wt8/Kay79Aj+Abv586hK8UcXZNVLi3yb1Shb3z/VUb8Q
XTlI1/zgcGA07wNRxhzi05QNbrlVvhu3L59Y+wpdi04UVfLYgfPGispAQnaXMDElXAVYqqSWghxa
RE+fAlYTkXjdMuHRQ4PKtUsztLG8VRQ/SaKsd6YiAshJ7UFXXxswGkpy2H1Smvnwtro3ZDAfE+y8
Tb3NSbOB2S1Ewkx7Fihfn1huHqE+/82+gctM0F1yGUzg+X9cAOlb+Nejew97C4IXkMldHg9b/5eI
X9aYhBpOoKyQZ7h1A8oVPhaRL9fEGVL3c4V76gOmh/NEHCrRvBnIAk0ilzXjGjGWvmxA6XuBXsdr
+oEmPyxziUH+PkLvFD8HTjwNPGygUqC7N9nM7c1E4d2SC4ZKOYECiEIA5m3V8alcrNgxjXNY+dTX
KEIBTMi9/yR2bf/rRgh2pJ9322ElOi3a7IiCgT7Sip0vrJJSChrpVoXOLAj5qVLqbL0uG4kaOqbU
f+4p6BbKEdkNxmahm+zR9jAoAnek4RoImUPq3mGZCZnDhJ6MXvg581xuVbGeg6IkmtZMMBY3v/DK
g7665bG4HX+yd0P9d4T/UokoHM+tnWWvnDSjfGO5mcHuFEd/d7wukEA+EnGBRNI1JHFbFtIdT6G9
MfwE5PiFiRTQjYPhhxMZ13ImaP4ewZdoemYY5sfrRxBiS1QMc7/BlyoI7WvVLZ6QZM4lzWbc6HP7
TRWtsO7K3HRObZRB9Pbh3o0XLpadwABP+kJVKBgOEzyBY7GURa0KeS2r86HoDCzRic5kL2J4gK5D
PPCF0dK3awxjsBZTOraLpeoSU4zXTYI/8uymamJ8EizFDN4SQAUuKxRTzjCwLDwtPHDksTpyVHt2
mHQNVAd87VYdzV+bv3XPzJdYxzL0EREeA50DGkL4+pWFOChi6lKhf8Vo91q3oS7cEi8L+zyyRci8
MfX9XX9sOskw1S2JNaXOtu3treENhV783IG7v8UJAK89Yr7D3wc6Jt0i/lvNXsHs/4rjhkGY+b8N
1otFprV4XCBexFxqxsFHslxBwijPn5E4Pi5ifHSuiUjD7SPPqkrw/8oFUMJ9LhjCbKkS+Sb3Lj9j
jGxJ6B4oKeCHvQsDaIR9WEqu2fZY7H2SEn63oh/vxW7os6Tceq+HqSBIjPbK3KYuW/XWIEBwE5Fm
PkXwnbD1GIYtCRdn5UMFGkFUEkSsdj5Ih3FebPrbb37UCeGPWdEfO8OdX7XPtroOG/cpfur9gBKT
+oF7vS0FjCgDbSC/wXML3AXgKZTg3ctVjrOwkcZUJBxtQYkwyxP7WtMj944Nj7alO1lb+rbiFXkd
ozv4bbQSikx9OAActjra8I6LPEaaY8ppehyLAKrFWBDYox+OGZUolKSfVLUxWQ/s0P4d3NKsnWnq
rrWBaixbFaZGVpT6EmhP9/RBIW2AyOSEsEZlQx71odxHNj02kk4urgn0k9XW/9LcCL0CHIiekn+r
70Iar9qbRublfErXTaQnI0Vu1UbEGFyU67arTr/YQnpgXEiQh6jp++DuC7YTem++XFGYJFZlVJYN
cxh6zwa+7YVRdKJN+6MZEFB3Hwlxb0Vrd7+WNPu8tpjNHDXjJLwUSNwRg3zIn0Hl7jpMqYcXUn3w
wSjjshliA2iCPQOP3eFyP2R3IszlX/67uPfLkfCVSfYxA4QW/uev+5d0oy2TI8/qmqhA43bzA3FW
WVmqgWwX7WBPASa2DwPwLEaCF7Lms23ttNAtm0Gvmwu94k59FV/BG8T0HVnfNnfMT/6mx9p3ek0f
0BxeMExdw1hmrZg4YFj8D4ybWOEIScvPQanroyV5q30DiKCsREdn2EfiogVKMnWee3O6a1uhlbGj
EcY24DTD8j9I3aM7RcyyUtKwflZY7HTVUf56JEXYIS5e8ENhFaZeeBc6az6P8/Kt7UVATZHuFL4r
P2DVpQbZcIarCU45z+QEhBTXjYL341uov3bLKa2iBNNKM4IbE2/4Yb9leofGwtNj2r6VXk+RvnTh
KdUK6O3irSWdaG5eTWCMnEl935HnDc/UwKq4bHA7DUW3iylEe5FVeKoqQBT+67/Q2Q6ZnU+odzMk
uFeGSV7N87IrTvYZy/SDJBuOCybZ9tfl6S6Mr5z4dGFf2gUQLdiQzlSczHhl5LvrwGxRul3ORIxa
ZecYrnE7WuRjM/whHH/gDVcyMTWbG8nXzwQUqIMjfsNr5lqv0KcL/P0EaElZrD0Md9gZjN+cPGuY
CLzEarW4Tlmy1g9WsTID3RJOBSBi5I4JPzKuT/uDboBjmMNp3hGf77f/3LiYI6eAdD+CJ721lImh
oNbi3n+GdBGLnKQZo6215yu78174cURz7AHisc5ViXzBRR/eNHx+QH3d9Fm70Fkx0jUXcNEch/c8
puUHRMADpcMWtss5Ym9F+23UT0W5s5LXJNSNszLNzssiFmeW00KrIGwky2HEpyhcMfdos0KFyS93
B5Fy3ay01z4DARDsVn0YOOno2WFt4IZv5xGWwmSmhTcdRqvQI8ejp0xKVcUvl570fvpIlYdWgMMg
qPRpdviVElud2LtGkDAmOhO+dOa9bqPHSsnHobPkzkQjuVB4mjPtmTLHesIuSSAPz12yJdZqRRuG
kxscF5sbDU8HdsdWTEuoaTbvAzLuiMD8GmeSvLcMfOZd/Oe5ZvfQaGpW/JrBVPD5I/SMpDDm1hzP
Wv2C3v+8EqFtWJorbQuYGhmpnEzvmFw1JHe03wCItduulWsrwmfT2GRChRuLa2dKw37EqnR2nfij
qRmAK/YDSfgndmgBTi6T7Sfb39T9m0DVSlcCyE9qPYD4mqyLSeQjCADwi6jkdizDyzH4WsXYCAp/
LCBiGRdF0DghO2Nx6UGkPuTmVEAyedaU+gf7iSI3i2fFY+Q4KJp8PLrcHiWT4DsDdt6vwQsCTODG
HpYJ8LZMIP/IO2FEjJtYtRW1m2niNXqbcflA/GBpq5OvnL5Rc8/Rwmtk/TpxbwEB2RErXiuaFcGq
KdTT/CUnHhvPf89zTVyt2jS056suI+xWFNOst9MusBJQ9pFfAh8V+jU5hduMpu4tJTHWsZ5v5IVQ
4cRP+qCikjAWfgTv5DtKlDQ6PiFJ8mogPNI/C4/k9aRKx6czFA44bBWYFAe+E605dj5ztKTHmK1v
PHEuRoV6L9/6gTbVjXPkkM/H1sCZLvqKJhQv2p2HDYW3Yya02biSU+Zp7zwhwUOOMnFu3PPeOi2u
/koh2Ec2GejnE5AnXKoKIGSot/thqLKhi096gGD2EC9itk87Ro9ftmYtDBlTwF7bkFhH7RJXrF7t
KmYEDXYLpbbpd2XrTGyDPZY1ncnfia0SQodZDbl10Ft/hDU1UPgEWxyRUmlnwZwAOB4m5PR2R+Yd
LzS8KQn5Hluy840II8Xw3WqYOwMeh+efO/4rhqCF/s2Pas5VMIXDpHyzezQYnchgdJtGueZ3xjjx
eV6FiEVkDekaCPnEKg0DDNi1DISx070vlJXdSNS50onkcoojGKPh960OgPqB0AYveoWpBBfA0wv5
Zo+6s5Gqsl0r2BmHs5r2ppswcoDNLtsTG3rCTSN3mHDN37Iyexne1uzQwhVLtQmES5yQArqYTq5T
w1w9zKMU7owkf9EAYXalXjAy53EhkC8EP6zi9byzOeARgfouA2DNvsPKlaemcJOpraSi8S4sHhRx
vSmXZW7f+hp+3oSyFvqUUE2VFGrN2zOfca3NOFTP/WIGRb9wV0bDKl/BjBFgG4rz4e8jhpjoAFwV
TPxwxdSoqAoee5EM94b/kbmC/6MSXMy9Aa/yMfGO/tB0O5GPpOEwcz2qFdkjaFAJbMHnXgcdotjh
VzOnH/lbIQ16VJXP8eddsGN8ZKAtaUVCQuMzUDbYp88tDbLzU6I64kZ3qx+613NJlhohCtjyIYtV
3BAwQavuDPwNTollecD3y2LZmoCvvZ8me+YRl+Y40FR60Pk6Xyp4aVZwx+3qSxM7FNlMC1d/dChl
qfLX9TCbrFo4m6CwYRAYUM1QwaQ8qFe0SIzkLtaBYH+pPCkV4umq0mDSJ0yr+3GGuQu5u+m96QSu
3df1Ar9BE2y1MwsgonB/IV6tjB+dDXh01mu+e4oALNDOyP27idnow4wC74Wf7eAbaBFEJicXdE7n
Vz0M4rowXM4svtjO/GTd1QxuSjAFfg728lkuSW+A9yp51hVSHO9bAPVKmXjlxmTDy8lr54ttgHwx
2qvveY3plT1v7GzWHtv7FqNadIu8iZvMomXJDFc0LP0/fZNRAH3QoBuwkMghuxNMEDN/FO1o2XVX
IugwzFVAs7i6JzbnAlcW0d8lHc6GhjIeEJEZ4kZ1hvtSo+TDQaadovqmLIrZP6NKW6AO/W8MjVAs
Oc382wTOpRqIGgefCkEPrEwTM9sdGhl1lR5/karEaOAioDgNBSyk8CD7pwx6zfVSuo5Vf3KS1wDr
+H6ZqD9pj6Vmtg+qkopp1d8U4BpYJiopRgkzY4jk0xlbWfE4PN84s9XaxXM7zE4ydYTqWhD5vnJT
st8qWY8N+laK/af9fu0eNgC4EMJJN5Smg2o2B2KhRYlSTu5EMwJH+mWVT9RQA1CyA0aOOH76X8uI
Uh9GKTvlXOhow3nVQ7YB9rQ4bi6WgfWNuFiH2LWFL+LKFLgoBI9iPaN4Ro6122BeMz8t6jbdS4BA
39Xc39n9Td7jBIZ1MeAsy9OwuVNIWp94RA8+B67e1BHqcy4uBy8DbCEoESDOiFUay3UgBKi51bUe
q+ULx7xQdjtbs48VPXTYVVJ25TRiALibxFE9x1THnjem6Ep9SeUy4lScUNrf/Bb8PPLIJUQNQS3R
hNEl/rajVfH43sk/IErIloSNIQqz1F+oP0+xhLQ3iy2SHLSe6WnS+lFGZISQRGlmjFF1JXPM4Zra
XdGA+Sy4jshMHw0rWffUYLYImvO7gYfUqHJjg9ePyMWF45sdJv87xdilSSdgwtwTd8nw5TOJL5T5
nnqx1+kR52lTV9Gz2UkrErIfNRS6I37unsVn1bqheddJ/rQ+zkK9Y3SkkoRw9MNHxImWy8yhT46P
QticUpZoatm8/bREAsMezosmfGzI9qrNYgNkdshP6vsE5M8J44wInNaOPjGUObO8wrEpYpVpN7u5
v/Sau/d0EcVhKcvMGzruAyFQWjEOepUjdX/eSVYm3NHmpS6qpfbS/70f4PQqhUIjcKBRZIxBiCqk
11f6xV8HopzA67QnzfboePDpTyhcgHnuh9ILqGFmGoPwQx1X4atsZEuxAwx9TFrj/lqdVYRJLpJb
8fju0mi488Ei/n4jICvzYxiQiMjb/kQszXg4Enuz0GvpOLlweDZyyzrWCLwO+u+YCh9AFsAuKY/t
Sx1fVEb4IShHlUBB5w391EADE9ikYpcO1gAobl7BFqwNh01uHmG2xsUT6GToKj3KmqpyGsuuUVxN
+t3CeEPhQpwPKeT/C0HqDD8SIqy6mWHlZwmPFg5blOGhgO1XSYYvaJCLyZjsiotdMP75EP546Oyu
KPfqHOHVo0jXZbkydmoPjTFneMQXVHFV3ltjtBp/yYha8JLv7VJEEckgIaX1ek4B/o1SHbVZMJIA
PQUBRLkyLTky4NhnbCkOtHKe9Df/2/82odWW+f8AJ1W1c5zkEKpAcrRRPzRJgxIXLjImBaGeowno
6ZTJCk/EOqzQqGhNImUX2UKvRV4MhW+bIrAdU5iMEK97/fajvpVa9rw6U0/zZvMT93ZR42fh2+vD
YZJC+ZysBD64kyojDNcrP/oGGHssKIH2iaDX6tQ3HPcMxQLnxVwxAXvf6aYeHLLFWv6HJKbbJuy3
8HT7qHVKw7ADeUZqaCt3ZysQWJnuCDUB5hfH+VgFu2Z1MaIi8Kca68pzeSYjlxmKqycGX8NH+IsL
JAH36TJ/yDgyM1aUu57UqJyQ9pE5rKA+Hwx95SrU7sENhpp30lOBFAO4jHWmSoHywCyKcyTgu0VR
VVWsCPAzjGxs/V2GuzInZlwFung4E9NffPrUn+kWxHyi6UdMwsb3cvsOCy9q1NZJI4Gf09KxItiI
xLoNBKDetpCeQlBy5yW/HmpKuekDj3eyAezF2wPR3/eNmecyOSFuDkox7zKwRYtLEeRxaYY8tzdM
EDpWvk6zwetN+igzTmUty84VBrrEDy8XAiR4bS1b0HpMghfus8kJi2bX15a5pydLp3dWT/Ds6i41
WtnjJy0fuMST09lzAOoM4k0pHBSq9ocelVjYKR9fTRFD3ABvnoG+LHQAE82/E2U3iQ9UvxKUsXls
Pe+6V3lw1Epol3TAh/Izoj+3USlch0/5PsIXiW07FpNPKGOLzQmca0zYoimX+mkSN2wXb/v3/Y30
if74QypCYKZIA/Udu2X41/FnbkcvVfWcNLcnAVVEyGSipABOdvyeqnhU1jGmCED8Ds1gaOi5Rlm9
FXaD5xkwJvjv/yxN6svjW2nHKEvJy8XfCQRaGkE2BCidvYxcgojknmG9zn7MFxuqWQUoc4Bf89jf
p3AleRfv4S5ByeQfVBqfRuiiF3J9RRQXBsCf9TsxFJrh0lbZ643w3TWzyiWG1tTZpCMaahDRnpKz
N30D7j1KVERevY7h/Ji+i5LH5i0fZhNF53qb642SZZhQ1Fkbwc/llZovKX/yAhC6Qz1SodjO79FR
ri4m6i7zHWJ78hKNyuShfveSmtIeV8jR5uDQtBtRGtVEyQtj0wP6EtkEFf4sffZcWHV7DB4KMgmz
KRmGcNRRILN9/1ULKDw+P4y97VpF3bRHurzgeq3Uzzmy6o8PHDqx+yJKSpw7k+TSNSaCjL+ZxTOs
eBkWRE0WT2rKC0msYQnnJSVWWgcB3idSjGGacNxNyCTJM38wwKjRGjd20iiq639kDc8wo0YL0cLm
dc3uTS0AaOr4jwCK7XVGvop+2AS+unCryoa2ZffIDN5urEM+GOfSlcQNfUJDoDmLyoJJL+NkJjnR
qQSyFfa8JXaObb8kSA/7Sc7oo76LBBJZbpo25SHcbHIuXpb/XjlEusa/Buo1PgsFBUzovjCvbPt+
6A+afZtTSltKhsQhnW4KzdH6phhRRoFIUtW3stdE1I3RS8uezILh1jZVTVrKHNhaEmbIo8H97U11
yDZwPjdW6Vcn/d6C8s7mXIap/poHFNqGOr7iVNNtyHh6kyBKQGE1UkjrOXb5RlzjJFIaPwxriE6R
WH8y0hqPj69EonLCC/NklO0oMiz+adNuDZkrr+zzyjXBV0Sicrgi3VAJADNxc5QsQ3q8Du0KVSZn
sWVysiy6ryJMMxzDjLrS46UMfaGz1LkXuXhuzOEEJSgxp2B4p+CCOxLECmrxzLcfCCD5umgLQkiP
GcHrcp701FXtbGU3K067iZQZmh+XvQ63nGvCUYpIPdCUIDy47wW7K2mW/MNCMgESp1z2wRFtZlET
fgoiPArlOLnB73vIpima0l5Hv5/EchKapanWyWmtalUzvc7wI3ZQcaGpHNSRWXw4qVMHpYPlHbZi
cnASDn/NLCH8VdIwkIDNqoGoJVfIyeMqhLJo6T7M39VUvguocQLoYTIUjFfyX9ueTX9Sf281xjFJ
rhXBTkNv8oZqsVUe7g23v7e10gZ49+YdQcPRvum2iFsp94RSMQY7g52+j4ePmXjUjv/CYyVUb06r
HgvCKWvw42EpUlVU6QSsnoVPmsdK9y3EjZ4oPU8SXWtrbB/V3WAwG7OMLCzciefPAopkk/cJFls+
1BW9CeECwBJvuhyVY0fty8PczWZ64x2ZfXXbpKqefRdHNnjISOg5NS+gm761i8NReCYk228T65oX
IH6/j7ibwDJ9Rofd2x4/AEUF2p95At2rssOUCqG6EW3eyESah6Fpv9I37HA6IeMgBFclt8S0djoV
o/uOgwN0l00FRzbAf9rY4zOv4JM3pJWCUoJRDPLNidRAjyFLvthqxjqnsNzGJv+bMCWCig+vJ2Zj
2zORjMRqzVJdk+BAG4SL6cmXg39DKW2uSva9P5Od2U6ontuc/gy32itlEysAB6KM0nxWTWj2FXAk
Xvxbml5+GKSLH93Xx1MhqRoRYO9u1Km0UpnJTK4j5/5pf5nu7XXzl3cCnOAzFt75dZMd/GMrquze
0BaEQvmj4SYq1E9DKkQSXju87bAfyV/o/+5HexgFMlKmCtqKTb6U5SANJMXeS1QnKKjhTX67HPDz
FtvA1tsXnYvKMiKfFAm5ylLuycnh/d48FLZKgCHdbFXAIO9nX5sNzzeRakJ1zw79929ffAlCe7Gx
9GvWGoOyGoNQqA+iMPZGKg1KGnnzqoGigIV7/oHGprYPJguT9gyLBs8k2Az6fpMboB/obTQKbZoL
wpbUhiQEsA4UE3Hwj17Lk8vnbVleKeB9XZvKZg99xqIadD2qbuEJZsmgRL7RE45K6O4QxTpOwmt6
A+qpnCJ0p4bb7H5Ptpf5MFeD1ObccVyKB06v/o0m+4MlM29/AIWRzwhdv7m9HYjakySLFBHM9PKb
lgTV8ah1Fxr62c7BJGikSKeCtjvR9qVKY4RLA2GXdk3+S6g8suZ0QA+VG25C0OmN62juOEyzb4oF
ctYMz0i1fyBOiXMyeV5GGG+6qSRUjkLbAWY/0pDkDiEi6t1IUu1+MAWnauHGZxfuvbu3XffnYFnW
497wwCgUWqOyN83eDLp2i3UEor0pApqc/DyIrfrzd73N6sFtFkzgVfxRldbUlOtoc0l7r3cpEhm5
dnYtZI0P7IR+q0a9cS4yhfrsfKnUt3Q00UwAYN2XkfaHRHTqjULbDt+P62Wb0GyWm+9tL9x2chaX
+rHfLWDlbzoQNPBaJnx31BJKEt1+YL3SSKC6FESQ0mRXZn52KiBq9xlgrI+DGifJCAiZOKO25Wal
VRVYOBnHdQFFduFLysxUyjZMR6T8MwTpl+t2QtIAC/IyiGY21V+6VmgkkwlT5Ri3qlaFCZM1ilEJ
EjJXloV/E2Rv1+LlZaJYNNKPo0h28m23SQuPMplpyJUP4qBr19VzrxHUFoSdAmi/qevBoGZX0HQB
XzaT/s+yKfkxgGxI5lm7ofdGuwY2cPGDzT1PCPYIIzovap9tkl+5XU/ZC8tU5pkFxxaseQjh3Doe
ZeVT3tGHJi5aA6Z+f7sIG63slq3zeteR5pV60S+882GLE6lqHSaZ7IqPcqWbFcJPQT1lUsOxxMMT
R2DbMJ6Lthkovu4Gt4e3PaptVUzpITcmFpyOIEEp7aGMcMD8P7HC2uerSPr2NmHd97r7iGzHNb2V
z3f4elIyyiN3wNEDSr06ZJDU4RS28LQYfmNBDZ97JcRhkQL6vsGqZHee4GmPqBFM+o2RC4EMw1RK
s/ViSDt0qlxzYQTHtqd3KN7yRI/3LUpOzZPrHf+D50G3E5fR3XQbu95ATPBXQQPa6YUqNVApMNgF
U7PjI2lQ9s5Rz4IhFes4Baf8hNxoIwqiJMisbjnB9V4etRhVQ+N/jf5En8gCq0w3mR8uJjOm1ZJV
eg7fqJ1Xr0edohcN47NB0huR++ADoOfU1pbZIoHo6FnMNRUPMy3DOwyQ4FhLyElUZ0bJfCPzuHjH
eVc7pRJ7c3ZzyhYSddGb1dtm52iI5DO4V5fNQ6Yw3onVb1TZ+8y2Z0IwENOiAjECG2jfolDKrlRi
pwzcsQ74hg+Ha08f/618c9Kzr3AShZAfwuEqabSuYyrgTe4eEvAl7hgPqdBJl/PLRiwFdqBZPxFb
/09U6z7VQ3F3QyG8Q5AJIqmP/SZdE9jYl+E41zMA4ilW2F0QTBVvWvLZCaow0ELZe64ASGk4epBc
I4KGi5qV78zntm10HI1k9tnnLh3A+ANaF+PZuf0XLfhWAkPAPaOZco/MCghuu6MzfqcvKTaVQfOc
6zmNPQtkMGT/f0zhT5bDet+urYQUaEbiyWAmRjgpoJ7kqJT5bcW917Dlcb1AomsHGs9JjJE+caCE
UljJMroSA5DE0ZRoXgr50J0Hbj4XTrxyWbwU7c6VqwiqtynayTNDbpSMZFwq5uDlH9W/u8kg9wkM
WPR7rJilqhquwhKYYhbibLuBKWRFe9Jcjrk+W0uViiQhta9Crfa6e6NzOYxbOD3zNyUvcRIb4s73
vU+Le7180dM3w16Mb+z+l8YNfM6kdBgxqJOwTU3nmQu0xMfg9MG1LBuY4otcZ3rIJMEUvKEYdNUC
wuGZXF9wIhPZJ1VdVC2Lwi89h9WUOufIejjSXXkYGPz7mxV5V2tT0Sjk/v97W1YVHNkiDr7uzvi3
/aeLnt1G6RQa14wMTzZ4OwLAaszQynm5SmxUBh5vdTBM/0cX+O+fJdJOOhDiTZcG9G43wapw1KC1
dRCqGYlmd3V+eFMNj/jQsaLa3zmrJVPuTCiuWfkut17y1F6nMx6ltclf7QtG29Q9auYq1z/snLkf
8YLCIuOa9mV83iyEF+LI5TdZkADM7sZOxl57xdwB47QLT5CArPJkWTNw5duzNIhwJFmSMl3u8C4f
3QqyfDx/Ev9kxeqDJZhkPJcXUP6uB/SnU03O7akRIgsUlyKrKJ2O2C5+IBPF25eJUg/noo0EN5Us
EfuaqAWGDydPhEN4lBXaYZUyxB3OwEiwoN/AA+xd20OSxspUGTrzYKVRFPsW+EJaoFoFTntP1pJy
5gJNauXXkscp6KHqlniUX0/nt3oKFSwXvMYweD7WEyFSSWXNhECGIcI4txLrckcssTbHyFTyWIsS
QXMKooN4eBJUg71+UGZmKK4Wz6HUy9D+ipaprpL0wIunvdCgvTDBtA9kprVVaEnJDRH1J0YuIkJW
bVmrjGepROwb92zGxSeOfTmJDhOd71q9GgD8kniCWU/BN9x4+XHABYRuMUbXneXdFFFtrRMD8b/b
P/+54gKXMzNCsZLLcCuV61FahPjuB9TnLHUvpd1bUHu/o+6p+YgQf87Yhr0+rxYa08gkgn4K0UiM
6/98rj5M1Y7rEXlPVGorPhfZtXrNTRgqDdPbDm5taLbQQ+BhGnVFgGlSBdCMrESgES6JHKOFEXDh
0mtl9gTK5mMCayVyae3ug2EKzzO3GiWsMgUSILNSTDyez2Yf5RwBrE4sGysRlxUT53uWtT5J3jOP
CK2DxzK3aBhs0yzHv3sNdYEjLa73/gFtwl9Iq1BIs3wGov/UH+A0r9zO2XiUsOLeL2xPK9GRDcbh
io/xkP6TfXjIY4XE4r9qEFwKExzGZOCN1T+k5oAFSgFRzeZ/7ex2G4rJf7qUMWgPoHbAvxwaj28l
l9VcNQVxPjTO3aXU7phJosBP8A6MLLusneZXoLazSgZPecNfFiUUzOsv4bR1ZzmyIRkvxzGE92Io
FfR8NpatUhLT0pvkAdNJ7neBtKDOmHBmxY1rt5gP5eoJqtVugfI4wwyqpSzH501zmnSRz2n/LozG
9j2eI1fxA0H5rlU3XJr1s9AIKwRow9pvIlyVpb1h6+/k+7317Z8wEPlBz+5FjRzXQS+HHAOKCH1U
xC+XRJx7fMTv1uJK7DJhOIgriQI04jVf52NvFS7J9mt5fxaL/TxjYvaB+tfMzX0L2PVRa14V6v/U
OVcsY0FIWJoRERKEtprR6ffX/UMpTZb4zbB6nzrRvMTsd2uKdIEKmFkU1uZmPKRpTFs2aEsrmbaU
XH1g4Ya0CG/FQUEphrVdMYitO67JWM0dICS3sx1OcxX9socghTOjLThb+81HDkVNr7ZzVIdMFI/W
BTgM2py/8aYVzAMm54R322IhFwUHGkBdGA29LiAZpTYosSsgAlC5X1IGe0pEjQXwKW0uNLYONovw
tDyRqCK9pYXpbI8qxTi8sqOs58mB7Jc9MX0VwXeyDxBFNuUkmjcW1u4zNH412zNsDMa4T0j+ng40
wDVcwGXb01V0J/voKH54BRNbs9m7WeTGmsL+cE/Re1xa7Yv+5X6Z4LVhrMeuNjWid5yCnhebRKTx
v1rGsyHVQkZaLHtavAoSKNn3okkAwU/UbvYqoj9zwgtDvOdsU8eW2Luu4D3W24HXG21HXhI/xsHW
c64CNZ6mp4vxvZHJs2xFzAf8k3g9w/66DyBG+hoX+kbr7RINanLqXInwn7Hflq1SSWY1eMR8Nab7
RnU+tnMR0gwnoXGuH6NzpzLYiMOgmU53PNiIY1sWe24+m1Jl0hVKKoLNv6nUcJnHhvfoUT2gcQIW
I5Ac5aHXk7Ge/W4iZnP1AmOUs4IMSQPHWJcEtVgCPTWtagpGsTn1T1Ise4k33DhIDbT4Gx0RLJzp
npAVCUuqVAypOkgj8P0Ikhm4LqFqelTy7e+lw4mTFJsUxzlHSXF4l6Sn/i8b3CFrk8HWMrCZ6jIy
heRfcGVQ3IqDy62ms44whabty0/q9AZl7nJ4/M2eNDTMToiEvLTrivqzCqTAYCQ59N9eTiqi2l+b
IcUvakIL8SlT9M//TGhI2fRHOqnvS1UboeQxGXBgFqZ9C2NaBCMvbmTHOhBgXnicZS6AS+8LK8sj
bKxfVX3vE3CETLuM+BVul8nR5D8syBYXpJ+xQael/d+IEud+bj1thyvpfW4FFDrtmFcvGuVLctEy
G2T1mg6+FQOff/CYafb2KnY5kCSRtS8ieInKaANGulLWI8iHkKAAAlYHnXF8HB9BMwenucSWw2oY
QK7AKJg/c0BtA9uJNfzkbHhKpH5fr4FwpNP2TJMYRGWBIpzJC02MuhN0GT1972Q0OEQExRjujnos
i4grae+QvlCGAjvL0UJgOyZszex1MeEYHrCLI/ddAwwjw0p6tYYqqS1R+pdJn3PVsCTeeATaV1EB
PCuR9/4xV35RCdLjfexrbcg+OcIej7Y/I5RHve5AU9mw/utSwZlQI4W/UDgkz4lZAyAPGtqaH3xc
iueCDbVUa+qI1cwrU5ZA8WqNfsFC5N1QL5MIlPW2br/8TjdI93p1IXhpJtGF5T0mdWtsa5ehFxKc
WO1lUMspGNTUIyWy2LA8U02aEd2r1cBYSrrTxc5snUyZFyBGLxLEDPEW82DOLeMlOUeLLG+y0jUK
oWy3IdKHE7IM6JwslAYNcFJumiII6QNquSfZjWlIAJEP4o5QbTwTCq7GlZjARdcwZ6+yuHBw1ns7
2aNRMShsTJQ1ICDhpxfP4I8OJAuunFxAWGpN5ReeHIBxEoUvhHKW61SMvkMBkkNsodA+AeTyeycd
xB69k5DJegNqbgRGaCA2ktT2v/m+kbUDm/3QyhTE3LaQqXO/jNf4+MQrXSGrtyMJ7hbhX0uOTjvY
vb47IcKj8rYPIIfKjv6SKL6FekAaX+rwXvk3A8fIVSvuCa88mAUcEbd0PWTRcX0nlam0SeDU3Qff
2JXK7NWJ4PMwjDU7dyyrqHsjajF8XkEhBmB8oaD8ynxkL5cZpJ0JnLtYZw6Pl3gJ0wLPS0eZdWdK
6LOmfj2VUxzC+CrcPihjxtUR/v134gelpsBipHX2Kwc1r2fQrWOcSiUGNJHf9M7AkMKEcxff4+xc
HUA1Vk4HxqhRmMJIcGethSWLCat72DepRhdzv2k4dij8Z09JFUz5S1l0Mz3q4EXAibB8Z9Tq4TPu
vHKZJX8RReT8vZOGaBYPLj/eq58efU+wzk1ImD4zWaX55HwVRMBwv4D50kC7s8gGkQXYVu7tsIEq
8R1l2zgXY8/D/cqU+5IVm/OQsQGB+Z1z4f7vDCaT9wTT9N3m8LbxZMJyvb/ttyjNpM7PcaTgeU1w
W4cOYEGqddFowlj/ogKKQuEqC7DUj5ad+tgFUtedYSJ5EIeUpFoMyPMlBr2w3Hhj4mXSs8JhJ1mz
NiZd3Yb8Jrz7Bjdlv36z4qlyE374lBBmNTGLL5zl1QHeSQLi601k5EMBGQXMyQab3cnCFBvwJPpb
o/PH9v8ivgKFMTtC9E8+tr437iQl0rM7xJHL24McLDBuq43HwYXHvoFFQ1XdrOPE+Zw4cth4V8P9
2ujqBZNf1NPWUnsXEbBFhkt7h3nVMwGaqsRGkx/S7M13UCJ3o4OOF+b1KDe5WuOBb3G5HuglHRGk
fkL+Bh1TaCG8w+DqssEOl4imnEIgpXIDyKKg9rZO2tj7xeW9UWiSawsndgK0ykXKlZkY+Y7UzU6K
zsvAtF43osuJmd+KRsDUWzx/HUI6oAhNOckF4CJvtBJVCTgGhAWLb6PLySLrC9n1yFdnGspSI8n4
TjzrGj/VGXgVmGEPybuYHM5MmOonV+YwIEanTKm6fRWbsa4VAcaIHzTcymIWOTIbfLPZkFIRvlZA
THh9peb60Pp704/NOxnUgNkfyqlQDdXHX3iMtcrbjcpq+HR9lYGAtPoN7k4wdxE2Nxen1O7bnwhD
5uHgvU6Nnyjl4KwK1GrGEeKchuEdU4z5fO2BaJUNc3kuNJDYLYSCxoNwT5dl0YNRn3zrVSCyLRT5
Xq4ac+gL06NVkCSc1VgWnCJnVvfOcHsx6qBPd9huvxgs1+ssITaGikMhMzqk70GTjhZBRrpxxd3t
27RM0NswufQCY4DXQt2VdOMsbUgtFbgXHyFuc4vywtuUy7Wuzk8tWmlQhXdXiuhU5mqeEZqWgjUy
BJww9NGQDiaYOBKa5TJ7caXyxrRJErtwnhVoAlK829ezGZmkuZbab//Irk0JV8qjK0UXlQ7bcjz4
NwAKCvzHlnXTEQZODJbz0LiEGP1Y2i7UKGpD8jDXaPFbmhqNnlVjDqBgDIzRutNExSIMwYifcI+H
jPIcP/8cO7JeR3TunIOSCgXLTlQkuuCNBAr4Q66R6e9uDwusTsIXUahFx+GC5yxDEZr8fL0Oh8zU
D3aYWEk7xPF0P5WqxYCnAmQccsH+ln9mHoi7E6+KiNL4h32bI+8rtTWlwGy1lHWEgwp+rZiaFoeW
GspcE4us9Mg4lzYJB3D8mt0ZfqLfTI4BENvOFCo1g90wdsQ8qzDFtE2Htteh4+TlpXwyXoYX/0H6
zU3wPTvZ9k3e9oi7jVyk7UmpdZRr2RSb8eUFkXV/Vd0Y5td0NHW/WDZVNhOBKazQx+g/Y5gVnXA7
vdg3Tju8p4ekyJWw2M4ns47qBsXQj7kEca4BFAPYP6sz8C4FjVH/LepDS8cFvZr3lAz6IT8zSGiX
vSBoq8P8DNVV2NOY32h3mABnO+upXb3jGDKBM1MLieWMJsEusHH7tZ9AEctrHZmTgy1/uy+AlalM
R64dljBHywSbMQ2mMP7NE97dZyY45ni6AdzXzuKhOZp8/KtR81JWqMay9kkDeroxu4KW5VSUUyw4
+6EDm0C1YnDHx61X2tuEdIvbQwfQ6JqlBpfZN3TFmcaIjDB+F3GNYbDZwjsmeGYYzFo440LRpJHa
zV2EQYh/zCk8bsh/haS7BG8cp1BkjoDEu+Su5jnRUQQVD3OOlE23lsBlAl03k0zvDTWkqQvf8r1/
shzVPSzV67wiYQE1hSrZHSnRuCWldEW34bo6g3A1taNU+x6ZX7+uVKl/9W2xIC7Rr1H9ubUfQ5Kc
9UXvy4bOpBigOSFg63my3o4Wz+ML7/2vrZCbVxC1wjLxTqrHFuWjYcjXP/26j96wYEsX+ETZuCZc
ovEUoOGNfW+OEt6lFG+2vXYAQ/VtxJlu/rEeA/XrKLHfThLW1GOP5oE2RzjXPFTCgPB3yaVVh7/+
FkWh75uYiYOGtF/iphyxBDtN3FwAykHV5ZTOBfD/OFzQ5kGxejx/+qH9ajnhOdPNhbgm3DPLlZ2C
0AFEGyPvJS7rdJDuU7tAbTOKHPzEoq7MgfOgC/3pYIpapEbtmYrNT+Q1sAODTfaYHDwRB894KsLw
B3cm1f9GbWRzsc3W/nAsiim9hYj1l9Y0mtUxKCR0ipJkIGrpfD+VOIN2Cn+Xbh2Cu9pBeouklJ6f
wJtXyu57/w1zCOsZHHA3ocwLRhY8ZI2Gj3HKfQCm+yKgd0/ybe7GbuKZABH2yMwtTBrjzMMGtQaM
5HrzChzslZujiPu6CFm5uRrn5lW8X+yRXmjSFmZN/Oqgw2uDZk9bpm6WG5odScw1YNrwDcdo5HLa
ahEKu8Tws4RXiRY3lWHB2Crf6eskYvNu6I+e/FKBL/I2uWNbr69yWBf/x//YBAO8e5IMgJacsfR0
An+C4ynMglHoK59Np2oXn2/U2tvp8fJl1hoYIjlho5Dr8EUM2XIDEtKqu7xH/TRC+GV+8WEHF6jJ
g99Dx6p/nwJw3E1x6dcpapjB1U17d0aS5mHVAhatOG2sEgSt7G089nWMsWqoEOmsxQxESt73N4D2
fLatA3P8Rt5t5usg97VhgYgs8hbbLMC+IOul0yIqf6PzjBOWP3w3E2Yb7JQvAx1R8eZMHHBi2Ucp
i+t8D1KRN9XDAjB6HVA8kB+tF6XXYr01sK6Wx5ZzVrZs7KpJK7C8iO8+Kc+rBvT+tQFUqbz8H29O
51n3anE/eBhlM3A0W5l7SknXrEeRDh2GZn1UZDcbtJmpaM6O6SP8BVUNOi9cw5qdyJQ93sDlwiIg
DJSLuEndFqwFRwY3yIAHngboK1+ei9LIjIv9lhTEkxvZCF7iG4ToKholMVE7V8aXGtSuwVKaYrjj
VLgQi07shCof0ycCGn+EnEJRTc8sO+MKHl+2dGyHmJDv5cPeCnwqJahMG+6t/gYO6H78TeSE6dkD
zPXqO8oyhD/kaI+KP89y21ef0lsNks1weRimzilbKbTr4P1gDpbKEnPu3xLjpyilPkpXQmDhJ+54
4nOBtha5IPlZeiMKgkxZ2EaBZf+Q38GQ7wM11sfTs6yZf3Cd99AOlJkBjn0h/Xcdgk73AtCSOskP
f9ZCEmRrNTL0feWLc6Cfd/PKQ00yK1H4R1xArBMZcNkE/tbCWwNUyNofx4lTnE7CGUmcikPWQxFU
VxXCeqV35Hylw5qO2U3bhvTnmIIKCR1ZjndK9Z3BTkbGPMa14Kab0H7OJa9HR7lc/SH+B1fwM48d
D0F6qQXoDwY2RqiBCXN/4mbEEDI2pDZW06g9S40GAG4ZJfKUFq0ydzR+vkBR3a0mSjhCV0O96Gmk
IVzlGyBiKR9yAcazpPbnQCGqjC7ayrpjP3Xg6TdwfmJJZE/zy0vEU2WH/a/YltC6scTHUhM7LV/F
Uwap9MnZEXTXmIp6cSp1nEYFtaXb9fIwnYFCUtED0T7ti0IuKz+FENkE0MS0zEbY4u1kiy7T07kt
iU6O+7lY7PeEsbmS9lMrP6Ehtf9lu4iEXmK56HLXPwlaCQ4q85Bews6IrjcBVwAxQqT1r13zkXFT
sPrf/joU+EnyztuqdIr0NkC4V1Fov9//43vB7LAkniucFU9GZu+SIseudu3+pt7UKpZ60MAn21gp
4mbHOS9UQX6Ofahkh9TVJCJNR65WpU44j/2RL1kIgUtzvX3u4URQm/nwcjl9sJgFcPE7D+qYXB7s
z+VBXvr4nWDogwEgdvDSLKtCRPjkKMPitCl7rGOYNqHkc0LXbez87tgwcgfYWRscAWbERZylsaXb
Zl/vwkTaZFkATViCmK9VoLwIQrjQrpEtjWq9ZaImOYrp1zjH7HHVKgtwMSJJ1NphPENsay503gia
At8uY9MLJoi7UkXsgX3vP+rrXo88NvcZDve6Up60+4Es7sznZwgQkf21C7PXN0F3vZLG4op1+z9e
+gZ9myRNEzJ/9ht26V2jCFFE3zO3lqZIgSxBBalqcqoe1o1FW4iHyqXG+bHfvtVvM8U1EDmwCxj3
TjuH8c1Dlj2RLCyBcqjYJAzzyySlWp4wKCqhOZm3LK5ji8Z4gy3VSAp3CwO+OZWrU+uEsmRdAca6
s0lM/sGFeTEW9vIpOZxeYyVYuJFI5PRt2Ky8y3j3/Mmi8L9+mDdUfhXSQjffEE3ty0tF54NSNtY0
Mb/yFfwxnRaAIHCPe2Tbw9vjQdHJrVlr6ibyKBFSTQCnbUxbxXZN35Go3tarskbt4DzxL2VCYitd
NoR2GEfo//0M6c2VOiBRZm157+NrN71oeHTkKoDLSwke0XnHmF94CzdLOKViHaJDBXL0dlV6lh7K
nUmI+tEZtl+sU8hrebsQCjJs4h/OZ4YscwHH3N1xPs4RpOWbe42whN4C7Tg0ARR8s40M39LRZXoO
XrV2gy8EchDub3VLHNjtuG8fMinWTXWehVPagskhFvn2BjQFHcZAlKqyFEXBrQ6PXCXfKCDwR2Fh
czjnxGF3FVKPEZOldeNLTKva56WcFcxNRNrDAw4ywhBD6/PrwckWyUJYojwvLA/puZa637XvAkh/
P3mgKSd4XcLV3EGTCYULE/zcdz+g066ZNXZMlPZsfiUa+6n4VUYG6HoanIkbXkyfPuthaS9l4cHM
FqdQSlNifZ+rlk4UlNlE+puZllBYO3Zim6idgA3ybekL8E3UFqryiZdWnBzA15c7yH3m2VP1GM9L
7g5OuLdkbhuPNHUVu8Qroy/Ccg7DHT9UYmXY178oSkZ71bJahDa842nm+LZuYyxkeL9+SapK6Gmd
pw3+knMQmpc6guxbZaOtWjDS2zASa7EtCnxjUp6gi9Oiu/7OoNamaO28bFkfoF8m5Cd8UxfPiWC7
dvUKxvUiHXOQup0e1Mddrd0UnltVN47GcinCU3t5J178EnA7wsqWxa2+SfIOr9unRL7tNOWgB+lM
CYburJ/97r3JOazAKT3yCfquv3LR7PufGVQNHBASpF0cDTI+6Qz2f8TKe+UPmg9nE+wDzwY/VfNv
VCB9Pqb36fCHvO17t4/Ic70VHX4Xy3eF0h/gRAFirSpxCc01wBGoUOZFTtqXT37+taxfL0xX4g+C
4UkIX3OadeHDSVPeQNZFSyXVBqnmgO4KLNNqB52b4za+mHzHc1KN6GJoUeicH/UMqYLBqqW54sAa
7pvJGu41Ywij5GNqnnufgcVbf/294QXU8++k3a0xqw9JD+5aHK9MxeDvT5+TOFKbawmpdB3KytCu
LTO2714Bzx4F/9PdsHUSRKj8jCWBwtRYskDAShV1eY0UZaedVQxPt5MNnLs1DOqh6jX91UdORwn5
TV1IyCFZuFhnQlq+zIaTHOyFq3PLRhDOpyrrMF9Ut3qiASKJdex4Y+W2qCk64Ne63/8inpgM3F/h
Nn1wMe5mFZUGDJH6/32kfxgvXwMryCOV12AChDAqqE7XSYa5bHsM3ZAvpClZHLALR3HiRYUkxC6R
z9K0jwAH8p4SzxyhQAaToCClJw8UbgSSzoKLO95O+o8VkW4dHOWgQfmxa0KRckPoU3ourenD/adk
R1klcyOx1yYZdJ4zGTAbzWIO7M1aLu4xrCsxETQ8Dop0ykxUqBN2QvyvYRuL3tgUs6/GNRoit18F
wRjaSwOWwkCBgIK9oAx62rRSVWISKmTP1YjqpwrkNXIaoNGs4nQtEnz/LNXUtxAKQ9a5J1w5vitH
VTUmwGKGdoZQ/P5SUZAlDaP7VXxc96FD9j5NV3Q1woqUo2s/GR/qM/hNHrQlJHDiTq6DvyJCPAaC
AA8L96oq9GzIiesZUfwMrZnNbFO1eTTrlI3NV4a+Wv1tc5mgDZwOdRXyfL1/POxM2feCu1l0eAPp
BtrqCMU7lZFSHci8mL2/OyKmilUeXYisCoisq3GthnjVgiI6DAaRdZWBEV0tAhHUTByAzO2MzrSg
L4yjrO8TB+dO6u4uLiGNlZWBIADdtd84ktL4XHycEs769SIpYE91u35NqkKy3qQWiCOLGG/NmcSp
lrZORmw7s8eOdTQs7c7ji4sF0FmCBureYtws4t97TGAj2tezOodEGY2k0QrJJ4q5tosP/9TCu4cc
7mW5EpLFHljEKop6hSHNT8PsbgtjJiwuWUDcKH2B19yE0Ie+ZrUgAFBBBFURu/yWxyuKVhLziBFh
4/3gR9xDdZ5W9WNGFJtF40XfX41wz1HzCL4qoiMCTjXf39WoqByYff80KYabE8RNyk2YikhPySUK
qqOowMwGuSb+vq6roAyVGrw4u2/nmQJ8LoRIEdNlOollhW6euWR/fVnIBLhFmoa8AX7c2LaOUdVp
pLvPnRKQdyPNOfN8RkTfnU8Of/EGlfSCfk6Z1TxB118tjqLTFUSc8bnKUgJ7rapgvE3GLIIP/XO2
M78GIKS0SQHvFA79JCm0eleW+ERCJV0ICDMVuZ5Fp3MHCYFJlOuMjAG6o77MmvRys69QLReZep2Z
QojYUpAMDcd1SI8yqCpeOB2fH84cMsE9OZOJZr+y2S/V/ywoca/mmRLA8b4wrz+k9fpM1aS4gL7Q
rBq8JwOhcbIb7qJD3lZPC98wQOwabDKMub4csMEY2zhoCm7u7WYa1iLqkxzscd6ReJRPXvTorKiI
7ZYZM6AHV0opzh/Fu4YtHuKwCIcgEbnPbM2/xJmGNT2VgufgfP7RdIO+1jpc7SyLmRnVFXKDoRkC
3jEOnCrUOauixqX+64X5b+Z2RmsCzAQovdiGmQBU8RRmi9TQy2XGEl3K+DdwZGa8T86PK/d6jFqq
vLgpie3mwZSjc/YPMifiPUDa8DIBY9a9eJX+ZG8r27i4T3/1N0jOtzCq+8AX/DE/YvmcyvLT63lE
wrsu/k56vQW0Pqb7KlFknIDa0RwBuyJQjoeiF6N7ybc06YSzRh2Vsn87I2r+Xlw5bvBgO/mhA+WA
nFWk9fMrnXnVzDVdnTdWB0LL1IQAjuh52G+rt1O4ba3HuuDaBpFDsRUYFPX+X93s168N/uXUn0EU
I+H6otem2GivT4OVTkCXa/b3POP7KNGFr25uaaZ25fr3zkTsDWVohYT4cZyoYm7GBo03n7fkQKIB
CB95GTal9BZjxdJ2iEowJvxCrvhZHQXfK+6nYwnzUwbuvO0Fdygj9PegENKxczASnUA+9olyoeAc
D0MYGKFec7s4r6cvnUwU2GgUBWYy+cISQwvxKnglQJq7yQGJI17U3IM79CZ9yCNVCstR6YQwR+Z7
PRiTVIVcWURput+Fgx4tPbyvSSTgQRvu4iDFU2lEBp0UtiNdVAPPk3Ppu7zoUGU/rgwUz9oGm5TM
ZrK9c8l/Rf246//GYAaY8+vwdODSbO4NDhdSY9VWMiitIXsPy7MlOEem2KKnnsgJUyg3rSo5MAF0
6EoNcFUk2c3JP8oaXIJGdR6k+1h++IOcHIp+L9n0fSeUcyLiiGxZCq9LpVVFtWi2NQQpHquJWRKb
7Ihpn/8RYMVeVG/xD7+flNYXBx8dkJtLQdLqm9a0mdnMXkgabVml9/6uJ5B8Xc8Mvz9y8WFXPWRu
uonXqmY51cnFV/++r/v/mlpr685YENN3QXBf45QrtdiYJNEbVzI+e2OHc7FbQqomYGN5Vu2BycMH
B869EMu3ykrnCe4xCh2RQ7QI1Masba4gNz7x4Gm04MM6W42A2Wa8WUclG2Yu/J+ISlkw/JL4o5QG
GtOy6PdqkDr/wD6X5Nxa4kcGywyiMUL5vLzWShILBRrYWSX3zD+pqvxT0p40NoHTFUnZeXBkegMB
j5LQZaAeVL8FXwNLMt0HTUhJsl+V0LCCsR8UJRedCWImqAeJMeTXaBzVvjaACqceDZrICN87vKEa
12raul/frCerg4FLS7jA10ealoejFJOTPRS6BWeud0K0cr4b95OSRFQ1d0LuYi79vS7FmFBokmQP
0QEZsfYzQON1iwAfOfGGpImHMFGUfdePh2syPBQlTlSMu6Zv6jakw4PxLeDD8NyuFZFV/xi5vYJH
tVQRCda85kdpOHCygumFhkJnt1myD+5IU1vTcbVsLJU4BJeWNH4iiQf57R8UiRXnmvo9mDz1mqo+
TiA33U2UT1Oi/NDNDAUZotb64fGY64q5ltoJQgpOBj461SD0XxOZvg6aTIzlezjnQO1H5hamCQAx
hdgAKa9MMmlYFknuID9CgVU0nGglhLmkw/j01JVKGsfvvwDz2RvvXyLa69siA86DUkQeY5v8agFu
pTuolSFFc6N5bG5A3k/9s9dRyLjZa8J2kx+5SgMD0PS6WMh4zU2YoAboBzkOwpMeAUljCdVZsbJ1
VKA0fJKMUgK/aiuZjp/3/ZQg7vw+9NcCb0JwwaaOBWpz42+dT9LkNi2xt5r75CdaWOM/fg5qewCf
69A9pcKdfgOzuQVoYnjnODx2+or+KYWWlqTEO4fTVobZN76hCdpBYx+u6fcQwhtJRtlad2n6K5eW
ZezIq+ttHCUnDxmFs2nTNF5Zlqo9caFXjnQM8bMHGLBWnji3Kpv6XLsgI+3PRIw40VZDCZOtXZmZ
IWqd01eaW5Fkhomz3ByhFHAScPdcHGmAowvoq5YuM/8gowE/fGZBJSEb1OoBTauqkOp13Ck1CZ8N
75LR3a++JI/K0lCgFebFNt+SAhr0K0jX7lVkVNxihVw5CbPiAcnVl/d9oOjlRj3wAyxyIlQYpgnB
3eoHvmzns47CCRcWAYHhsowYm0FvgVlE/1YtgCc2jgafYLFgpCKJ4t4qx0X4qsNL0+5RQPlYOPBJ
qzGqRUHe7UZ7D7MDdqXMxpcD9ar7rXrgCuYG2xy5pERgfHgxwKzaVWzOhZW5HNXKkgXacHmlSfFa
Vaw9/KWgUH3gKsCOX2F2zmDIV01bslHVDwTrpD/Eex0mW27hvZ8qB92S7BfDX1SSvLXGPYHZKbCH
30d3jJH08e4jcFKxeuV4yCsynu33DkbUJuIYM3UJioM+gFffH5JI7Qb0YTBtpYjumRBmPspGPm0S
mMNVfAhCoUOeV+cQHdKcLroHyqGj4P5EGN1KLD8MamMFfmKtjG7//Ve6KiPwyTZQ2jXfeQBYxwBs
llPOfNdGaUvvhDvgipHGPY+a2R1tjfTTIGbPXTtGF7q4Tg9IcpJGSoyRlDOWQjyUeNi0fCBF21xx
/dE7cl0KuUh5BxhlxUjIMkeHJROziVvTHG3YwFssU2Lk2l+MScNn5Kh2EO4Xi48g822hPz9CtZN8
TqWeB5YvQqkbajOnJX32FjG/2zs1ZP56+DR46n0puduZGmOfCSOtWb8pG+cLwbPBA9E6egoOMSSg
rdWwywY55jeeRFgbUqRhwC85fDVjK7UMH0ROpZW4RMgBSelpIlrKy8Qw6tXjitMF3urrKdbhEjGA
RUGmM/dBrgurjfuzTdey4PZrHWvCGrFbFoeVlkUgh+BhFevWXkxpQ+IbkV/FCcmt3Nlq/2TMjaON
h7u+dESjAOflfGTGowAB5J7zvW2QMZ/lLFa029uRQR0rX73Bu9uUN1acW4TynpKW/wepePuL1o3E
EvP8sN4i7xCvLLeHSp8EOXYCT9v0Mfhk7bnA9HT4GLCfAXLpI/DXdUDqUCwpZ4qV9yPLH3fw8h8z
T2iVq5+9LWqfvOxDbLIelAoy55vw+PVJTgfD8wiaywg21L2e3N08d9OEwL72W5eaUya53br80UII
56YrKzg4++ndWaLALQmv9xBTcuV4AV0WHh5qkOUJMpZ74aWm/7harC0Yf1pwA+7FQ6MAgDh1f99S
qXR+dOLdJ9LvNW0rW59nghiAEu7IT4lO6y9PBwHWe1Om38RqvhENYVDU81LPjs/lrUqE+B8FQGz0
IG35NZe9CZ2A2ZaNrxZ6UPWAG73gdBuguxWN8qIFuO3GBhSrphzjqPzpwEZuIdCrhIusZIvZvfMI
m+m298KSg1raZ5bZyTUUBr2Vl/Aa+UXbwBJiaClWORduqZbhLhhMWgH0HQ8Ar1nafVrATZZWLlw/
BsBv3CEz+Kt7WOY1KlBygxuct95pnwVyA+ElreLo5i3+s7GOIJmvogEkihTBruP4dpZfQmNNBNVy
3evpWPGuL+2ti66uIchC27OZ8fw2DT6SZeo+ckvvrXi2DmWxu5q/Pkad6ort+pJrh24WBqGxMRVt
bcBudpom3GKCeDeWYOLz4+wNGTKwI43PCORvP+LqICxwQ7fAtam7bBNTyZPnwYjPzF7wLn/TjpJc
obL94U5bnT9lxAiqMctiOCgIfAWqNg9bVxhFoOaasBhW/5j7d/0gI9xuzFXHvm5+rzU/rajQLoI+
fjM9RNXJSGeC9WuLIOKHa0QDunIWCMY8LCb9Lcw9PwPPmI+uPnqBP3oZn9C6QPh033XS/vMFlj1m
KSKjwpNwK+X3FfGUkPfSnxGNe+RiNPi09jn4S9zxzhf4KWo5h6C/VyNxr8KFQvkGC+vBdlhWcqPg
GUHteY7wK+Us36RnxHsTG5/DAb1Q7yJul1fENZiSfN8sMJME1b94HkMNeMYbG6UAgOGoL4yYM8KH
6VVMz2VmDFWE0NqEsdaXMOFzzDvXLgnZr1+heC2ZiWplORSIZsQeRQexfYPXe0XHnujzWyRu3Pdd
qQKbP/ykIgTCehlS50cjHyyICWE6PP6vvxdQw0Ta+sdIyuokcxNeRaiLo/MDozZc16/2JRfM7NnE
XifsTGiIkjc6Y+fIkWaTNtWCH3BOtkKxygfAadmF9sNQXpYoKaYi0LkhEzx81rWYp9xZnpKqRhvN
n/fCDLnTRlQhZF0aJ475R6psxN4x1Xnh8Wvnr654ue+yCAN9ML9GRJBBxKmFxf18qnWos9ZSEzei
Jh/AktWioEvh8/tvuErpDgUY+eEp0oEgRCapmvqAsxHgFjhCGoH8kSTjAWUcP10P9Syqwd70Wom9
gAffKKt/yIrTVG09bB1ldEaD1o8xOGkNJK2gucpdVd0T8YRy7OjSTRdT0uREWiz0vEefW/CUQNiG
T2y2VtCK1XX+BZCS9sM9vWCgbgyRZroFwoNTSiqaw/ndseZ31ugvulMyOdKk9Zyx896U93megebA
z8JFD0elqnlNceWsdNHzV4uoY3L9lQ6no6766jP4Vrkz4loWODwOdpRvxUKsJuBQd4nlXi6w3rjh
0isBMC41RwMj1bP/G+E7wir3vgMMdERxfC0Nn/YjwdWd77Y7cQhvrFgQAetisPjpZgvcyWxUIm9d
wx5hHOx1YTLh8k9EvilG3CbbiFmzhAyLwjlIXkdbA311galfzP0rQRDjlrSY6JWIXWz4dCqFhtMO
ohc0+A51uVCDV8Kx8jgLbdVxVl7x6CQqlzkDJ962K5CszeaCxsKnYpDxkr/7L5dBdndXbFSMHMz/
6ATIJSqoA0eMBzRHQDlluy3JjMB82LE+s5jXesAjikMCCxqby/4dxeGoVU+FaDjxsLhNUkl9enJi
RrTRVu6XPRmcYTKLqb4sV0FUO0+jpUG/lcFz0UXAWiv7hC5KuvUw//3Oq4pbOt50qHXogZyPmuGu
DFqUxthY7eJX7WBkSGyzGeY41pH0FNmtKZ/klWdBqMbU0lfp+vw6sD1HC1bHHPEMOZdfK8gaQ99p
gSQRFHnV8j0CmuGHf5r+cu2szElRoRHbdoXgLJy7YxylfUpWwfyWfFoB3kwUPdtlaX1D0PPPS//4
lBe+nuFojWtK9dTAbE8cLQUhSYpQi5GJvYJBhe0bUw9Y0PDS94DqNFgslxx+sI41iSXwDbU5+54w
ibSww+HWjjjPa/pTi/XgBCOqxZakU6Q5vmu/LsG3BXieQhluiodRrcZlAamj7Xc8DoscFpKZxp1t
WpvSbUVYsc+hrdkFOZlU5JJj2IOZfOPbOibTWmqGWL2r7S6jnzuZV3WQXz19fS7eGUAfdCTxddpJ
YEWrFUeA63qOxixf3acJoFsoOIhwipj4LSlvtkxBa67diJ7xGzZgS5DtHXa2vkIZyfjeUSk/TVjc
Pg9ttt2G/+qD0GH38hxiyV9C8j+kyCsiQ6eF8150oB1X0s+BkRT/Z8Dfer/NPXX0O5BHT218zTM0
GlVqpsGI6r7/Yy7YN+5Vc2C3lVon/OxZ4tqy22TkSNdqstltZ0jOJ63N4kJwLjM9aLUB0aYt0ZP5
y9FVt52/xrgGa9aFSqU30CFTrpM2yjGmbt7VHAtrlPQkcW39SYdAA0wo2Hg8Sh3/1SPpK+ng6+zY
BwdPjljbvcoV6mRAlDAGFD0OweyTnMkcvQCpnz8kMT95er7Ayu0Cz1Pb5aQopLirlfaZQ1c5Ck8W
YJ/h5lV3taZ+j6qO6Gz9QnUVx0m4adlcs+d74dtFZSQZ3lEgic/q13ZBz8zzWt1ofNTSEn74YpYl
1KFlvJ7UKGT36yRIkiOxDrco3SmqWhBZuNZhM4IpUKzE+c0BAe8zPEoLp9FehAA9oSijbtA7pchB
bdHVGFxKRs+Xj0igh+xmpzWJ3RK5kzlK7Gwz/jkBTvMf6yKGYxe0539VIsfDZ9kGm4YyUVjpsRK8
n38YrMpSqED18gdnTc1V3Waqx0p4rg9fBGwZT0HZLJJUzsOD3YEXfHRMHbTmtJiOvtlE6y/LwHm1
0ez0xQdw38GHVtrr+6WQz6UQt8jvzkYX0JVBbgpb1AtnCnZM5p9gtswxYJ02CwSSNP3fNhh2iXhg
YwXqD5Dz+ypIQ28Ksh5ZzOsTJixEMtlHw6IqBJFELKx1FXprb+L8PY5XnofyAoZmsEAnez86VdTB
xxye3Kxv9pZXM3AcBpuFch/UtGClEQ5rL6hEmE/JWJRoXCHMGI+Q1R29fShDMWTficFY5LvVIeKr
elk0E6eOzUiJpYvMVx3Hm//3zhItmNrnEyR9IcEd38U+nMpUngZO114rlgoFWs3hqFrggBcjluoC
FWaxLupga/I3s0Fi+giFBX7tl5TUW6FEMqoSrGC9FXAy8nZ4JkM9+hHCA11koRkPhcOXRSrOwR0Y
4E5ryDDUuyPU+BWb11Ss0HUZSRd40/T5cpf9q+t6asbNHJKoVAGBP7ZEO4oGcM0e9+V08jWY3U9A
5Xl1BZSfYly+KwLMhVaaPveu4rFxjSrQTAtFcd/P+xSRZmp4FgcyxG1pv+D5sZ98OxI2C+jlFh75
PFU7gfqJkg3P69p0npR8PPn30zoBHOAl8n/5D6pos0WMnq+RW5lRS/9UQWaaaas4CArPiNUnHpzD
ZeNt85QA8V6X/OAt8BnJSSaox9L6fegtcBf/cTMwFKUuf23pbBv3U/Cejn22QaH+jK/jP1e90EEC
SLUi1d24NiuyTp8k8nlDDm9F5sOeaPhRzTnfW3DOrL31JmGreZSf/KpE31S1YDs8l38tW622leji
2YjczHSkkz+K79qIkbzMb7YKFbbJ7BvpVX7YqHpxNRWVqMTgKpVr+MLpqWp7+UR5RZ8hc9vYnxpj
Clpdwe06gNsSyedxw0eHG8WryDeuK0gGxt7yPWnn22Cm0kXlkm2uBCJGIgXQMVGEqwuFZolaOPF0
hbQuCkADKX5r04pmfcR40kKFtakM1Q8hGxSsRW+c4J+WIusG1FkwwIPA5DfUYX+alOD2AyaTCESB
rqXXNCCnNO3OCQ2PvLWJt1GP04YpzNSXC4mPi+vvTniI7LAVbOdwaP1TimBZdhAZvqOQHHCkt8XP
XTLg0OwAJhr+H2WKd1gLM9hTcZyLlr5sDSV0imbRIcupj7gFaunLfQYCK9IUFtOGtfaVCK3nvvmN
PtvTiAyzH4qpFyQVhsMidkXt1/ciL6RXuKwOSQHsdVgS3l2hXhF1cc/sPCoTSh+jE4GnS2jlRN4G
T2jmvbwiPKucn1z+aNjuws9CXQ/QoNzm8CYcFZF2TqMVq0jXmAdDSZTb+2N0t6y8JKNRVNMtCUIu
8dOnXhvZJLxKbJuh1jHHyo3qK2TYP430iIl7qyyLyeWVTwXpvHUKavES7RZuD5clGblRKcy3Twjk
qRvsdABbHJtktdMnMGEpoKghvbvEcFap0Y6O3l9ZhEWjr/s7K5IWpI/BOAmMQS1tuS+jErJ5brqP
9aAswUYIL3uD6rQkx6LkUaKyo2TLCBy2TIi1tEy1+qC5k2pVGYtRdsobkRvVXiJ/dnBfjihwGGqO
t2nG9H1EopoqzVYIV+afL1nfp49FXXgQHXKtOjBpWkXRsquddKsI80WEf6pggtpDRc40bzzD6f6n
XHJoTZi057hFpQLygthM+0oV8CwvGctlRpmyNuEKUTf5fAYCBfOgKHKvTaBXDCg9d2HgSFd155Zx
Hv4bF/3dNXfZctr/SMkRI/hVePa+rdsV1cjku/GDZSxFcUookMLvhABdq2YB9alauzZibTS5//pF
cumt/hpubfpKmPp0OBLctmTfxlAf5kINmI7IxSQxUeMj854C2m0bQz39mQjxxd0MbQSAX0Eo70I1
3NMcO0aboe/H9F7yUbMAIa6YgvaPQA+id3jS3dKbedVm9daqiZ7L+7mBEGc18+J16yPlZv7JrnTw
D95imjwslWXnwlTn/yPM8b7oVNFHrEk23CfwU21cGvinKe0V5sm/vZVg9WUuY/SkYZRxju+eHikC
QyymQP7nH33N2Az9sCGHl+m1qslbkXRCS74iVFpWe9VbPB7kVbasmWPpqXWawCAh9lnqHbzy57mz
YvZSESdF7uGvmCeel1/dF+vjMnvX2mUxDVov/X3FtnEk0uFfuuNL8I6tEaUtRstZEu1ZIDjqgNqv
H9Yf8guudaNvt0050myY7lI478I75qnGrtKOUxpLbyIKGow99Aig0MWD0ssO+CkOWet+Xc6/58nZ
kO8kbqTuzA4jU6R2C3BozowiVyaGCNtw/ve8n9Ayg9Xxm6+k2alaMGvNh0faG6+Ix5VmOs/0s4HT
SM9el01S6feGl4SJdzFL8bvbNyxLTXHqSMJBrPop00EGYHuNPWEFDz695quyFjj36PtgF9Ogjb/y
lt72pmcSiB2rttWXDjJguBOgxfWlIvX1zQRKu99FIrB67EJqAPDlAIOQ6nSp4ZbmwSEBDJHLU0tN
PkrQQUFEu7o+wIdMPo3/cXQQIyiIjKHeMgPCRQiQk6+PToCGIjwSMGj3Ay/8xRpIQgslu6u4czQ7
XdODKxLIVRvalkmqzGHm52isoQS1iaI0gDN/YIEbYcpnmJXGsjruSTCpqCkK+e/oRVZDT8Zr2Vg4
IqVd1hSlygUhSpITPD6+29IDkxUcAHK0FLR+zC6GsHyjVVaNdJMrzgWXpLvvqZFg0YONVxHxd0qT
1BUz0omEzeYnEFN8ZLkri7KBLf5WmZtaIopUfV3cZXHiVvyP4uPogS1hPkoKZ3yHj7gJ6DOmsStB
NEo6CE+yMwh5BJwPvAfWFgDFALbm2rn8C2n97BiFnIW657UwlLgFfjRVRGwrQaA/gQw9LWRd157B
4levHTSDUKhkXbudBwSaus1CDp/9hd8FtBrTw9lmIFyWKy5qX5rMQ3WiVdB8YhYGUT23HoKoJOIF
9IrtZma5W2C0dJK6+lxHwkzd+HF+6s/LZKl9icRAqzEfKcXAOmXpZ3c/3yX15HT0f2Oq5RB4zsmp
bkj4VHFn8qj+z3deNrak47iwO0wCqI0yhxZZMxSNjMZ4CvA/x4ZD4ztN7Wj38iVfHUaGx8iNLhW1
Iyhaa4foGmDib2DyPKUw9CHtLSFmJRTwINXgZA9SqMmqhJ7xQaCuvVKvrPxiDf9qM59r2J6NxEcU
Bd2p16VB+Zu3CfVPqmvKl47UnSwNFmJQjhvJOlLZaslBwi7vCgAO15gI5QFuajills4cuKYowXTq
MVC9Xqd8Od9d3nFjA4kuGSbWpss+a3hG3vSJNYOnr816rRSvJLs8nctgutyeVW9F//ZFY+LEEcRk
garWfKvXvZ4LyoA0uYKWfBGApmPINyo+PM+I0UIiBPyM8wXl9Y4LviGpJ3lPLlPn7pRJ6vNkc4R3
fHfnLXYR46KkwjXqIBRwaBVDeGCG9IvxqWGXAfPzyptRYRcIWzIgi9qVJKHsXEDIeNij4QvexnWs
c9zxHa1uSiCJYl6BdfTI+i8YuqjcPl7x/gLB9sVdZdIvfGUjd+n6uxj8aN7lpvAZJfky3gndt9jV
0WUz2bXh+f6jIXsf2zMfHmDrvl4xzDMqG21xSA62E5Nb43YuXD67xI2JM3AiwGjrghjOhE3G836h
VunJinjUFfIy4+bcUpMVcvi4T+1N5QFhDuGbusUrCj7RNhdvG1gVIbl1f8SQhR4cz6CQtbhBt3z2
INwB1heJ7XhA5XM9iGovuZMAf7/uW8AwZf44FXiQ75aIQr0c4iYl+kY0L3E0KWG/IRXS/MLQE2/H
RbtLORiv/L/nwuuozznoyN0oOzR1c/BabDJMPu8jlYC0ZUe6RAUd8NjghVRQVvZpwJF+Gf2h1bCE
1mjInH7T/EGNGLcfVI+gXDAANlpFM4+fyC4EiVU1w6vygvUnP8ooQydwZqJOdRLl7UIZuxd5vteC
0qU67nRr5Elm+mGxPVef0eI9EHKghHtOGGzo9VsfEneUjL3EQzpTXFZeNquS68c3oJLXoXd5RyMA
G2bXZdzcNZpVVS53NBuFReyZLtJ2j2PWotuJRtRBwcVHMmK1zzt+PsjEmQlIDW5GwfJCIjSOhnZP
YHWcLZr3EmJ8uHF3l35pWqXDrOsfU/8iqLWefeYfwPkBJiX7j/by+oNm7WcpwR4Y3uubSmG5zSHg
/noRWIH8NVaXY8zVPffGCWYGrU0gyW921ZGMl/al5Y14YguLP33L0AFI/F31MwU3RnmwsbHC7VlM
6E8xoh0eIF6gThb+5OAeXbo6M+VuYuaV0PGJHtMjNtRxnQ0TDtBo63cMzf25PeGjiD14uycST1TX
2n+H47hwJYXLUmBdzkKxZpv4cGw5nU5hMJe2LW5uw6NX+Gim/QQzMMHddwfVjOTA+EzIM7Oeoth2
lvDTnOd53BeqDiyOyoD0XjnvMQOqwpcmolT2QHMvgIuaYCeMhE9KnNDmUGZS6heBI1eYIsSaEnwL
afT21gQ2yVZwhHCwrgQJP9v61Ho6vV/p/wI1BSYbD8hbtm0Y8WCgXRRoOxENWXVFkrM+ht9m8NfP
VswL4qMyXtsb75uA9VlOGl/5LmPv7189kH5x13f+MviUDlNCaqFNi2yS5Tue6ar9lr4XNimhLki2
5v2HQXYtlBh19eF9T5QdLnqXpJJEoIbCAY3qznruEIBwi1XKhYXnihSebvk8RrGt2pp7gxrI1FJg
aq2Mu/w0hKlwVX49b4ynY6mUcslYpRDI/1PqoVa4gFcHJjY5QFZ26w4Y5XoUn0dDmY3HmD1bZoey
BaFbqB45dBcm339V4H6YTG6YZAV/xhqwHqy6r7YUkuXROQmyAnnkUsyhWz+mUl9bt01f6wKwOrEN
F+HNkl007WPaKbAxjrOkAsp7EebxjTqA48NaSiPGEqLfKz4vDjSdIL4d5E85OQXlBJ4qxpZw6jZh
2csXMHOjEn52K9IoPUtYm584xxPNPUE3qZDpG9RxqkCLqpPzeuss8FNAmro2osLQ2ViQPmX0D8fY
HkrG1ORKhK/f2dDuSBgmo5Vf92zzkdVgmxZ5YIWRNg6AeLC12kTupqvtBnlsHf1Z3r4OxwE17r5a
Ceej+TPHhK3DmFXXJ0Xbf1aO9bIufinKzUaEGSAnFWUwHiq1lfkc6slgpPjllg+0uvx46aCn1Xp0
adf79Tl5So8E9XeHg/D73l26Z5bTIdet6QmC7o++WIzfXIhFLpFfupU7aBQplKMLs81BEKzGOVyT
AN/aslU6thyksE8mmjLAuNxD+zfcyyz8GB02+1g7dh5X/QOOahfzPN+x/wDCsi3vH32hLIYRsO6I
cmdkcu3OWDjAmZqtRk86SCXW4p6pur6qD+Bsuz3fIWDtI3F0LqAYs/oMomkAWeOc00WCzlfOsxfw
KNgTQCi08F00RIY6yuKDtdf8lJIJVOQPNL8jhulft7vxZdQMm0sZot3HBpkQJN/k81Fzq+/kBdcS
9SBm/GVtrNmP9rnnsPUZ/sJjCnmMfV4yOY2R4V79cMddgG6dnJoft2qplbsWXpef3NSeg+MrPORh
/GIyQz3p9RZJtHo1wqoevsNdJZLj3mPO68fVfYR3pKIKnRe6NwQsEvpgC4OULYw7ae1+vOyJI7NY
7/dvV+DwnONiEIGJtbEiSl28JDHnhRBezRXLHTYJ3wvjHvzR/fj+N7XGDyswZNitmL8STN4Rx3FV
tWybeFMvyYEuzhFOZo0mvgNjfYGz0drYf3cVhW8gEF5NHwojHVlZ/UXQuDME9upGiRMhCh+Du+U0
oK6rhgZmLBTDmCxUD7MCAXkdRr6eu1PLpMZABFVKSDax0j04VPE2o7hcOfcsaEj2Qnq/isOGvySr
IhrBFTSd/0rUSGJ+wJgusGcNZZdn+1gSk9/lG91qpu+GleuHJsOb1rjsDgyArvxfM5ZVr1Sc3f+J
9a6dwv0MDQlV4ToPtl0Fc3gW72ona6RLN77c6mH6j2+7fuGfc97aub45JIKqFj7HYXI5vyusxNr7
kpafPzaveBxGS7PFyNwx/eAvppXafcBQElPWMyB1MDf5uGgcc5ILXbcJ/kyEb4WdY/RV1atRHsLg
M0vqHnREFmrWihGhchHdia56bwp7DZ5KUXX9G8LdBDx18vR4eyHmTlGRDPO9Vnr38wSz59v59dQv
oqJTfUqURXUx96K2CcdnGO/IY1kUl/h81YZ3JqfaGwiRFjihoCyuXNaDKmaGHxY2OiNuPtADsF0S
AhEThNcEIgqKpQGRff/VE9PGleEuP70zwN4sAVhdj8bMx5MpBlZdZsytZROW5bfEpQ56yXKc62hY
WbxRL+IvW5TRseMmhyJZ+uRFj24HgqMkdiWf82lIcMZcsZoFfzqxCsJx4ye2CA4uNOkDbukRSMiK
yj9cvAR2lnCsQior2bhIOb0Ep+N1+B6MPzMBXkHhSpkS1JI10VKKp3Jd/PTqv2ki1kx6IHzHQEup
7lVDWimKitoInePcBAc96NXHUmmad4afCgzn5uOJ82xeM2P2OnjbMIsMRX/AxX9Csxk0HgaaCnn5
ApMRyOmQoASah9aqvCLfI0kAJbB5DO2dsZqTp9QM9WQF/tCSWLHyrDCKfxrqAWyLakjDbXFPWWHo
Dj59Omekjz7NhKzOR1pHYsYM+ybaw8c4jymNYGPGsqRw740goktMd6td9MCbnAWSbWYD2N1WGblO
URdmRCVov4CUqHA1rgqHGXbDEmCQRVRBtsuFWVByw6pm0ZF+A9rbjkTEYnlMEkrjWyXduVClMddD
Sw+t5EvXWj4pHy2fb1FnvVEj3E+5N5RGbEIe/DOdA/F0Z8r/ITqcBRX1YhG0YCIVKz3JgxdrNUdK
ZgUeH9GpkZymkDTLfntf1BoFPCLI131GYbzZ9doVKoTTCqE2U1VM6gNa/abw7+F1SpTwoa0HOD4X
lk4Cq9JQiLZ51NlRjk/K4nEi+tOFppV6D2hbN3TCEu/Kmo4iiBSPjlSSzvoA7X7YUsR+3JnUgAPQ
faXYPJFnEvsjvMQ6xuctXHouYba5tDDz0b7YjBhy5xR2KUZE8SlXqz35A03YhO2w4qLyah834CsD
p24fgWk0StbS95ifZ9tOD9iwZFrxJM1aUt115eUiEqMNQxkmD9JxV1u3flpmIT/YAVDmysgn8oSE
cXEaRuWNhagYGj4+zDrpulYWnOP5Pm0NEIY4URT1z+RM71GIQ7H3qFFQZSy2wCP7Enkk8F7Zi3da
EJ2Ly/0LZThKo/wO1OUWMWLHKQYbHLS7t34sOtSmagSfdvfkua91aTaGzgS3wZRy24mXEpGS70hN
AZ6mioFmz5mEHVM88fLm3bjxTfCGimBaEne+cc+vt8rHXt30AnAEaHGbew4dx4pALTttesaFLUdS
RaNB6jTdIbGSPYIUt6ThnHSF2QcTppN79IDQkePHtl0tuoX3CoAjd4LCYrgDVSF+BT6tXAohTe2s
6xTo0JZpeurNPmUV/tuc9o3eTqeVM9fdpypIQSh9+YFBYCT4kKkuqc1UEGntEx5aaVC+CszuZVlm
6kTbPxD110jfMnQ2KFzAouYWmPdHnjJpnKfa3sCtMkRXh2LNId+AOR+NxpiP54cHS6NiLcT8UpyV
VS59dpojaRLHxuJhIEwrg9sDYsT5n539Zmz23EbIgVyPtbDhxETuMYL/2MN52eOTR1TC1jyiib4m
gJfeFGHWS8UJ/JyG8LpqlPl91hPUVV3hKgTz1az3YtUQX3EqTBsHpKA2N9PWGHXlmDNuoJyI3dLd
aWtwj3bHtYLb039nkofibORsezkVkNY5EoYI5UKDAbDoqkYlgAZKdCHMgm8qqrPQxKRAz46sKEdH
7o/QfegMjoARljpdBbRNTYXtQpA0O9oBymdlQMVNt2pZ0UP8LdPLeKs9s+8NasOW5STOb3C12fci
AIUOm9cdubuwZYnHYDhtotZDmmIKN0dp5ofhrYjtnCnsk6yoPvorGG8lDZi/AhcvI8VogsPUKNjC
dYNYbmOcpU2Geo8ekhAEkFtrKdXzdKM3zD1dUaRbWLPbOWVYkndU9LT+zgw01STaNxjiEdp7HbSK
94bmp6Zq+/kbg2xz0CDN4vv9VHmRM/1+ksPMgXY4q+j6lq423hBBVnOhgaMPfZUdhuddLuDYLpLo
4OcdBs52xVKe4W/O2MWS6ECCrfsyV0X8Q2P0EXTjREoil8JHE5O0JCxeAa4dN9ZoPQ80kK5O06xS
xH64JpC+BgmCcPoYX9t7Ba0m6EfK644l9n1C7OQ68Sx3zQvnUDioaPGRQy2kTY2GStG0CuSYwHxa
Az0H97OeGNlumGvas7xLm/ZYFrY3xv/XFin4zl85YrK4PUj0Yy4LMj/pE1x3WlWy9QrVvkLP/ufW
Nrm5pN56hNhzeYTzR9Cz+9edhcIN0Ta3/k8Y6tNXhZti29BX8ULD2lFNIvvsJ3GwNEcFkRMCK9c/
J9YV6ftEpjwvENvNAyzt9a7aHhAEYv7eK2OklKFe56GMe2DI3LFPNxEL9J+cwsiJB8C+8mI0fnQl
FK+2bxoBsor99n8Kj9CviYALX3+lDgTEKCffMdBTNWdLeYcVPFQGSrf4eraVIksMdrg4drq58qiA
eBG/UKj+QjFPzDieMH12SgjoGMPEGDHvAS3d+GI0p9cjHytwT3Ei7U4nVmI8TI3/t3Eq7UOGfgYR
m5pqUdL5mDFf+1/Vinpp4fcGsmaTURFwt2QLhbwNwnTocv6gQdiMh7gvNzuEOJ89tyQ6V9EY6/60
c86UA49TLIOY0aVQ5uW/Ga4T0aov97z96lAWyG5PBCG3DCkqQOb/eiSab9DWixgwtja2/iEFh8Zn
O4JOCMDNsEupbwnSNzAe+mifJ5pQZYVWLdsbU/bV+GKPHqJPR2R7x3D+kUknRPvlsGid1d7+OgRh
LJ0ZVDhyS2D2I9wXNMuoWD0PmeqjRlRm8WChtfSXCWywPxfwJ17qkRyBTfNmim35E6VNRo9/60U7
WPsWzHbnUO2HSgI/2JCwbYU1ayibInnh2HXrzsaydX3/qQf+LSLlM4qup62onNvzB/PIQwxsomjd
7wQ0spVZ/63r7wp4OXHaTpf/oHV6zRYPpjsgRT4CM21Oh3pJzfObCjOp2rTJqstHUU6aPomHSuhF
cFjxDwN/S6IUJdOFNP+aU8V/AxW4YwtBQoXltunrb1waOhXhP0J3glJ1cDaDnoEnFDH5fvekQdnr
sMWiVLkNN+ARkybeLHfM4tJbmPOOAK4//bDxhGEjKjXYLcZ9rQQkomVCcl5lMOq5wlbvLF2MxbK0
CtfOhkdboPERf8Q3JjD1dHwVgFiT/B8qVMKscqkNgl9Hj2hEwHtpz+hasLaKdo8EtBJsRpb/csl8
EVs6NnZE4ciMA/tCsx6OjclzTdyrd7qR7Ig4oGoiHrC5JkDS3YItJ5UIQrErUBVP+kUlHqMizvRe
oJaG+zLxaCsdE66KWUAQOL8IGmP14jsz5b+avGJ54/JmqpBb1fJ7z0swHcLpH9qofpz/T0sLM40G
zMAwhTmj2N4YZQbPknIsUqVgbkCs2jq63R77LOJUH5QceeB0PrJp5I5Ituxgz738m+KHIzzJLiXe
pExM0movrRuJ7jQgzY36stwRJyEBh97Lr5+Di9WQaJr8hGw452IDVT9IwXWsBvEGlCWArfFnyjDM
RqWeo+6qHnv/OPCnbEtRGpNaMjpXh+MhM/hojdHIBEi06Qa3/9z4jp8DJLsHYXuCe0fN+rUARwOp
GhMMadeuVccgv7qXCh0x+C1NrdPbpg3d3oyIRrHbB8OwtOFtVvqE1ZcHHaTC2sos32oa2fNd4X7Q
zi9S35E82NYsCNoMG0WarwsukW4w2IetXytWictuRas/v90tNan2jLksNZzrkLMO6lmflauUB/Ny
uZd4km31efcad/jhj/VxE1PomiI62np/cZYONu0Q9KbwfWNSdohfnUzsHbYr2rSF+MPjhcq0AHPF
M5CK0vm+rc0LAYZpM4LCWb0HLzgH00tNGEtzXjs6I3LAPD6DGE4P2FUbbu12z5E6IW3j6w1kw2ND
sEfUx8jRP6MkArtJXfEqQl4Mb6NRVzyvagyid2ucoBuIdlX0ISCSoy81L0Xv5LJTzOwW1EU2eyzr
65J9ySMfEX10jkr7uNQoudE8YYxa3ifu/TbCy9Tw9OjDHoQjwomwk1EBGWVHDFeBPIQtieOjb8j0
PDsQIfM7U3EXGcH3L+hEI4BQum3pr6wt81A+yxfwKi/BxzBc451lbLQB9YaqxdSG5bTsQfsOTIQm
WmWQFCSdcbZ2TSvL8+lsodXOcUMFlB1eYJAEOA8Wjwg3t96ECP9NMLAPW1/F2jwuMzoPuSzb03Q/
Ellz0XQ3oCoHKGiNsxtUBD6R82diYxGPnI4KUeyMcsknErrWruqhjwyJLQ9pTe4F1kv5cDJNLcC4
JXD78NB0gNWcQx7/Ii26Q540XXDqFQDg41HCnRDyyuHFf2slVCIcY9eAnm8MDW1+HhUqX+5PyVUU
CFbGQwWlIz50hAL0Ca/YVoSsBua55dYTbrkTFUVU7QoLc3JK8/KQTuQP4V0MC+9IAiDmuTJHcqBL
mk8vL1KEUfD014sksSljn6xiUVD26oeUjx8jbdtsB0BCNajgEyp7Jt3fK6OrhjNb5llyZb4ynSNK
E2YXzGcPu9P0Yarlns+oHNL3xBRRt9+3CEOZezOzmt4bHQmF01QG5FJyM/sgXOrXWKuYMVL2d7s5
EWFzZueNPknLjoxXxZmjVoogkwj7EKuPl24Olvs7Fla3EbCfGabyF7nLcfSvqAL4Fh3Puf3FCl+q
MNrU8OCTcSkwziWTvYwAVxYxXJFWUkFt6RTeWjisdWnX0EFxqMxvhbfuzAVfcRLy7ohYgfSEOeeA
+M8tE0WlRhUjC61SDctxu54ZmMamhX4nXg0wev0gihr07+O68Mys3RrkbwIv5RPTIlzwfRcPYfMX
KS8C31GhO2nLbzqD7dpQVW7AOzFAZtk2sbfD1PJ3g1tZ7zqNR71cJvdfdhkNrtOwa9AlcDYgBNDA
TUU/bX1EUS7q4cGlMmt2O0B3fDwRKWhXvd8JoyeCqn/v/F68ZJhelSG0FznlxH1lDkQhRwHcCnUJ
ZMVpHFasU1ZJcMqzqFKZpczg2AhdKqr5+EVN4j3oE76+R0NVbAOW3dGtSeF4w6HgV5xkDTwt09oP
uikjNxTMgSTTPrxTzUbYkBYml0HdIcELZ0nLx4YRncZKsgCX96cuBS044tg3zagLpwcMdQTtKdhq
pZ92muxYIS5W93YA+54y2fIOkrfaeIKVKb7jJ4wFrwGDcrJszbmvwwh6sxUoWzxFI5gaD/IIRXQa
2woB7TGefPkkcQ4EA/WoWH7VAGhAe/0febqTu6PIiUQKb8qxTM5DvfSoICyr87M5sROyyCm5Kw69
7BCgWi38molHL+8/PRS0V1VkvY56vO1eU2TOMiczxlVqnIfcRhqiOOZO/7VjLBzp2+PUWpvoaWQt
hsRNWpYTborotm8AqQvx7SLy/HFqzSyCAPYBIXAgPM3Hax42fpJmogKyAW+4z8b68QfX/peSTPZ4
8LyQJKxrzkLbMhOLkVzx5SnRE6TwzXLuvTzTFCCT4NdptoMvMoRmi6jRTd4Obpx/WVQ4YOCIlmPg
jy8s5UpbromQe1QGygVzNicwKwdNxhurjJzK00zcFcaNe/1ohTwKE0aiWpEAKiZmg5kQtsBb+Ezv
C3/q5KH6KaO3c4aDpAuKY+Gu7sf/eYzoMRJ0xnXYU39tDJiYHZ539DOgvxsKDRbnBMxtJzINgifZ
siyrm66ewdqaS2uuTD3nf/mXAv7eCotoHSq3HH+VpFP88n00LVaVwEeL0vjI7BGORvzjdDF2z9W0
y5i16N81Rti52x72FDwp/8Z2GWzikUa5LbBwvFRwAmS0DVOGRP9devxW0zM66K8yHX402mCw/fq/
aHYxDnJWUp5X1wC6zgA65j4cNfgLnPqKgkGbAovaAjULwDq0MsbntM13R7gDicNpT30m+tkwviuP
DjssHTWedbMukf17RhANEAC2JSHI707rQOHcZUjhH3P/ebXx4/2IYTN0FdgZXCEZNLaKgY356M/f
grDTtT47N79WzbZx4IiwJdU/pjXw7toFLuweSN8UyJOoXR0rfSaagQqnl2NyXK6+T5pEjAz3370c
xysiJhn5rHU8subW0tUoAZbSZJ9G9C710doX2htlMnBKYPRHEMkWXR2jSx6GQZ85tmwEHrDGyI5D
kfcuXhw4vzN9gyEsvYOG00/mD40Qdt6hLj6EWhmwjA6gkIIIgg38atfYxS9E5iU/sevZHzIeYD4n
v1i/34ZfPTNcFod77UY2+RmXJPGvNeZTSqiYcyg9Tsg3BtTEQ82+lLlvZqMckNiRBr563bGRKayk
V/b52ZhyxiuqlU0QJ7alLWDRiXlDpIbBWIreV0ugxEmeCHChwu8HY5v17Fj77naNvcEnaylzhbE5
BeLRDg9H+rX0aKa07+e6VXInoI5XW5tqWTCcUj62CVtoHeBtI9SSIVtzpm/QBstfYGclvVWmNKRM
FMJtNlJEqPL+jjnuJHSdfJYL9KP6Bf/E7HCMOrcIA60jv28NsY1GLzZz0wx9e1Hiq/3MBYp0CN+y
8yKvm3BeQqz5WCmHl+/uuiEt5tcfZVDTOy4H/Tm7MZYVz91zWaTBYHSVT0SA4GK0KYQPVtJ2oX8p
Fo5zcxYgaWb3WS/1kihVIU72rPnU8gFhMXS9Ki4gyQ+eFDBDIS8ok/pY84tAab2zNCgTjWhccGHt
WoCXLCQI+fh8WK0d9AZ27QZMkOk1OMIpQMdvDPv2yRFyKnjuDiJdkG8FnaCL++5MJuX/zQLbeZVD
mJygO6teivT/7JEs1Nb4oWNK41OGP1xD8kYNnoZcbfGehmZpSmkyYHGLXCaf9GRDfVRk7jBBnnex
hTKaYBEXpUiwJvasJ9szeTCAseFRBu3N5oe9NO1sr0G00Cy+7lrqwJ/axCgp365bEApRQx72uVKC
2X2h/4tW+Ir2EFhN3m13yl+8066VCgwJ3nooPVm7+yfYfI3lYWoq+heL4OHTKrJIfdMJdWUZ/Wju
vafrtTtvT8o+tskjbe3vU+2Q6hsTem065EVktc7X7MQvBcH4KL6AI8vUxG5zgMJSvuImhu247+ID
/zWmMmu5gst68SuoTxWY2RbEXcFLCKGOnXpr9SnnvnB51dtzw6u0MdPgIrAoxNePq6CNZZxQcQAX
LE+05RlVOfPBlrD0EsvQfks3Z83szxWNywxtwQCCvMQpbi3liI3qmiMJirZNfbr4U2Y56kPBbZDD
EYWGSm1/3zwj+z6lJZXYa1tDxka/YoZcffUD6lGnd59yJyjLL34VpwlI8j6YXbKeMHkhtp4tH2T8
gfvJhThEeIWYeGTBEeWYlv0LSqT68qFsU0N6vP4dzbI9pz9NeicFQNmipMpz8fvpJP6WRA+FfQxu
idiaBOLAw/CYLDj/llWc6kjK1BvT1AjuljJoCJmeemERj40qDQ2TTNAtDuZkzRiH82mqMcPvJ4Fs
e8W5CBuRwj/zgnRw44t4cyp/al5R52EFnyeFGz3qJVVeeI+COOjkgKVus8eGj6ot388eWPz0CiFX
Tjc5HjrklfG8wQ2l+PPfNOBkpV9yLVUj3CwyDjQExVxDDqV546svsaOCZ+2Vky2iDKAd/jQJi6P5
YLM3S8RUdGfCEHcnmlV3uu7q2vKM1x8MRWWGs3iWWLWBDEsRtT4irAdg2x2Hbo6hsaixQ3Va1jfP
eg0T+P5FIGA5j/MSBvaAEC0v1Rqae9jK8ZBaeDWQIPS5hTmWkSUo5WznV/cBO7yfIBCukSBzbdzR
0ODxGXsMAyvgDGU0AfqM038/Fgunbb4B1kYP+QH+F0MGTKOYPei4jwPcuvvByzrjymM4rhZFyAXJ
ycQuOKLv8L5kGmaIqwq2k6OgvVPWx56uO4Vegi0KEkFcMFf6mcELSUeUln1NsjRNS1BedMA+DRi1
wB6BfZRfp9zpzBQaGs22PvnsKPoE9S27jJ4Ec/+LRt8Asa/pVUGOMLi0SbH+DwFO2oXxwan1ZmMN
eS2HXTS8vRXT8Fg4Qv1+wznD2eMKMw/yyVuzQRCxMZ2bNBJYXviFqIwappRPF1MeDMcSUI2Zuuo9
rAw+LCAQNpBaqtmLLTIKtY6DezXZzJwp8hDYgBB6UfEmUCZmXRn/8aKy0e/knentf5hGpV5LbL54
lKv2U+y44QhILG8W8H2lv6amd599H1iYbd30O14eIxB0lNYJcRWSu0IdQfq4iCYaJcGRt79DGf58
V2A/IQnSNCQ7fEgg0sgyuDtbrbTdzX8SqazL9qCW0qcBUxLokPsHyLcosGBy+Ba9xraDNVoK541x
6CTIocnUK324ev9PbHc0ttWdoi1aKZAyxmgZ6MN+Y9L2i/L1agAd+6azv3cYbnw6n2ZFqZF/xmQb
7D+ZPZskgLfn+d9Bn6T21EDwya2SU3qm91ZqH4kATiieuHjIgPQFfhJKf3BoAiJWtDB5KdJIDv00
UBjAAtok1F/JylExfyDeeHPnuv5NfzbThMUeP0IadWKJlsUsrKEXGAP4KGMiNgW0+jrYbnQPyE3R
X58/5FqTw/B469SN0TzZWqZQ8JJeZB9VpsKBa14yl2ZYocA5/lDb2c0I70qhJXqIiPMUd4NSp61A
homxSxt7EffZFL7BwTKQTou2ejhrS0ZM9xKbOA7sxhjqR4JtyZAobf5d5nda67oi1bEinKfF8qcY
FrJtK4BjNDI3H4tOfrPRXI6hu/RwR1PZTHpavFbY53A4yKnOsE0LwFCcKhlRwWs6TqrmFgRSF6Wn
BP5hD8DNMXVIF6LX0LiIrqSP/WNceOJwGbr7c2VocPAkUp8zaT7yArnJ5I6scyuPw0FieVz5zX2j
OAQztfSxYeirVNmE8OzdZtl/RHRSUdPI0m7+ug+XYKFbJR1bKplvc6HxvOO0VIqytze76jLFvUbz
2PZHq6SAB9N5KWx+mEx+lGpNPJIdAB29Z4odh9Rptv+TxbI81X4JIROqFidhPblpImWVMvA878y0
WhbVP3oodBff6soHtFu1ZZbQYZSQ5KF/CkPcIXCEDE3QBO0nav8U64eo8rCza9tmU18mvdf9D6tv
3A3FPG2hKdOe7mDBKeSOar/jjJkjzKhty4KCCSQtS1WJIopnmjkTX941+aGYE6xTnonxuU9bRIeB
08Vjf8n+oomJdXBiZI/xc5eGpO2C8yyA204HF1rI5kx8pySfr5+CTctRAaR0xuohcPsb0Z3miINQ
LgPsJUd/PxwMHkZModFTV1hpHr+wnoz586GPFV65RYv4Gv1sffzCX1QGmtiiHzfjiRexbxth/twd
zkGIyv5Uo5vm3M+541zLuYIZs0HMrwnq2XKqdXVvpR24Zjf6qVNmWr7RfNkET0I/yNh3kgzucT9A
t36dNUjMiH+2WUI0kK7iRPawkXk9AjdgJNRhdIYrxjeecId+TSIEB060a4em64wePCxYb2F06GK+
pY9sFIG4TQKA7Uq14QkR1ykpOOwgG3A8JHp4w/pZ45Zdw9vrONsLsC0IBn9MBb0KvNOzl0jy+/LN
8pL1Xey9+OaMalviMvdkuZ/tvGKNp72PyQ18VTfhC7f/9YnInp5y81lCql7U1l2vib+5M2PGD/cm
qFMljssRUUsf63dt/9/nGgQxrDzfpmQo9JzZhf6JbMiZEHaSlfq3yMyiP4PjHbvH+h7Ds3f7uQg7
zRLY7l1jVeDyM70qyEWmaJA9kIL8hZR33eIS94Cj1s5MrLUfcuvWGBj7fFHp6KtAEy3V7o0PTzJU
rh/0UFBTOBxhvwfJ3A4bGKRkY4fLFM7lbaCXMl+p76sDK2mkcoxN+L58Xi64NBDnrDl03lJAfkKR
N5hNHsXr9scvb0HYFdmlfXL5mWqCKLg+tcUB8bog1EosRSkaySjpqBG2/2XfUJ/E6/E86Zcmv1s5
Zbg2+N/RLZWuyGjNjeOsk7jQMpKQFsKEzrDUEmibEBULkRPLRHbQuqboLXoupd9JQD/q+OKexk6J
ffxEu6KGKkKiTPQo9gwqs+zXsptDYRPCHe6NSjK2nCPxYVkocPNLdYCYpU1vZ8LHQlfEYRqRPZG0
0zcGVD2Pasbp4Vs7cNWi+KMgZd8euSkYnyTl+h9tkpocgyReXMo8fy938TtSli3YyZ1IveExdGQH
LvoAMYojAFbch2QKlJF+acPpdcB1g3wSBid9qG4IES4ZqU2lQlqH4IzPVHFqmeR7atIExakXabY9
en5LvbtEF3/L5LvKGezYVktuJyt9Rg/A8bgWfDjdYUuRsF1IQo4JtZoBd/4RyJNCs/wYnd6TX43G
WgPtYVYBECo0Z0CucZz5aNWgm8inhyljeothE3OkpSZCo4gtd8MbKLodF4ClMi+cuyt+03eeUpwg
jcFT/lQQXLs246FSXVvZH0NqdyysRmWTiB3ucyzAS5e61ES1ndrZspoQvprdGJkJWiN+rQhYawj7
0YpAqJxOUG6bQR4ykt1iX6IVgs8054QfM3UcDzTcvVlQHrUtjweuccIOu3Ydu//FqfJqCWk9ijuX
gCB/nLNmSrp/WFgDhRSsyrsZH7Zbvgo+uO0kNc4X++TLL0m1ei4zc3i2SCcLlL9dcM85z5KjMHwH
uPFNWiynyCUYJ7S6zn+BfTT71wzoc4DgB5vn7RtUwZ5HGx4a93HpeSu3xU580ZfxqCiIWBBzWY+N
7Dcz4lGmNqd9dSEgs9drZvpjR/w6+fWOFlNELcoEwUJzn8patJ7Z9hI1+wXwEmrY6gVNMWzpx4Lo
pjROFF1iFD7G3CrdfBj9EhFarevEwGnQ/k9bX5xEMi2OAy8qs3sUyaZ4lw/anFnMjWGVB7ccdIKB
SXcpjSbhKYMmVKXpv7VRLqae7XWk3KP6SXycm+G9DHH5MyqVUiIcX9PSakNhUTZlVi6KkrpDvzZ4
WQf4GC0VcWa4E2PTLaHZnxwRFDrMl8eS0MOfGqhpDj5rY78Y6uL14b4OHlHVJo4tmmQCPfbBeCWZ
ZcdAIqJWcu9VXQy0i1h6Lmonj5cRGFHiinSIQGpoKdnAUpBs1E7es5kbR+ZrWa2oN2X3SZHQV4Va
3UKCDKCp+CsvfjU2cxF2VheZJyLsvnLOTywY/dqrU0HkXBX5kv35yPWFRo9LtzZe2By52K0UsCBS
c6fkBuGO502sEVrZj38e88ZZYPwZL5oaBDMRwrOhN+gCPG5Z6diHkeewavwabh9dD86yQAKaxADf
w8QscStvmGWAoTvdgCkgN8GDhY1fnEBKe8QoQ65m8AXfiIyQDvpWnNuvapH8PHzEXQ+S07ah2z9l
4v3dHAei0KnaemFoORNM0SSRsTOmFS+H/KuP7l7vrUelgPHSpoHNN+vJdJe2elSBRQ6ddh6aS+8D
pnu3iIfDiveUXEjuDoOm8TOvNP+k4djfcPDMNVtfLROerjDxW+SvdLwjNqlzsnqsL9lnSTCVn/re
IQb2nLPidxRvUG2ghkwgdvZOyxstqBcrP/VcfJKihVhgZGmKLuS0fx97Wvg/E7bTrV5i4NUkb5tJ
NGgkFoPqg54h1+VwYXalhb/bgKgOwPcv5FWz8vEd+GkZ9m7R2R3j7QYQ0MZG4xYYlLO0vCf98mPd
eaWWxJDwmUE5EnO3HnrWV+JndHHI/H0kbIdPD91gtgKfYI2pHFAAXtIRJXd1rJtTNhFp6goZeM0k
C9zr/c1+fOc++/lMc6qibEGCDTQ1wo6pmxCMOp6TZkh6g7HDdPk8nSKUAbTHpniSQc719ia2InGe
hwmsiMzUucu0mcgRBXqiKTlJLMmeStI1iezFu+A7DlhdevvHTeII34dwYd4ueOnAg7GNEFVup5gv
t+7QU0NtPbkY7P9WNfeJC2aZtFtROBXdB0IsQ44mFF7SdZYMPSifeqoVsJS94rGYhFCbYz7k4uIV
OgmtHK9blY7DSxIC733h9mOt9oJCo4Cn3qfzHU9E8859LvbkG3BSKJ5OJH1DxGBDhtnRljEz6vPl
aIADZBwl2wLawFWcvH+ROxQMBD8rSLVTZYpwCg+UgIh12KXLRcyTGjjIbXPdlYTwY7juMgAqrSDC
NnWG9IT6kB/97VnSD2WZwozYj5SMDNiE75RusIf1Nc+McDpJu42bwgu/OAxo8rh5qHPi0N12YxJa
Yml3swWb/wDbLZni2mtQFbEko9/N8J+UCpDez9Dt0aDrU+pDbydoytb98BC7bGqQ5ZsGv2fyz/1e
2RaRvYenQElO+cXJ9J0RZbmCP4kK3LgdD803/A55VVERiUKR+AfnW8WYRt65Ok5fKdYsqpBd1nVB
U9YxSQYWg12Ky+P3SVxJ9GeO1Yz4tZ5rpw5RQSh1H/F6zexjA9/hUbBL/yvGDyyfmhtkZ9aiLYY7
XHzF44l0c42QJwV15zHGSOgi5NlFAXd2FL4nvhLLukWlTiSCvsaBBLw0z2Hkv9Z5X+J4f95sQNjP
L+g0+NYRVV/mwOFAlNQuJrAts3tbyvNf/YFEFYszk/S+6x7lNquBJ+55IerGTIIQOTBJlDSjfJi3
LRXrYwu9QPDr5/72h7EHBHVCaFviabReEfQNwQchca2TGAj/BCQldjaOXMtYvoVnIkpnmp1oHrBU
j9EqS036AOvoOj8jtgmB3oY2xiBFzUTEQbHpvn1R2VLNxfBAxyZymAGBhe9IL5VQAlKYVnZjSdIg
KVclTD0zv20UyDZoD++A2snYWBFRXcNK8/SlK5wJSNA7oljRTu9aXHSYA0PgY9cchE0ciApktwiX
pOVETDK6GbTWCvg6sKHLxpKNp6+cSY0fY1lEoVLOA4JPHLEJzVGk956bTb1WmoDb68jmZOU7uo+v
AsTFGX47Y55HYRxkglsvgE0N1achIOOR8aN54OIq9u4S0yD0BhiMZrN8/4GoHPAZ9c4ttmf43M70
a4dsxbUWwStszlhawm4jWrfQ0r5ZV65cGgMGZ3qzn5WrNw5kE8Xg/4VJg+zKaErcZownk3pk3+MQ
/dn/qvWQ//vYPOqLsOrHQJDalYK305vH+hdyCbaMULh/COSIwWpwrmjDpNEk6LCJwMCIqbnY1PMa
HlDzPxKvJmPW/FSOjUu0C72TdeoDWq54QbpTpIJ9w3hvBdT8evbKfIKLEi0GoV6X0Oe1p0C8gin5
pZIFs++jNcvJkRkTel1/YKlwI7sWDmnTV2hU8oKL59ZrU1UlP3h+j1wMYO13H/x+i8DK3w71kYpx
2WwyRoS/uIzOtrZm7NY3l7o53ZVUntOmmz7P7js6LuJr3LG2yQqa3egEaSIfqgHnY1ngJMC0IeiL
6wYsTdx0yKOzCUegPYRWk6Cb8JHcxpZTxjDjADPWirt+JmgN3ejSk1dGGZcmqVR9ni+kxijXM2aP
freAtS6i0pK3OfPuZijpMUGuvVlgLWe333QU4PNCFJH0IRAFT5dRShry9+YccQxyoEED3/pCIHTu
bCadC+cGiFZn0LDqgn5Mls5hi3W/26n4YX12QLldJcHhZwtLnwciSTQSdVsbycjnmbEDr5yJknqS
OYLQjA+VJttlCDIKW0Cu31+8PquksWoCZAXqEoitBsbsxk27dpSMg2YLDHEZrtln3gu2KpjduYLx
qmOlJ5W68uENL58t7tpGUA99Me+Qd1RCUi8cReIEdI/vtkcfwh1VfGGsDopdsv2Ve/Fcg+vc60dW
Mnk9FMLMlOX4EMU8MGrQBLaXCF8kVI1apthcRntA22XCXMz/I/ULss9rLZ1bcS37mTvimt1u6ixa
5RMQH+NJz4uC2TTKBqRkj4ARJaGbXL0Hzk0EEQCIW8qi1Y2aSPeJYd5z7A5fuMtB2v1txQbrT3LK
i+XssWRTKXf1Dd9lRl4D3jDEDXrBcAH+6IGzlg/kl4zItwF4MRkNRIrrL0yOydUMbhRcDQH04Nxf
xaRv0q5wcHrTMox83/WNzlGPD4pV4fYLFcxnUxuUAGTLFbC+vAU3+z5vMXO4yVkfJRwxOwn5TiJD
+st8S4H7P26cK8AAHJxvwKbomqj6LhmczE+D16ssMZzhUFYD09DvEItDQU9WSgAWeXblh37cS/75
FAemI5CVyVCOtRyaZQ9vE719Cgi+x01ImlNJ+BS4hh5wNMP8JYCEUv3/7Tga+4aLDlAKRxGLEXiZ
4QArsW62RQFLOEoU0qWUdJd81/5nFtUkhjWSerNvYfN91F2ZoNC5+lwyDif3HbHapDOZ2ML35qqK
WbJfrhVMyKlVTDWgiKstSyYLTY61nREcLfE94739vnuJpAFfGJJXK1eiAZ4cDfO9SuY/lTR/jgWI
DwBIdpBFCKFzKUq++B4HjY09er01lT//CkPh4lYjZ1+po/KITchM5fSrBxo5ijY6UYSSK6qjfAFT
yyxHEglrnu6HkKLrZljU9f/l5icpIaNhZEzrVTZFLIxuzZU49qpwiVtQ4goJtEs/I5n4RyKvz0wM
hvZObcXpYi3cnaboZXczCPiwN/l8C6CmW4EI2EOeM4W7J+psiDz/nyDyD8VNLh05QdFQpQDVWDoe
y7tTDNfBxHvYO9dyF09kN/ZBvdgiBBUWnDuQcu6ugaBIWIeoR5tdUJDit2t0QGhccqaR3QaciDGo
2Wa0zEeUf/+BF/Jre/MahH/gm4+3Mwd87NbeJyuDfRBVA7lKAnriWHa+GGccNcQhuG3oEOVDv2M4
khtW8BKnNIaCKulL9cEytKuWqIN9UtSH4I9mzqB3De4Cj6bKDw02gPUQUYvDEug/QkrJBYVNtEue
oGujYg2jzSQNLym/6UX/UAMcQyu64DDCd/Jr+hJV7mlchE2V9QqYdLqcvmwN+at8Cm+MB3idbE/7
cmxYxbLdpPFneSJka0LxeYHszkvBv6i+EXwYYGfoPhsGerqXCiYpVidDq5pjUz7kZyWyo43gJGHo
AyihKRaRukwk2FkI1nElN/V95ft818Op1KZ8VDCgb/oIEK3xJglQDxiUzn9X0Ql8xjGjUd7VS4Ry
iFJXyxA+CjNpygMsqthRwkaLS86SujGCKmHtTDtzE4xx7h0RPt3jHrK90pF97SGg3XX3PyoxxOIZ
QqLI3YA9aF95N4FPBmLa3Gw5Y4OR0wrQFEOomhwOVx7Qn92SWgWEKD8JlbyCk9kSlKXwSR3WE0tZ
XSO56KtTfFJf/1jc7QqnY9evrgZOs+tXSsOP/hdgtWeBIEAvwFiWjTqllMkihWkE1NMminbOOoJQ
pO4vmiY+P1gJs/RF7GL+0F954d0rkZiVwc6TuZJNDNmEbzr8S6VpyyLkGtD0V0zRRQfPmEryLrsN
8fMKbSORCyldp9AuoaDyIPvP7FJnNrNsNO4528y3S6ok884yjzLo6xhzQvGhioBhmXJgUDr7Prkz
HFU4AjDCf6IAWD1bcojhNUyQvFpCvfW7F2hHHUqx2yG9XjXRgsQxFq3K5rq2Z+1j9t/RIJ4sBgxw
7ZmOk7ACz6NMEF9xDmEW8Dyv4atZOBnmCUmNIbwo2C+xBnYBJHzGcYOtCz2uoM6b5d+ycTIzz9I0
Tf8aeKrp78XgjyeHUJmAM8oC6uhX1qqCnhjsY1xsM6mzYMslu+X9LbX8MQFYjdICSyDINN2wGEv8
8QdRCTWhb0FQMU1QV5nzdkngQu79fd+OVZ5RA7B2bunvi7hI2C9o3PHw0IqdpUjSRm5MTfjfXgoz
/T3cVT352/md1csc+AbTrwr7uZCTMKNFrfiAWTmbcrU3MZ+2U4kHdVXa/nYLmM4rcsMAvrOvpdbh
rUMRm0Azo36nSoBAEgKoXpNzLCUqJEmMQ9Xq/WqFgftXrJQrVhd3xqibjOiIVAggwA0pTUN+v56h
ai2SFHhL+ijxGw2mX02RnuNL6MoqJHnWJNLbJbV1iv0a9s8ZWlqrJjglbkQzPspqR9jtPE+8fxZM
JLEQqd3foNx802AmXfFRZIKFgMBzosfnfqNfFq7OmYPcibFW01iTNFhIHa7WHHzFQ7HyeDeBVSgg
Gnulf5MvBFRhBGHm3ZmTPljtkdak4RlQWyof+QjzumFyicddughDLLoYTE1LsWLtD+jP7vxNvsBU
ASz30dgQTXdDgP2v1BbcupwocPmIOgtrG8a3QDeSBWJALiaMaEVF2CddH51TD6BhvyyLrZHPDsTa
NUemVNDj2Y0hSszg/41OPL2sZhJ0/JJoP0z0QDAdG6qJrCVUtEg/Zoagj29leed37Sih2V9wEBoT
k8jO33gq43rdZmBJCuO0O865+lUEdVTvGhuhryNYLXPos+uLCIk4Zijsexvq8PGM+0KvIqMc7/yb
u7/NTfYUpMSpDfq7PTWyxt0B6s6PBNy4Y8JqKEq6RR/EvB0NKAPL/IR3U1CLsloGTrMoKrZxaI61
ffU5ub4SOAOY+OpQKLd7dJl//B4BZh6tq7wtzjFAMNFxTJN4Tbpp/dP3+BawQIsYPXZ0+pWZL31+
QtwEzg598gSJrJYlPRB3eYNUwpWcckmHL9jBv4vvu0r8MN/kjJaJJ2n70G2ZKgpQuEPSSIrHLpCl
FTKmyJpyUVVZxbHJqufl7ieKDEtDtMd6WFwM21b59DlD5xI8COE4RAFEEgQwVlyfPoaamnzObiuR
bSoxc8fhZUPrYYFDNZxKKTItvwUgWfKFwU3Z+56pizlaZrN+Wc6qfeB48JfOb38MKqSttc7vVPP+
zgXRT8UBDnzJTXr1oBnCijqeA6iUyvqtq7UqrZiQDBAMKWoehZkOSJEg425KK+f3H2Jcnu1GIDiC
a+oMm5CLwPknr/A78HD7Su2gKQPQTDGHHCu0Q9369BVMLivq9fJ3+KQOh91tuGaSxCo70JybLEu3
kCecgJOlgdoAe2mZOabwNNTtsE2F2yt99Q9qf5E1Qm1M0NpBUi9z9XjL6flgEwmF8c0hrFukx6c7
8HHlYrs7ex1Oru0s+9z4qfy7nxiypZlAZBXJYkpr5b+ybW+VAM7lgvS03xk56BooSIBiKH/Hh28a
AMtNgYyL7KF33nIUFgGzjmAtgk7RxPy09GnUy6l73hWng6kjKqmpE93u6tbdnpONtgr8T9yGyHG3
qvQ4P9xQR1SFsPBUFTTTWc3dvdsrylwpgXo2ildIL5BXn1CFFEawzKP5ueM/+vJ0tm/c8RSHxw98
DpIlq04U2PKYy7KwxzF4LlX1X8qSMAMNloADLfKazm6RL9tP8SBJnQ8ojhn6M2vjAu6gn5Ud01sJ
YVR4eJFjFbCH4yGzGi5GH/3O0CA0vZcBEvHxiVe/s9s+s3+OFeF4hu4o9UlVoPY8UJ24huP25KRq
aWDdmL7iasW3/lbqzF2mgqlCH6dy/DWlJxCUJI+cROSJHqlYKTvZQfYL1l4HO43MpWtIoFTTm27P
mBmdmm+I+B0towBiUTUrnGDWWIhgyQzT98BftAxXinb2QlKiKdTFsViLj1q7et/ttJPvAyGW7yEW
nxwayIZlVyUxnNr5j+DmzSbSIwuZxSU0gdcswE8+cZ7JuEgqgSMiaFqtosMPQhngEOijqTdf7A/v
TfE+AINw2XrLtLv7g9ixf4hrWWNDuc9ivJbANjwzjy/B44Ssm1itNEWsihr0u4xKA+EexR+lEbrS
iAkkktgbVnyeuJY5Ef1GabEWYrL9d9LwbzSsR3lr08SgXxDcQ+FY9nxUXVqTrwlTndM5O3RhyrXT
rmBKEZ/uYRcLFxaf8czMT9yxHZVbl0kmr8Qa19AUHDux52Dxm8gmtGXLXahVMR1G5xvXGegNU4m5
3PIJHCjBfZ937Qn13c6kMp/jkBX2TQzUVS04o8Wl+R5Vq4adLqQhoXMvbJlKn/zpLhtgjhiEL7Za
P3gWhhJTz067MosfiIIp//Jxelmh7oO95aSPpTEO3szZlw9NwPfxNFU4oDTZw/WsNzWnnr7Y3A/S
WuZwdzHzyQfnhuQIYPPTHFSQIDEK58YROsddxBkmev9fhg9Yam+y8IYY64FOy+YploKH4RJFy1sI
WtAARBeN/hklXC++cKfwyaaFzadP34vpYGiXlC36eEma3lOhKIQoyJABtrgXJrEslfKsmW4BxUgH
ixTd2+biGMwJp/F+Nj4X/4+7iB7HLcVdU3To9k+duWYNbxZ14Rx32qD55gxBWUn1JpcQt5eIlTLA
octc7jAC3lXaw+HqSyGy+EfgIPcBwy3HPrrgvNrp8xCCum76o1SpLBuvpLD696WfGMxDt6KvqekZ
90bun+5mCRTQ+N3D47RVXeY7f7+NJ+jXVlWXcnKUxuS82y6Um/K8e8fDnCDYjkcSj5xFnWmHS/nG
NqPKW+uPKxbjXrbEk+c0kgOCZyDWRW51k81Cdr1l8H7oleo3EvpxerQrukGnze/Ve1jHzqgRCKzQ
RxVVcIuqYRDGEluv/R9JGojux85pK6bS5iRMOfAYcx2h9mHeSBT4IGi+uhRNvAMPX06/iFZGpPD0
QnY6eszMrqv4awqR12EBum2RTkdNBUc++iI7BPXm9mldE+V+KeJ3XaX9ZLtIQrzmaSo/m/acuLg9
FP4w3N4oHGYNIDovbn0n21DkNNAnbfPh4/M4gnNEzyCHzjntBw7lnZdqUba4Z82yIFJ7YRb1pfR6
xFTYiPFX7R7/zwUHIWVONssC/UpsQlihx1n5j+FNrLwrhfZt48sfU3f6iajueZeSmn/kWK19fSRV
bc6u5l1DDEVHThHNywyneS8ur3XB7Hu5NnqNfKSshlfUM6zh5ZnVuTdo8zNyBEEwT8qbhVnLa0XO
fEUJ8n7wCQSJY7tMupR5TrEuFSbbAcfyPNexuxtJyIv+5cYAJgH3e4/mBAKnM6bBPlM/9/HGMu78
Zd3jdMODy0dpfWIwdrx4GibCFIZOZAufv0qrl3utlb1nuJDIUFlSbXkbaiwIW5d6nU0CpVAY8kbS
gHjB0XLvqvDDClvEQI5xDFRZOwG+lXbLxSAdstKrnvGxouE1lRoKNrhdndC1ERB5JZpXwuCusGlW
9GzClSJpRsnT87THabkBUPG4U13d/+NW0IzqAh8svENmhX1fmfk2U3XyyQ3WtMgkgAlEYkK+3rFP
JtZqRL5D9u772U7NkiBVBFcXWkBODgmVnyFr6pDkpl7bYpB15rICUXa0fiQsovfc1gGw4E5CBGb9
GzCR+8HVWcIeaWRozEEsnu6VJDedRixOr539OaZQcjQ58DYS5SzFEqKCWXivCUR0A5XaEAlUWKIK
ZAk/bMjJzM8MIte8JxJR62xLvKCQCEn28Z5uMxtyp3dVDpxV7+rPPWc4giTTosHzHHx/1nyMWSfC
BUizTvI+mzo6nhmU8iPyo1xDcFlxthLm8wPKX4pgM2U7Y46v7FJOC7bzme8PM/ftHR+0vbYRPG/j
INH4UOXzHxFSkq6pF7rZ+qm3+9AnJPJY67ZbaxEE2M1fWJTqqh2IGknmzDO7BwJHz0VgpdDiBjb1
9ZXn1guzzgksAmq50j2oUPEjCVLvBIhvwZcL+I7tSUaAeXlpRCHsBz0AOOstql4x4v0yLbqSsVeM
a4J4xEZAjL7AgMJUZivU1wQ0xwvpRCsvx8m9tdzngKteAiXcyrfG6/r5IhRyT0eolgmFGLTDKO25
+FVnjB1BeEPGvNIo7rVSCfDa1enKm6YF/qVtZoHZO6Jvf23KPYzj3hT6SKlbimC/6vfAjptBTuI3
NwwFa6Ma1BK2+WwsmbAlcSTzifYi1U+y0gwo7KJcwwZBBrKTQr+GIaZQOjBUBWzobgaOGjUnL9Xd
fPRU01uG2Nlg1nn11tmw5j43nw9uhC8zKwd3FFyt1naMQxd/N+mKE8m4VVjFOjxplccaspsu+wGw
xIF74vgsivnSTFxU8zBZ9rTiaYCnFTshj1H1DEqZA5RDwyc/2O/wGn0fHqsMx2bxK36Vc4ttwxAi
mWgr0DOD/iiyYbGJZCv7CPRlQs2O93vSs0ld7lOT96gyIq5r8ScUJuPk3bFACN5pDVmPlmR+bAF+
MQnkWHSSln7b1DO46I5H/bcIcudsHryKy8Q+EkGUJbHi8dUjfF9M4WSgUD2TWTfi4K3q4gU8s9kP
Ly9nYO+jR9l4J6S1uFgACV1bc9tCZkmD+PWHNc2aWaZON/yxjw+yQiFue4BVid6wFE3Yt/Vg7COJ
aKLws/4DqARgWz8C9xAarJwtKEDAN0uhnqTl1Zwjnj2CsViRc0xOHTaJycqYvBVs/xegcAihFGX0
qrJI68ugs2Sx4/r/2bp3CIQFXM1rjqGDdgYof71YlNJHYbdgfFp14MkDB70kRXNeYAk2WDpkfFxh
yvPuH5t83iEhUhri0pCWUwZ1ZSxMLNhTYPkSLXI7rP6W/M5pwRmSh2a5vOTd06t30bAtzbH91o2S
4BnEfkJLeXLl0+2uLvTR5OZbdwb9XCFPJCGhE5y3Q5h8jORNqXzE4Trc13k3XPTXTTmn5vVAhEdP
o0oBia/WUO6dnkUaN3/JqjJ3BX7R+wFLWbKalNzMjoob7oaVD3i5qASp2YeONKVppeCuD663lCMA
vN8g5Ihe3dmTnlCpNRQyl7sdFbkErBFOb4U5id7Ob1ZwIXekOp+AN4Gke1iIijs4HzrLumUX7rEz
8YLPz9fZ8Q08hzSUpwXC75U3PRU8BUG9Kxm3t7BW/ptA0K43qSP3mUYv5rIIjtqnyuqwveJncGZZ
/LiZIomLPA9d/ry+ec0A0bpuvednK7a/CxdhQ0kfK9qmkyY1ziauhmNt2d/jFK0SJuJJObuVA3BT
lS7CJU2sSKjS+MjX4aNTVb+NS7BA5WyiTamcPUNoRfrzQ0ENwLa6K6onBk5a8p55uJgRKlQy2ro2
fJhs7kjki6bUMp6jwowqXmAzdX6Ct8eEY6hXJ+00YccHA7X+CD3nbXT64qW+4s6tEFcNrCTGwpjb
zVilbqkQZHXD5Ums1TaBRG3b9dFelSCOOo4rgXmnZKGTJT9kQUumv5uKwebLnVSx3/qbmTuwTCa9
R1j+xgIEWM+IJQayb97cdwBTQU31T6fc8O5gPBjMm8CtqOX2AaOaBOYgbODoGbepxtZlyEu6G6cj
tNkOdj1i9g205zKoxUgS+Hrx8VhKe2Kw0JszVID6nuZuDwXgApyce1VqQtMRD4vwe8SA47VkrAd9
H54y9sI2MdCrCViQyP5CrrqhATux4JpWZwYB3yS5uQ3mIDTRvchc+ZZiZXv142ckfGNsVdg+8aAy
LRwUBm40MBuaLvVpM7VU0ybLpV3BNfdxiWYVIuaLz47DSWuARBllH7aIvXO3w+jehbUUyh7D2j1P
ZlkYDoC9qMghIhGXVRTxK638gizpUbrMbTvTpNRzbSLuBR/JCMjMMojeGLY6MuPMkJJklLbAyYyo
WGWUXxWGm/P4MrKwLNX99GBrZajBVSluvdCF1M627vS9ksaZnOKtiEPearzv442yTGbbfZj7mTpD
RVQGRhC5Z8U1QfOypwFe1YpRpafqSQwkOYfeYFRCRILr4aNLYWVDlYMEfUFlP7CRHru9z7FRvpWy
CESqSchHzoZMzOnfFXQhOn8n73szniTUgGwoFRvGnPv2CMnSFI+tgHOm5yNhXFK7NLoNfGSoWJ7R
O9aswV7n765BJOHrO7FEZdzpsaW9FRcesx4DDSgObgAcGQ685vF5pHJFekz78CjJkN24zm5d+UNE
ppWW9pwlNK6YTmFYOIJYU+hpIQh2Ps1ZLk/ljxfncgAfsus/96djHfmgscDlaTfZvOjrxM2Df3gZ
xt9SLwyzzMId/TcCBT4KIvH3fabK3N2SxRuIqAQ7OZ6A62nV/af4HQBux27aHhIc5PQAUZhZMygy
Nu2SBnrP+paW1P0KUNgibBUuqzaItaaHYETaxamt4jVfBUHcUVH0XgusaxqWcbH8huncFJLNyXZw
rsovxzEJCQ/qMubx3MDqz0kSf14PLjdbSxSurxp/GTexoVnIMBAA723wIUZE3PYw0KlXKEccRda/
qcXrWZnIi1D3muBTBHDdFW0EZqo7Db8oqnqAV6AdG6ru5VnU13l42tOI9OWEOnO5HFTYihEqGAJm
Bua1bM8BjO00lBMLaOaKW1xc8bqjmhtpW/SB+jGgvLfFoMZHqDS+esoHGYyaYp2KINzHOGY6r4SK
4VITOxQXJCqFNTCF+CzVytTeEmgiUUxCAhWfedMhm4sQDqAei9rJPdiqQT9ttGweX1q+jgkmlZNf
fSd7bX/pAIkuxK9qGAJcQbq0D+AZoAuPkrEQFaPTmbKwTE4xB/anwPIVdZzysU0IHu7JowQxNNhf
bzkJi3EPWqfvQi/uAhkNKyoJViiotAKTFMmCQAg9nOPG9jmLklz09oQTjmntxoxlBIbZwWahX2+X
pXR7vvzOeGl6/9pyIcfyYABQcMAL+PmJVi4f+1DxyovPlPRm7Ql/KCMhegdDSDJ3CqAl707QGe6K
LB8ZWsHVTUFkswG1ck+JqaBrRwzAq575G4J+mlflnXuQUYUP49Sr+O9jgCNq3VS81LGzaujJoMGJ
23J3Pbml5VvaZRVHm31UgQOHnddDueW8NbskyVMef1q6rtgleNyVXlGEEbAQsW1ODHKnRZiYu80f
aE2Gqu0YZ+Tdo1ZTXGqUClCPYaCjMFO2ONktk5EDN9QPSDt1vLKIYKo4KvqiRCLCTNRcDqz4J8Bq
8kFOvP4ypa3mC78/aTXoAVLxITOxqdvwFlFsUNgBWoHWO0yolzo3HS13/1wsppbqjRf82Dqg5hCg
iFnkw40mHmCTxVm7Agp8UTSuCwFlq9GRcCxE7+rxf8AgMEdcSBgBYZfhlwHU1wfjnlcsA0QitYLt
eTG5ZakQf5LS73zSJS0tsC5bQ5JncmZBbgognHaXvoGrtc4w1MtyS2Vm02n9u8g5Bnzn9AzXb1r/
cmvQefK8+0Az5YV/OODa8Qi71UqMYicpAuP8oHE+U+tXrby09R/5uDjoxsektcS2nFS9uU7GmgFP
He+JZ+lGF2MnUZG+VEqM75vu6ixkBtgTBbmB4f8GkxEFqeT/B820FvZxXVxxcTL+2Y5XbBArV87s
p+Z1f+z4hh8xhx41xYK7nYDnlInJb/xaUSe/FvX8P+GzybitjmaIqakFA2Oa7SBHR5RhJoRZz3vZ
hYFY8etsJoSPaO75Uwzs5t1wH/nyYtuq/tFX8klze/VHjEgYxoG6pLt7FUaA9JZFAB1zQeX1evJc
stL3O9jv97dM7hRC4HYq0IGVEAjfVbJXSP1lR/CxDzV+ypTZlDlFbehBzGmYpYZlcLY728O5wUOK
WgUofa4YZxrIz7t1H7efBHuGDtTmyeChAk8KYqJ+uKNUB4erndqPQ/dxLBPA+3rVWhtr2AmmIg9x
YLhUB8dKCZ0UdbVjk0l59fNOA/KAN+t/A2tUzQpkXDKFMebV3Fp45t6AcgMgOggSMhFhk+FKefiv
tI1QcZ3gI7jnAwq/xm3Q8mI63ubHv5rY5+0tLqDx5qJ8cGakOUDc1czjmmcA4IOpbfZqGoERJS0s
jC8VlgtU38zpNRmjeaAGxyfDTlCq4I4ZwrWRml89voMkSJd+C/11jo4y1VlaF18x0HWHGUZG8LDe
VgT20yPwMqoOAbGkzn3Haj57nIBzzCNIcVQSOgaGHgxbssWekjijnsStdW4yZwUu1gOVZlYyHjgQ
HNU19/KfrE6hMYN4XL/QxzV5z2Eb7/aKggW+ZsAROAK9Lw8Hvj2e2d7A/gz3BG8kthAdPiySybDH
VF09xI0up8g02t5rirvZbONsopuLDxgKWd3S95KHwiHyTDeymmSVg5d6Ze9hdvTYiodEvrhjPShH
Yo9NmMSuvklsA6KM+jQ2xx6ZTqJlXHG1QsOU5uNAO9OpxmtKJW7Kmfk7FS8yXahEkffwO51EF74t
3taGfggEjNARiEZOQ9P63UwjMY6iDwznP0HP4tRVUvG2Xkw8VYFXwGxNS6OZLaxgA46AbCBAJQK0
r3veHLHiTE9Vglyx0T3ZmyUAtPb0FUFsQ8ZeU6VWW3/3VxOtz317UKTrGr9uXpcOFqcts0zXe/Ph
a/7Hxe5uH4PTWrTHIqNrB72iZGwGg/tFYlpADfo42Rq7Dsr/b8Iyk4FSTV41Nw0VRIvgKug2IVHO
YP44h+HxoD46qcQOuljuTYKa5h+f4fdkIUZ65dvuLUeVMk5lNNChKpnvkrAZwVFpV37PSzu/EOmc
EXXuplecvGhaMPuNk/ToZL80mB2edFaoefl+wcuvbUXCvSg2vQ7iZNV3zraBnViCK71i4lHUswS+
oU4+bSKfMKTf7lLZAcKIgfqYT5YzuPfvSUUuMyOrgOenuKrILrmXLUynb9ljuqHWvt654jQPZZZ3
F+hJMy1qk0S22nDlPbWeYH7YaqUWRhiFmTpFsYcwGFrn2OD/b07GUAaMQQCSlCi74bd1NETbahy+
t1yVb/zIpkROBkRX6CqfRnj9msRufUZUzvfa/L6dyF8ArD7QhAl0rbW7IfbpyAhIpAOtk6XLiMZt
prDr1nzQNSjifB4kDK1LmR/PtAc+vVKWGDMLklSo/AFCQrYmbiYjcmv0+BPXXHct1lKQSuu9n00d
PWLpt7NU50TsWnIlAr+zdKQGM7KGmMqIJe1wMrG7RNoDp33s8Rzbjx9IXNaog3VVkdr2a4LOFpHG
z210fQEduGiWQbNebyhGZFO6lp0PjrUi0wlmQlkEpk8wKZXEwD1YjU+5oT7caXCTmJapzlnRYP0b
n/Svx48m525QiFN8ecc0CD7huTtydsAQQqMyEIUwldOXdpwccvuEmey6Vx+SD8BIP7hHZbrl7mTU
mEZK96JaEKr5pyDUOMNGXkr7ntxZ3r9DOZHjv0i1sfkSrbgXR1gjP1983RvY8IaV3jEK4+yNX8sN
1JiI6TAAzHUaxAAqZETv2up/D1mKWRfmJqmqhEfcs+mdf+ognYPFZhiJ2/lCd4ZAJFGmzTYQbgvD
ho1j1edQHZnCRfbtDeXMwkpWfZvtOud5k8M4v8Hj6ccovj6ddrWW+kJasPQjLawMX1EySqJ1Q9CC
d4CBQCHKuygZgQ3lpPCj9OTvQLApq5hawZ5EBHm+9RBixw8eIXvk1hqJ5xvXMxfuFHxEXLi57Wag
ifQAbjjjBxKqScAagKfNz3n0+a8QCEvL7eMDsozrxks8Z0o88Y6ZSPkimI+Nm4xnZMui4AoLJe3B
Cz4xiHdVYRXxQRdBuZ53e/yPF+QtMX5bM1Rdl4NnkiyfQ/L/AdpmIjeAKzMN2+lLbIEo/1GzvV0H
G817e49XVFei/xqP7CblgR2mghpIGazH/j2ExIHIx9Ha13bYwlCEOghEyeOcKSTDPFIS5mwWNS5S
BdbWFkvvwdDv4ql6zIhEYE3ikERurpkcKKBgaIy7damg18/6M+3EM2oyl1pKQtQ9yIV4HxpNLg4x
YkEisih1g65LY1al/C3YQiP32MPzAA5chGObOBjfHRgZC80WEbs28bAiQJrszr/6przfZJfuPZBE
vLW71QgGrkPD/uCXEakVF8NW4rH9PaqVjfda3+Hh4HgO2qqpa+OdruJEXqj1cXR0LJuvyyCA4F3r
DGalAfYO9Bb5qtzy3FyWaEuEmEziRmOabHIZw1O/hZ0stJwHGewxByiHAHEwQqa6ZzyrgaqZYuCf
OX2OtSdQ8n2u3j25NHnFUu/J6drXsrER/+lDCQse1z1Bj2WhNW3Crzg2Fw8RhVijpc1iFxw8cY6d
3Ru6jVd7zwQ6PeOw9BoyqgN9s+BRtaIVN/ZFDhFynXytJlOq7TinLQRiG75kjjU/P3/wvB26ks/h
ybQahGFFEUbOMDD+3a8jQZwWJOyLpRVAEbfnrKoegGZC2XR65HhIZmTjMIE9utE5Cle42fksESXi
rKlLRZoNVLtkb8yAVVJ5egyA/xDhG9U3m/lpsmBoR83Y1k2CNkn8t+hbkIVTjxEPchfoAW2R4al1
nIRlXZy1dpWPH90Chg6g19Vxaqyt3pwZlD62I6aJZe1iGaJlPN5nba82+r0Kb52JIq+ndXrq0aQj
F82eUtAMXuHOkm93hFCou9RsCNhNmtM72gHW+6MIB6mh1RIi6pXBUDYBMii+mU6aZqWXwm3rgOWr
ex07XsTZir5aokaIAmpm+ReQNXPpYughElkJCoDUMjbE+w+ZbCJx5Pdv/T2wx/gtBtyN/62fays9
CToiSToUiucjauMsWwUqvcvMn00Wzr8XMlj4+B5iL8Jf17glW3XB0lxum30MhyPGbBkIxwdCL9/p
8jCKlxl36qdUVsEwECXH9XM9DnMPwSv+Tn4+cZ0n71ZAzbhHdd9O3VjlBX1IycpeEN9G4XYO+Ct/
N2h2NP+pTx4IT6UHQlfYYiGA4GreJ69nnD36G5WhkzLcqX05LSQL0SQxCU2u12AQ0rslpxjTD+2k
fmJVrqyQHGEaer/CukUuc+erjqYhk+aWRVRLliCJG6vlqjzAeRb0vMR6Oa/ulP5Iim9zjTQ6LXyX
GorSmfIuYqbyuDxqscEvyUT31H4WjwQJ9p0WsJV9oj2gjlkHOcdrifNHI22QuYoYX/zWYCxx1J9H
6dFfkf5m2SWbt1E03GxyPZfcpA+6BEL4nNMx+nYEbeluCFk+lrIyyKiJ3xFi1wff8uYO5ZuPMnT8
pMaLv57hNn8shhfgclMJ/LCGttaoLE/sOn4Nyf5Iy3AH8meNxnuEQFpWp6PWu01ohM+n3qRdY2v5
BfzgOMFoX9qGvS45DGs2CylzmecIy4DR1Rx3YXPzfz9qzQQeMqAWlNiJkZHL7ObLvjJMsvhWm7w6
5afHLDXgJ7Snl036D/vRq4swCDyCcx4L9HS+pNWf430mefqBeNoymxFvOxnF7MchNFX1nhbSS/yv
Gf4yFNqgSIjfFc862do675b02464jC05870w4/Fw0/NemPkewVjie0AvJrQGBnsHNjCE0FDGWfrw
t8v0bF5ztCawijMaVmTv/IZZH5jilCJZND3Vh8jetJ2DchvNaQQwxqJjbaRH+uo0Pq/stfE/3QOX
lKB1QRjJFOV1AxTMd9HYGNNlpm9/r3Esc+k3H/7F1Rykq2HEXJ+1w93+ThBkUU56c7bN3hn+nTSy
qwJRNUBzEtSzHf3r/1X7vE6SfevWlei4+L+0puwJLASyqw63QKP08PaRAKNH6Osil2bk8gNUb/BD
SMMt4HmAmqvI9BTrqmtO3MnA5xRzSxyhBuJRiVr7btGPx5OtnfiHkbP8vn9uPaJt9xdTjUCgRI/T
hrGKGTwl/TBK49vFqofzW9F1Jy9nQnqEZf8bQXleYVZ4glNwjnlkrqoOF0zvkp21wqYWz4WzoEEm
iEvKkoJ20KnPPhW7vFDxOCJeYUo/ekl227IXbrRjjK+VSFNaZWS6HCd4KIBCuQYZgQU4GnsZJK9t
PLhH5wBcS9r0KH2DvsnKYpMNB/O9Br94AR2gU1vKPSZqmDr1EayYOiKJsChq3/H9Z6VzaFIM5c6Y
eR3xOGtvKEVpjxgacQhSSnLmlczh6b2cSoVA1H2/ArgUtsTT/fifOshxF0tqKrc9SUGhGAK7THNB
gXy/noDtgHPCPLc6zQ7g/0idnwqdUJRJ1mnel7Z+Unp0mZTINj0EiekrmT4MSsT/0qO3q+9aXmfr
DiplumjfXaiP5qNsELCaI8SDEL5QZFT7OtfmM3SOKp3Wsvl3ABbuSfpxIqpN0a9zk7HuzYvOWPl/
45/hSD9pLzhxFGbuuWKwNMnglI2SzsmK2TRKQfCdVO4Z62DF1+RSsPYfXNqCoX9jPu0gFpsZNyqH
KtdgufVULTxX19FzaYlrmuAiDiapk1eEejcbXlCRNAwJWa1ae6zvoRf9L7eH+UIdniajbb27AuVp
HAm4f5NCkTZJa+mwAnTd0K59iGqEjnBLSouw484pGLDA63iy6SA4EY2SoD2xtjLXo1QHtCFEXIry
UNpt+A2KQ+fSmsAv9a0jSDMXUo+2LM3tO5PNnanW6zykmSXD2L8PFwfDeGl2dlQQM+aFPsHT6Jwv
D6NP2GHil5TRVqK/6JL8GoHWiziGEWDkgeJRXeNzFOh3/3Ud00eiA084h8PHTP3VS0ffHnTp0MNL
GK3x2QXE9BW8uvfNX1gxdq9YFbRSipRo64lCzPrdEYCeQZ0T8LzF9cMcbqcX0M7RPgheGISXx54T
nNGHmbm5e6ez9n8w2VlHh1OtgtqKgfdcU699WUlVgINGy6YBl990Jwh9C2PFdKd7R9g4meDRo/iM
yVRwV80Mrwax4o7dwuTGph8/IGv+0NY8Ia1zv9Es3I1mPlW56IfA0GyPYq/eUR0lutgBfnEHN0Rb
qZQsaZGQYBm4Z+nso9e/cGDg+keHKR1oCzmyAWP0ghhcUezbAKlPy2hPZ4DZXgbdonhvkDEyZxN5
bBvqs2vXNn+598On/gM449KZ5rFnEPcIfZSLHy0MeX5HWyU5DD0i0XycWBiEE50M4wGzV1sbHcy0
A4wJKEWI/7ApaHfLfmqtOJ767BwcEFZgjv2mJMpkkYskNNkk7kjnksq8mwMmLGV0cgAbHJAdfSHN
9mJkOonGsj6USrZkKaT3v2AkaCWyxwO4WfBiWdne1s9IvU7Bk4wsgGAIeU+SU9MPE48hJdjevi3b
GObvFnY6wsiaH/YMzVwAdUVaW0/iJLDSolsRY4bxkSYoWKpGSnp4TM/I+PDHsNbBuUfEvcFdz1CD
vSwRltQshZevGGXulIWad7NkSMB+8svjCts+VQ6gUGWCQwgLBitsC6RWCa778yX869PlZpQy/q4C
F8PtBsK4mzue5fWWxJHycLCKGU9hZIc4rIXlUC4gPy0cfOBsOcdHtAPqUTpTgGGEIOv7Ig0xe6Kt
ul69teMW2xoHVfT/EExpxY6tWBlDgmWxHLT+n6KKtfFtTrYDLE7x0MH5Cx4Drjrd/hQnkIrosjaT
PelAjO0F2SqYc6HbMa49ujecmgwqXq+mKAixQylTXj8Kdt8JibOsmeNSc9fhvdlFmuqYXPsGmZ/g
totza7JJEsRtJsTwEeayTiEYOcK04WhlpPMjOlrniYCDcWYYpCdEa1RPwoxBt07L5Y+OyRCYHq9k
ap6S2OUN8FW6tdN0LqI6/ELjjtlKW1u00dV7chMizWmYjbxogAVFZXuTFRHw8MVhDWHVb4Icf0MU
DxEyMhOB55W60rgVSWV04nEZ9J7tOV640IWRY2AjArb5UIJXFu7103iQZ87WU580X2JVA0+4w+rG
eyQZxTZ069nO8a3vLoXoTfrzQLqBdCdPJt6WIDX3cfLExbhW7S6C57uLDyurOlA+HaeV7asarAFD
nLIC5E/RA+YRJwsJju5ZQkyEGn8Y0tNlAPiNwPkFKlegvmRCCaIE4kjn//UKQumkcKEzST8wXkis
+AOgagYf8LEM6PqYt2eyea7Sh01dfa07ew7ZrwDllHMLHLJ4oKcrgcPZ8Loii2pEowbrzkv8oknc
pomqHk3FjYaDw7yV+DBHhGN6UVZK7qABrXC7rVMifxGHgQpgpxNSUZGV/acuj1sgb0xq+Lwbx9Fl
h0mmPBohc2fHhC892ygHVPohsX8PK6MhymF2qKi2R1vJVJZAi8dL3UyFG3Tf55Jp4F9S+byKpEfT
uXcRgCZlLODO9g6TthQsIWL6rHsLfTPFvz2fsubtk0eKA6xOf2avrqNgJoCsD9HUss3g/0yT/Y/4
xu5A4pjRzjW6MTQv9XvDUsP8ffZ+eApguDAcTcPv++/odkY/X+KjTCogTtUVGnH0RFjiL4vB06Qp
9XXGp6HR72bJoNGoDPvoPCt+XDX+Nfvx61lr52q5KEdTXcD1N/tprM/x0lYUU6VK4qGj0LMmk8MM
UFYkpQ2dlR14HHB8at6jIIMGOHh0aSGQSYB3jX+bRJ1O3gBfdEXYbCoeUN4yHKHMDqs7yGZM8qU6
9LjApDWKGaphVNS2hq8D7pFK3m+vlbJP+A5vO6nXF/SaX8BVDRhxJIcHkDPdPExpQ2sE66k01+IH
bJKePC1SKgz2h1R5ajNcvGfBNHuwP1Qhkv0l0TMUFY4CKgYJYa294/fBGte2rGAhK9jWLEx298GQ
6+Ot1KfFHH1qe635C2cdNHw2HyI8TBnc/LBVC6gftib21xl4GVxEStjtGY2O4jN/ihYUiNIPLshT
xsN30IMToyANWkryo5MuEp1bKgNnhJ9mYrRF4duOmTBG5LGasTSJtOWW80wk8r6BiXNkR3EJhfra
4denr0L7Drei5dhV6yN0vVfpNBwkm/eyK44J201C38cAx5yV50NUemOl6pNg9bRMhWh6YShMvVV+
tSV5KINAvJTwQpfODpc0O1rkyvCmsw760XBytNCQeaHsiSsklvbwYgyKvj+1vTXbADrIzZv3Kkm7
RNUDOw54fRjiUOtHUTbyYQZ+gOT1L1ZgVpSU2g4Esr493el+DmozPITfY7x5eCna3nVBc9UrnMzW
Rz8A8owipZ2uTacYnQd/hqrujdIRL22Ih0XJv2JXmqsl41COSg8DnV8ZDyYY63xfMjSWqwCDPRA8
Jsp9+IqC9z7dyEvP7kNWQICbT2P8BEHOj3ZbpIlM4rcoaJQSqeDBEmz9VJ945PdcRNDDwOh2j5yn
LzPLPT3aVSoa5MY4tEGJv5BjDB5kLTQWs3vlGftWGq1lniVmS+cBnNXUF2sxPI5U6kTNT0MFG3OV
5BTKhuKQq4Nc+4/8BpKx8/YNajj1TZbAZAIpK/XNK9PehtoSYcHARRYMztXnLGxEqkgeyg4dnUxk
JSt0IYd606v2ntTKcCBlhSlI3Aq+AWJ+YHQozf0zehIZZvHXs/9u8SLvR0ueAmnmM0cYs+3VJs+L
r7EGGrwpNuCAh4khulkkRLzuIB+iqITXQJ+6LIEn1YTi23c6nTf+sdh9LRZF+8ChOGjUlAdsnlXh
XS8rd5WBmeF3pa6+T1hbrrM1jLoPBRZn8kzFoKwi1+Buyg+8qHBNXqe3onMqsZ65iy7irjbebCmK
Ez2R0nI5WZgKtA6W87zEwzsFxN/ULNTb+4Pk5DcoROLSvGH8EURKg3DDv3QS4I77uqB0DoHDUFzG
IhBLTdIzLMrpsI6mBXt2tsJxVYiShMVlusfKpMBUJrWrKpcyVkHKmfeRalN+Li+AUMRTTDAkR2T2
yNuWG+4ZzTSUs/fXgVEDIVv/Xjgr53Ih0cIN9C6ttWi7AQsXx+wP+2FDry6S1mrMc6Rzl8bYiOIV
ivvTjYO5k9yp0ZuSUQ+YkUfQpGqaNZR5I47+w+dGBwEhJWVtdqqHct8lIionn2z1XwtU2V8dYAQ7
npSDHz5q6Tv0mvnHASSIG8leUQTqhFZVsKIiSNNPLzEGT3R8HdMezWc1uXGMw+UMBSTUEi4zyIwp
TqV5KvMqiDUBd0fxiEqH7wPIfT3qTgMYH5GA0D8i/t9BzHvnXTaCMk4Ubv3jv/dQDJm535B4IiBe
3Ypreg+sqaNWNaIQIo8knFivH3z5O7Z5hyh+6BvIVOD40XG0HId1i8eOLXSaipqyX8guB4pBafFZ
R5JnqPaLeAfzC60IVkSCw1Kd2YiGZbi2+5c7mr6qRalif05cQhR9E4RNxkdEyC70hhBSOPqvZHnw
3Wv5loT7O91H7Z0zGzzsN7ulwwlktVQaxhDmk0YtPALIifhTEsZifi1kbVf5+pJ7FLgZSgqBxLxE
RqRbT/AZzSym5GKAYZA4usqYD1TdnyTWU8KiAgnKHjhKGvPzge3Xz3FCrVhZyBNrmNGE0CmT6mCw
XM3N+WJn16469ELNPWy5xnSPJmDoFCrDp/5izamuc7gVLPrJywmtUjQtSYrXXXXWs4HxerI+Q+K+
C4Pfr4hk8N4uQm+/iZwJkP5SdOT/pLFOpcXSrBWx0NoS0IqcFRUJUbyVu1L8DuOmQnTqlmzTYS6j
WUNIXtIOjNMrwoedqktj6RC+3zcmrzR3zhqYrWIEP+mtPnyv5nMFJQIJtLpPHBLQ189a8u88/eAp
YNndNfdGGfjRTBi7IpF+bL6Fmb5SjBn73JrCFzVRKp8eUw5yK2qWF4ppm0CzulJSstgWhxvk6zuY
zHNJ1LzKAp9Bah6KkhcWmV/xayYWyWIBWbWOYpCw4xe3Ppo8SAYLsd+OtxArwZcYrzvSd9KBMRK7
nzuYFHYU/bC2pnmrkBY/W64MwN8l6FEVlGFOx05AYcOFjQw46gRlSVi8uCAX9bz9PgbyMfUUTtVD
l1vqC97utUBHhQl81PqBKhpz+ZO4QuAXNGiTVQSsLAw7XlS3BIrjXMK3pWeVEQudjgdayw+p34I9
z5wS5Lpa5VGl+GkXLwM/UNuLefDu4XXp/UcFeCY2zygycui16Gfyhb6q5nB+Gj7HygBhwYsgL1Vu
KrqNOiQJjvrXWxUfnlKOJ+UWvNFQxhaC3+rpbwEwFM31sxc4q414qFtsDT3hADMSIi67MwK9jqxH
CGqDEgJ0B/9DL3BafRsQtKwCViI8h4EhvhYwRx4MhfdWWSrNpx1ayQbPrHR/n5hXn5cm4VS3t0nH
WmGo7aPoW77nj5SAAzT4yQWvixT9DUmweSdq1dP9lAum/RfobvaLBzd+NQToie6w3nT4bO5a349M
xQXVtACw958kL/EebRaquipvpj1KPwH94/46SICI5W5bVNGUsVrljIE0gTduJkhD17jcPcgrywQl
Xu/T9Mt6DrqWVC6fGXxEVxvRwq0a4slrPrpoRls7wgVw+QN51uX8sNSXV7mMh91ciNH9ogapDz1d
jHZ6/De9aOBUJIO+X/kSzHHd0pHAywH06jQyUteokxunWAntrq40og1Llxmmzm4NRG05FE2ywaTp
WP8RmO06n8pb2DBHeZV23D1wwP3uVURLRk6et0/4FplvRyJL3U9xop2hBR9IqL9pkFgyuExgwl4+
5qD2z7stKlQvv1boqii7N64uKh54RWi6XazvXnpzBK2p0HTXh7lwCF3liaAKcNdoFyfgg3P/6Be2
iUOWyQ7eznTymUnZC/HsqRU4v4ZPTKdj+X0onkWUWVQf6/+ruXD5uzb4TMqxWKPwapR7wt67o5hM
lZ6F+JR7sn6xPtnZjK10qgjwOB5yf0R8LMupQO5LfTG1NXfCPl3Wp8oJlaRYFIyCNp/XqChydeGF
4eqmLjlEWO2xjbpY1ofIDy8xpO+pSEG3BfE7JN4Aw3tph962Qvr6KdUTO4veqYINx56SEcfVD/Y3
6djLU5QwUIus/rBNqGuuciG1vKFYpwh0y7psgVGbEuR9vRi6mRLYSGLdW4h7sChMJBJx9y9hQRBm
d7QiLp2SA7wZGM7egUnEyZvlobReWzYM7a8IUn8KBbB3hqMFe7MQLmPenryH5cpCFgxPYrYuFq6y
b79qO58M1XEQo5+CSDg+3OBH6ickPThHHd4e9M17kDPVXzPBmLTX09vtV04YRXENbwV6mt76KTiM
fIjAQg2KaH0RYDBDcAE1ivvCdJhe2UJy3tOwQfLC0OeZx2AhTKwVv7PRv6v9g+BpN08bbZ2c8yd3
ykbT8jH0U5xfoEjduRFywnsHUNNm+2wJTTE0IvmZjdgtQsUAv4mroxOxfMmVCYDwa6wa2MZXVOsH
8FzEniYAiNDyAZgERFsRhXD1TK80iUfcgeoAXZICfeEhIbuhLXJ4XYAStGGeHjkqdV/zsBMqg0yz
cZlPfOpksjzH3PD3h06Wtu2jQDI8xMW29+DYHFykmcRHqmd6FowPD2m3csGSyieNlCR5EsnzE7OO
ETEvCWplfzIFgwlp19S3zmiwNfMd0P09Lhtnoonbpi9mle91bCifz3kCBcx3fih25BZMk3KHXtkU
kxd/gmeoYobaRCDkuzgDEnzw1VIiaF71OudJOhBNtOidMJguVRoGH77qNP3Tt5pLNQnE9Ee+w7CN
2p2nlg+uox6wpELwLOYYmxaELSZO7th6KAFMJ3bcXPf7M2WcY+zuLSk30XUb5SLegkS0CxnEXqLe
GU54ISdRU9oTGP2gHKh1PGGtfkHRk/N0bIWWwmtQY+iuE2X0HyGHrl5wiaKAsECpXJ3Z/CvM9zOX
CTyw2qAoEWuhwjJ9krR/0HFR2GnP6XQnP53bdM+HMxiWXPs2551Kc8+wCN7VfPIokBtORL6Mybtx
igHgKeY63uBN2R7Y5nqfOMcj1eZI49DLlelnPQfCUaFBc3gZIVWxDKtrxwDsQwc21AYp7ff1BS2j
eOyMAcTxNHU3wLS1PBSyIA38bldoJ4Lqi6NZx06PRV2M2+6LSVnH948406etooqMgWpaX688j4kz
Z2VV6JYAztSAe9vKuoggtXCAhGd1Virbb4ciDq6yUEHDMlEVCuF+5+xuIFEHy7QrGJhWthkm9ZNp
cXc5xszJDPgpVOZ6txA6JJHKL6dnzvD8kKmo/mX7e6K/wJGztdCIrkICWy6p1kqOJsign/hN+b2h
yuxce/p6WO2oXTxqeSja5w0XSwAihAoaqzortb7Kj3fzbzX1dihWeXBkaJMgjNDCd83w6VBYFImq
bZFym1ShJQF6nifrjKWxaOkJ8MeQxWS5PDmfKz6Gd3W2LY2uwVadrFg3c607dIIoj7N1rlfjItmb
xzW10dW0ohmGVlmFojCMAnrHNkmivFKXzReR5FJ1nVcQJqKQiu5Ge5/iHe39EIiLFSXNMWQdWXr7
mhJ+af8N2QWhNcEYFp880wsYy5LCUAOVcsxz6HpyGiy+v/wjKshUGcIWXmAI6w0Qqg5ZgDMd4rKR
46TlLK9s26ZY6VFN1ckYB9oYMbwkuUWwoJ0yltH1qXsjmLDQ3DTm0X4gaJ81Z6d1mrcB9jauR5BE
mFHXgpoqf20mE0jqC+QV5rzC0R1/+SL+sUYd8f+XUWcCWrQu1M0QPRMHLKo4Zq50ZodCIpOh0ZWQ
KVOcKS/Gc4m8OjgA7jD0Aw7gF1x+tqfo4cIVbfs0eAjO3fM2KYCiwg6RGA5GaeQxergEa6mWzNS1
+yoqn5ShxPIWHRizMVcyWLgOTzR7yvfs9mj9lvs2wN206cRS7Ofrd76EREYUVbN8yghUXEMBlfF3
f2vefLk9GvO4ikbuODR246ALmEki6FO881WjA5mq9Qt0bPkm84aggWhtBDiyeC968x1wKJPW8sME
ay4iA6Q5PpHhzHkt9bXdcYrlN1rWc/AQ8QjF7W+3Xo+03FVV2GpRpFcLMbcwLoORXAGbMgxkXeOL
fuq8Y7Mg08MAIUQHNdWOrCJBMYRoZlnbEC5/qk5zkxj2hLwRRHL7DK1ka45NwJ4rsVxsfCdLqOi9
Zg8uUdY3LELVDVdTrysNDrztfMPDDZCvQRJzvHbYUmQ2x34IvQ2S45CQE4jfp/OX8uYmtl6e5Gf5
gyzfuYUfVQ1n8h7tzxfI0Asfn4RcMM4DBB9gZF+h+TaDH2dTPLVv/eP8ifh2dRkovx0kx4DCBfqs
5GJS7nZBo3qJPh6J0sKDGyX4TjsHi9dCNVesyHY9LcJJZAr4FYH71USSFoNWHXtfa2qZf/LFP5+N
it6SAZTQeFXYSLhTxmlQmZiktUghbwaj4Auu+heMWBcnOdEy/VQJ7Gcl/do/yyEaLxKtHUBekLsp
mwA9Gdkc6tqj/fqHrrExAcvYeuoYOK/zZuF2p+bY5bxrT3wYgNT1QcWuNQ2k93QK6oP2CAD/t36T
Ovg564aOl+OHAUW2rEYMjj9lRV9kgu1B6fYebTnWLsgIPD+m2jV801PcGVI/TKFzQu9LiVPylHuK
ORv38SbyuBoEMne2wTs4c2MbYxLcSmRDuJ9Gb840zCP3YHZqjX+YhLdQUhMmyEVeDvMND7fgbv2w
hCeFuFdqTE0u8aP65HZ3msVsUr/E/oOjEIzX3aIT1r6Yd/VuehvA44JyNE4VGxKEZBS9opseJbKJ
/DJdVOiBggeNidmfHH6szhc88P3PY6n35E0eL9FzkfclmEwssD/jvc6Bt7ya5NwBtY7ypZ7PaNsI
UN319cdKu65TJ30kjfm1TMXU3lVFHUf0nURDTCz0zAe7MS92e2YxEJziEk5EVcXQu2+lLj/ko93V
lh3vnFPepAIgLwQRxzuNDYAE/emQe6XW3na3S7ZvAMXUXQQubnpl6nIEerdB4os6cscUZbeU91Ky
ouatxLDwpF19yWbNIz+QfJ4dVYlDI7LjSSJskA7Zbmu6c0LSO8/PZ3JAgzA4oJhTZU7QYNALcrwK
Wp74ZJPzbawNIJqLk1ukMvcnW3cGNhhLV5KPxatX73Zxq6k7bH+36zKzRqbHYJ9vaIGF9eqDyFwl
cIJyUAzA7ETpOhkJ52B0A+EoUw8B8PVqyB0S+mvf1PRR+Ln9mLhuBqpy5bygb4ACONjUx+m+vgfo
73JetxRrJk+SYTio7+gve9kLL7dWdJ5khgS0hSLm8qZuBxH2Aa3GKT23UAYki731hfOUJ9Bop2Ge
ppBYbsXE/HT27EnMUs/jibc6kAT1rngtJteFn7juH86XQSN0H3vExMxRbdMWEP1Jc+ksWoT7GORT
PMQ5/0dmt13d+cVfnMJOWd6w3S8SipeQcI25RG1ba/gAi2jnb3We2UpjGA8ZhNw8NApbTzYY3cpm
4ocN3lNpo5GQe0EX4LaN8SddsIgBc8nO7iBF6DfjaX5mNOsg7NkchjRZOz/JTgQrTOiFuT+2lBVp
7l/t09ZdQRNL/D81y5l2ipaRpJ70Wys/g4Lrf++HQ53uR56psbikxHBbEtsP8zp/ii6BL7zpFo4h
2J9+wszK406QDqhfu2AasQf8ngk8JVD8ARKMzerAZ/k6jVu8vNQNgMYKKfCMVrM2z+/sdvVXSxfM
0gadiCGUXiqLpBOWhzJ1+R5nrsU2eTGFF6zRXcSnhIfFDjUKm9vUlCyypykHG+o3MEXoNL8M0nvJ
NfJqelj28T3P2vpiPF3WiIOKHiXzSrpvy9yFXIeKL9Tcw5aPUUPctuN3OL9LUWDNVm7DOVT5D1mM
p1JFKM/W/o5qb9Ie6WqelSsw/L5/0KvOd9zndkLVILHEN9dpefInElidqgwFqA3OX27+/cCWLYe8
mIWEBhqs6W4QNN57rIfPRjfyhSyV+itajbZ+2qBbJ3D+ujCkQKAEGVXlhN0BstRHKzNBd7i62PiG
jU1V/5xVHbkPqexCHnoUw8wZCvU0F15ZW12jJINBZI/NuE+saDXsSG9lGp2XLQBXkKlvjf80cLhV
8P0P7IoGOc9ZwdRiQfe8eY2yvCCLScOY4Lc/c6Me6hzANZaIBtXSYlAyIV5UYAIHofcrfoM5vcIv
TRuTDkcqv++TFCFo7hKbouV/acJSYNY/RG/XK7O6H9OtQeMXNUtwcrpVsblK65FtRKCsSDnomItq
YvKf3Q5O/0RrsPyEweB4OrENJukzanVgzBSpaqvDE0gzf03r0G6EzA4YA/K9P54tvu9iAjerjOos
KhpJG3zILf7QWyDZIFizsNHLVXkOvUOqhxsvF9Fq5oP2aNcjpalCBUKINsVskD5pYXaZxc04DdW6
dBsVBwjSn8cM7Sz6yWeF90oLaTdkUOtrpV30Xl5YRKHm/y8TTq6u7gIWhH4aoFU76wd7UMR77QhD
g8mzX465V+lOLW8SAhl1GhPp8XO4VJQD+SYCtlcgAG9a6Hng/teujJwbYcmLSq32B58C4UQ7bQpn
KhK9FsPFteRRhKftONlAZZspJhdTh96M7tiEH6oqxD61G1cMP1leuDBrzU2ZaWwxXd0PRxmN3Ie/
JLa+7KOpqnoxI9xGahfrEsCJbXa8C8pwJ68gf5c9EN4PGJgsMTKulbJ7/GVCp/7GjUJTLq6l9E3b
ikDpLRdsZsjRNDz3PBRN+ufQLaorOBOXOoKxztAqCwoQhjL4j8M5BpUkOjo+ZY5bWyNx0i0bV4G5
ebtFF/x3PSVYTzTYRkO8DRM0Xu1Xp1prgtDwh9gGfD6PdjActRtgdNGKkQE5wZ/unWk+rSK/VlVf
DMrU5RTETN2m1dDC4FeRZgdvgx3zDvCwyYKUySelpss1hASCGqaWV4kXKDb/IiVb7TQhflfjJej0
aVw1rZmOxIBdmuIrbzTmZcKMTFnUgULDxqpF9h0tIiNEQhtx+pkSPqOUIHL72+unNZN2uz3T68hl
aH2EZi4FmQ/2wBCunoThJ79U5YYX/xSaL4D6bqGKPIu4ij4OZQl/N0dticAFqW99gwjA9dcStlIb
uh5q5lJgfkTpt1Ad+5qipThT5ZtAfrflEAPHtB4C+QCkQjSvRo4uqzvRESYRX8v7+8Aal8X2gRGV
lnw5syJel1zeToOcOqI3IFDaC/E1+jMVSGzVarO6jk5zapSZnFONaPbFkTS6Gz27o7RLDECG63XD
mZQqnnMVHeUXDFHiVASO4u6s9EXhreVTHR5MmilEXhaxk8Q2F60Dc5izHrN2pSS3wVZOq3uQuEh5
yP08KxoCN5JbLwOrPWueUoJixu54EkeBTrM150tMSDmmkvznMZP4Wuk25GgUOdrMP7C3Y36HqP0B
haIymahcF8dzWE4xjfSyCBxEXnnbz2K0vJhPR0UVcHH2le4JvxFdNseYp95zohxGBWY9a+g/3WT6
vzICphe3/ZwzV7phf5hJjE6QLVLRVEiZTLq5LBIjCGeiBrCypIrBKNML7+9kwVQXkN8TLkAm8Sn/
UJpOWkEdOaLYnsLjhaoHt24EBYSiUA/YmWmXtGR+CbXaHpX8ix8uOjsvOCFawcY1L3Y7NqtDQpmE
mG+YqUOUckehhk6BH5hCo6PvAABx5HsryJq70qjHx0CzrhSfzQ/jbmPBinr5hB+i271G3MbsfxvX
gh+Sa4fyxsZcSV3dGa4pCUt/clfZZWgzEj+nCBj5z7XSYeS/h6ihNbimrcBZaPBaZ2IodmWmn6fk
PFzyawTAjjGJCtAWl9pCpUG+epC7TJ73eGLdi0rJNyQd0sbx6n89bOM6CIofcAIS5xca06/y5fkh
9vcRhfcvV8D0W8C5Dx0OnxrKgGbh7SWja4Lr3MMcdPMkc2i8kI/1U9MX5ifFMP1p89vxepmRG5tQ
haxBQcEuOeR4zOts/dPJSnSAwP1Upa9ixZpcMLASBU64bpkBeB9rlI0aBOhixVZGdY0wTMUOkjpK
cuwEs9Jxn0kGBZdO9Fv8ZxVwiuh2n1wl07E0BaMuZ2bUFuix9DuHJUcR8LmHkHlnLBCRQ2flWmgI
dQ7VOrTE56S05Gt0x4/q/JMvqFIXVFbh79OAenmFm/H/fRIAJg//h/2niLWwvk5yieJnfOeWmFAg
q0i/h0P2DxcJdXSzLl79Ql2h2l+V1bJGGr2ze6WKtcufKxwNlA7B5gM38/2WaBv6XmtolCJn8KJ9
4bhV5K6pFftE2xKxWa1ns4nWs6VhBMx7wkCtnqOqAcVt0K+Q0f28Ljliigcd3Ua16CzDHinDsbf2
QSq/wNtr+v4vp4iRr3W6buyF4PwKIIEYf4Ks2oAFnvvPliVGsI3t+dUzQ1ugjewtYLtAyXIqSjea
cC/m3XokAMV77QOCCsIzK9fo6gsphj1Al8MXayqGlAGDQ2n2M31ESXTEWnBoU2u5q20FW2gwrIbj
b16ZgrUwLSbNf6k221yAUTsdOZfFe0RDOg6ABGTOnDXFvLdPa+iDzzUFQKyzZbX1eObj7gwoXDP9
6IA6lVceeKGD8D3HhUHaG1ZL46YjgIouLO6KglgGDhMIszbILaCAG+TM33Bk6ixZg8nsnTpY8wGj
8SZc+rOAvaQWJdLpbsCSgPBuKzbgCXplWNrjo1orWYmQp7bstLU/1u9F2tDDjhT2oyEHsPIpces9
/V0pqOGOmiNP7F4IGPfvgICRTxqY8ozU1ReIag2eSuDVgekvWs+F8f5u2HdeVJklwbUVnp5IWni9
KwB10xRZC4R4aWTt8nKCZSkZR8Rl35EFmefjYv7Jrx1p3UQOqYUZ3agnUi3c8XuavGaYrI1rjJcz
S7HlJzP7Ih19tQQIcbPZGaAluepaNEXBDp2HkOKAZsuHf43VtSFiXwLckkeaHGBuNtGWtY5lGYu8
1GVJEgDx1+c/e707kAlVdtErWZ1lnOxejV26K3luluwXYJUciu5TomRIs64QCIZ2O33hdtMv4eEm
4V3vPHvs7FUdXoBme4xRvPIzI780QN7gXOyQnLAl7jRErLJxSwkFtTo4p/whDiIflZLct2YwMWWo
BfppEj8JR3IuCuq6QUNBphNeaCEC052cCswYwoayrFFVfsQsrOfEnkRIb94d/u8tym38BnFg5Vjw
lu7Sbpj0yVc6lmBfWJb8AyHI4bd7vXgT1hcpClovfeaPXCWkJjT4R3TTPeuKXl6+MVozpHsQVhqz
d+ZoTf/sOnA5IwS/MHqyartnqefDpUHgJUQtO96NmXGhvb263vjWBDgEU/q7XmzVn5w1vsIxczw5
rt0+BOo+Qq5M+xGiGpsVVs3NawPJLG5myzYbtSyczSGJrd1OFCyPGGFGea50jfutZiAdnhvoy9Nu
z5o1teHOFmrG74A+2ei/SGNF1SO9Ocf6SlYCpVwsU86msLMcVUXWlwwihPM+IMz/mPcT3kYMubyc
uUwR7Zz5dM4+6bO0/Nt1yGgwfDPlMjI2VusOfmLllnEbeCDo1B+17QtGLaAQ8swXtwBnDs6LJkNU
tYdFVq3d9QZvD+WGJLHyEjJmP4oyPFrLPYxEXmc18JRhe7v0Fuz9tGsw7JuxM65vZ9v/T3KtXM9x
baYS9upsX0xAvBu1nsgXgRrjGNvb90V8YHefnkrSaW74Ce9MkSgHmf43K5e2CM2jkvut4Ddb68xc
UKNt6DzPy4hqcbdVHedeosajm1A2BXh2YjpCvDnqbGbTJknKjs6AsHxIQPl/qt/kMsQwcwmW2/RG
yQGtN6KuI951BHT9/n3T+Abt3bVZutaeYFsBpnmBg3elN6Y53gDvT1yKN2pEuKMr7BAis+CASVbT
UMX8AbN7HY7slX9VCcqrQFp0aLbAb+Lr1wGvnJUHv2A6Is5tu3vs7iCMd1tF4RoMxxgrUSVMtHil
QD2q9kUyHZgaIoT0LkNlk1Rua/6UOgXVISFAhw+tz8Q2nVuAaVb0ANrToJ/dFmMX+imFNlE5WjEG
dZRAwNKrmd5qTN5iOwqU6TywUhhMcG7rGuIjwJyKxHH9+dFeZ+iIKfTrymlFTfdxcnxATizL5O7H
J9PD2kRNFqp/WX5ytswkTxuJxRqixYKvZ0P6BMrjpBaxEol989EtsRa9LaPIu5L5j73CAs1yV6bM
Labl4FE/ohx5+VDKQZKN62TfJnIAIDpFopi/yHdMv/Gy+iu/MRD/T2Letkz/wkISurEDzKxlD8fB
fo3jdVHspReiQGf8Waz4HEtAARljrLPlU2qoBjdrxdvEuU2TiUaWFETWuasgL2bQm1NzUkPZVBw4
ZNLfNauAx+zQgTWtH2zdUgErIvGojXwmAlB466SsziWhrEcHESJUIQliVXRAnhMi08Me8YFpUwUj
P0rFXtHNTyO/YDfxJGtNl2m+qrqRlnesD24VLPSDvu44HCJYfUtUnxjvHBl4PNJJottYs4cMaDK2
PQaT51hNvlfUjh8dOwIv3pG5yoS/Toq7+JXJJ7yPGb+h/tGheqZRseW/1iYdfGiZd5Xnkuh7hIh5
Kk0OZdn80OeWRrfla1EnBl5oOMq8vpD6N/+j0h6ouw+JKwh/GMKk5atAKrr9a7M6zkEV4qh1NpYP
YOnnYPcLAXtzO/87LgsoZlDlKh8d7BsBCoCBM/oeevuCcI90dm62QfSEWu/rBWDH9B8SwN/FTVya
B7yfsvF0CZDQ5MQ0goWxF7jRqqSRQZjrrXURsSE7zpyAAYSZDXbBFv9ddJOFHzeABu3vzFpulbae
sgFDKbu8hV6rhiTGCU2ZfqsDuYpOlPRCujyvMAiiM9zf08lFth78Qrlnh7rfmBjDCkJQMTJtmyj+
KY1VccvVwf6wb+QQuJ9YQDb9iPSma2bQMXI5jXeITVj1HNESLu3MDxYPtqRCugqO0qB4bUAvUClZ
FXSIpZXHscteiCFmLFgRSiJUjgkAeDfU3J+e/0SikqojUSOnXUZ66QhyjfwiGwHhOmU+9SDB0tox
xqumE83JwM0bcvQUezlG2Xmuzc7MDWXbSq/RksLHkx9ehlD8v+z8MkZEOk0olZeyLWH83ObdbhwH
HZQUADm6KDmqiNvsd9Gdm6sl8FZSPAR9SHTs3Kx8gMTHbyOa/FU+wpf82J9M3+8kyAXQAqLxQLDI
oOx0e6fahUSoga4oV1+SPWma8s/1j/xtKkMaD5uW0eyQABgJ3Mq4xcLmXBsTI0DEd2tP41RLnHDs
KVmEes3Ea42K//uw00QdksVrdBihdwFmMFsrootcRkcOyB5rTJa++IeAlh7Qkc8sRtXYKlZzdzHD
ZUMhlPIHNiyRGJ2LObEWFa+zIlgt3bGyd3l8zyEolZdCKZkAy5PcpzQWaCZ4/J16tmsqkrjQsiTt
Y2PmYTJQKJuqx0cijC4dxdzldpg/wHEoH1PXqjsudAPneBqq6Max4Ur563bXTWA4UCP3BPfRtw7a
ChiX5oIOsFTWgMi0dOub18aW9cGaV+8FYZRllli9wFzozTbCBa9jCgCl67CuyYw+6zEw3HCWr9Gt
v6j7pB4jwabVGhSR0M6SG+vQ/jyJKG846HpqNRLchdA95zFIk7LDC9A+SjG2uEWoo1+2dfiiEpWw
o3TmBXiBW4VOumKXs4fiCpMOmH5Q8OFE4+FE7jIt/GTY6p14PPz1TXLsYi7zDz5lfInH30WFYE/n
8soRsGMAPXdrSx3585W5YoSs8+FH45fOLKPsD8nXeUvdYcGE8c3NrZT5gHJTDmVH+2INN5jLto36
R/tfmP0LTfZPKaCgteX02WJHmJnBI7AtS89w4nC2TGHxCHqMdEeyPHbgrv1OTyL9h18VHlwVtXUH
DtigFo4PkZp2ZDyJHOkTVWZjehe1jDkD5FTeVzmX9+8nnn+BO6Y4V8pFfW7QdruqkNq/7CLs0yt9
mqWi4/FUz2+tCqNweaOP+iXHJD9OyaGUQ27mgbyIS80K7ZsMoGKT0pc14TEP+LIqgblshKeOeIWd
ekxwpqGj4sDgfIxkWZjcBUbOzsjZHMQqtI2dM22m8ZATPv19Gp3dZ/oqvajOfwaXx2qogiPTWMgz
TPsJN3si49zUwgpKM6jQjUga4METIn5kIR1EQetgpGdH1ogQYaN/U469RXwOG+er7MixlWQvqNN0
+3razYheCCaHtzit+dikdSYltu06uJ1BGLIEq29k/HcJ4rnvqw5Wh7cF0ZB6nhZFfYDcT9QSvPJ+
VgcxnI/2UsW5hQlTFiP8cTdcP+9V8WKKgFSd46Uhmk+LHCLbMSy01ZL3h54dZFf8ZC+QbPbxPGqr
6aOgK6E1f3CTkjqjzFBOA51XlR1Q9T/n34VxzGspJeiw5fsHr63UhB+/jeUoW1K6XiDyuEM/LQCi
SUZzROirRYk+n1krZARfO3RlnnJdbXF8SVKSiObgNWO50RjCyKSOlnaUGTz88e3HNfMVn48ZUB7A
Yml6C7PQ772kYQf9s1KFK6zy0eoicCGkzI0sBYxx5DFAip/e4lSgAWzKZlkhiP8B3Vs7oL7xHgxs
BvPWInFwBRV9JhcZhv33kYVC1OuOmVaBpPjHlUwjm8lMPo1QMI7N/vFpUqGkbtxkPg+G2rbsjD2H
ZJ2YG1H8q16OkPFyWqVBDEyw1q3uYb3rAhwdANTE1TSQe4XlYft6vlnNEhi9gj2wLw8VktVv98In
+3apQLKz+nY2aqg2jypOHkF9N4bNtffFjIJJplTASACKxTyMS2Aml6/XvLv29ValgWn6Al4Cop65
XlD35P++xzXNFKidx/apA53r3DfGEns6qHRLEFQb4tY+ukXzuzmEekA9+lxTKh0wOBn+SKGonkAF
SCmMUuKOo2wwO8BbUex4EVZ7TmG6Edr1Vlxlcoc3SLlYcvOI2kze156/5JX54hP6X0fF2B3oleDC
T51lxoK6IvbCoHOiysoxOreK9fkbG78Yth16dFNE1mM/QCAqHfJC1A2hyfC3QXPz1mWPLpXdFCH5
YcFBgFmU4tN1Qrtp5swEo8LFUPHnTIR8Nnwu4zIvGI1yHUvRR8W7Apg0NK5j2OQS8szaoGF0z6Xz
zlN1aAXcNhhCpvtiIb+lbWjVgUfPizo4eZ8Ia0fCH5aNEYj6K+7aXTwjsXKQawFoGb4l6PZalPLs
+tyc6q9MI6WULuKbkJqjgWgurS5oxjUyktzQm8z7QWQ7K1aHUmGH7PTlDO3r85jthYUv7lPGpAGH
LhK9426yoKSs9j7G60TlAKWmNmsR/b61DWMk/og47jailX26ty+0P6seqr/QCJZALjIHid15fy/g
xqtP+eqQ86l5QVmWoFX6jtX8thgGFjk6TeUuFIbL8o4xjg++j7ianu8gDgYStkrXRYgAklTH6ntH
gUqvqzwDoppbDlNuzltNrnhiNjX1ExVqFJ615AxmImLfUASuMocXGl029q+sJVYtIgw244srXO/R
LvccAMbbxtUsAp/ftXvLOw7PUih4b2thr2qugI7FF0965Uy6UjZrsHMTNYBc55QwBRqScOrf1xyZ
xh1K1/z9pNZqRsCbjfagDF0xDD3ldK9cSmk4V4TTKpHwgei3OrdWKm9RFPEUxrlW5pv5/BV9jPig
8Sy5/wZ49OdlD3RnkBV1YIKN5vQXow6zEFK18bVXS6OuC+2muzoNi64huIVS5uaRefL+KtAOsNis
R6oQMxiei1emtGzX+jf1QXbvYZGa79En8CcOg/GC+jeVyczcpBwuyNMU55uH7mHP2uRxe1pKVYmR
fYm+TCTvdIGzTOVXrsGq1vlJuSyWhtCikNgdGNUnuQhV8ZxbGCPeZocKxHhCa05RS5MX0AWgHWtt
lMfKUhd3omO3KTatjP6o9B5AI+TEbfFIVNK6G4zNX5L5ZjFPkOjQMrGMKCXhn6Jqczxe9FJv6pSQ
wvz9dSBzSmWzI3ogMBSFW1yvdDoL52r7JQs14R2oBjOgSIvJHDOmTciniCoFj9Za+CbeH0WZvD7s
ThAT16Dv9OsiKF5GjshVs7O3pXn3sJJh1XvSzEHaceZX42y4fSkXwb4YgpLFTj6/Mv71iPgUhJuv
vMsi3TPZQeGLbpCcuUVxchI9VcGPOeCxFlJlykJIH4f562Fq6Z5rL+DHWVLwl0SKC7JP4ZzaWovK
VXzdpidmHPpUvWIfxPpi0/kx+TaTa7hLmOPMjE6AfBl5xdU/o2nFg+9THbVJEmroTd2EQb1inqMs
p2DlUFc71u4MOOUXFyUsg9+uW5YkjpNUjn6HXioxOIHFXbJxfnI2lf9zld5+qbaNEAGm8dw6qhff
L5H1rXmXB8wGxzkEdHLlcRorTG14W36f0RtkuJeaPpQB0UxpYLPSGAv0XMMxnQ0JEpJ0xAgYNa6Y
ocCpIZt+yio3wy5Bmvt0iCF6SZBW4GSOxng6sejPJks7DqYOK0YzCPnOT+hxP4GVtplenMip7oY6
4NVC9zbcG9GMDcEVqqAQI3ofK6w7YGFvTVl8O2luLY8hxcwo03hiLTr9QHZIQzojGUWznHat/aJl
8edT8gnkINKOIZ/ELMpSOJjfk0LAnR9Na/aO8Gl+r7XEU50LzQDb3QaxoKIDgbKZKnPS3hnH9aNd
J02ZaiB9UPTd9YdCzmLCP67tAXFuznicoKP5Wdpa1zmUAOJMmpJCUmQKACD8AHk2LPhDPHb8cxGF
vx1ZuaRAHRnykn3RsMB6udGmkY+ZOtPnJK1msaKPqxVD4cQvKOFH1Zs0MGbmFGeHq3muJzUvHwvb
qYK/4m8tPkQWYfF5BIJaRIexPuYvBZ3Hbq+/PDm7q3bjaF0+Biogh5LLZ6LiGqNhqc9SjnTM8bbi
4wLjiJqjJ+Kkyd5x6PxSf463eRBrQCc79kxevmVB5Xz+i0mQLqu6AqJ1KzY9K+dglaSApV/JR7Ov
c6iutJyYYRTAbB+5xbRt7vdi1iZXMVZRc9H4NQgFBTDVdrYIN2nF6qepwSiecUZiRl8lyBhB43fz
V6YE4c3e15Y2VMPmJck2Rnusp5JcAuyj9Mng7sOe9Yr9iSbSvUHhEpFE7qoul/kIBbe0XaqKuxvG
GCbR/s1shXtoJjw9j8egls+16BsCNQ9PQOxPcuf+ySnAzatqsg5JSge5rK8Do5kktWwX9v2A18R0
lYe3zriQRFvTHGPIXsHS6wdsltA7rugJgY/KUnEWJs4T0DIvETsC888aIODld8YhBUvIM+NKTumE
72Ojsn8Dsse1sY2OHX+vRiCZjX21U5drWLd+cr9/UXuJ5JATt7O8m6tUDL4swVrX++KD3vksfVAP
crVy5EkgVncdSqY5AeE538E9H+YCrg3l3A0DZgDVwUAW+7guSDbFmgOSw+2S5yh93WH6vWopRkY2
zwM26+Eu1W1PyEqbVJ55epGUcvJTIDP+nIKu6dRmfc5Ea61Z9pabXwYj7SsjWE8r+ZV2F3/y+o+v
NXYA2+R5kyu9IreGYutPMihK0SFZZ5DIBvLzgPXmkXtBfYNp5RONa/095Ixyo9479svB5AO7jrDB
wTa+xf8bCmuvBg9J5hG+0nmLQDFUPLOt7stJ0sGEa1Mf03t20QuwEMxqAEOjtwVCxOz+m+gb64hG
Anh0Co8keM2Sa4T8jv8zjB+CH9O/Kxz7tswo2HU34KVxoxBc366pReJ+rkS3m6kIUs9BjUAuP5sY
Ot38uTrcAJHcE6AU93hcY39NOJc222HHwx8Fe7m9NFu7o7NS3q+BzCFvHpSben5fvuZrEvg77mXn
yzTL+HPAlcB9CkE9tMAmMOKUQywaynOdCrIXs8Mum7NFHN4z7oJSRvb93dyPrxdQQs4mG6QvJtZo
VoQ2vwnNvXQDfuUOv8qrBBc6Boxq1fd7un7GyxC6m7rozrbW8HE41lGw5qy1NpE4IRazA1/q2k3C
YYUMrhnABZA5rNgk0fCpEu2kFq1eipd084gIyMMHfhfuY5vAYDlWEn6WQssO2BnNcV6RHUHMumna
fN9ijg3YK3qIbPs6gDe86PI8wVJZViXm+cG0BJqaQrHt4IRb7+7XZk5bJYgNXQt+EkfM73xxHlvW
TGiOo489UNhBgEMccGvx/FHRE26YgMyY36KNqlGAxOi1NJWiaClyufcP9+MPrzm/uU7knIoZSbPb
+wXg82ILB7vA/yXIXoVTRzkGmam4PJzG5Ki+Ve8skTULVIPV1nQedlDSUbZ/GyV/fG6n60g32kY5
QkNrNGG8k8Xxb55TVbVHntYytSk89iT75T7mUoMJF5opG55rsnueRTw8fv7dtzSsqdFx+I1Ip2tw
sCzODbKbggqTG8E5+aRedpMFj7bTcoMLwROs11myhatROz1lCAgcJLUyc0mZ6jbglpf5zl0+F/+F
Ft3lJlt606rO9PmnWWSkaramKL8Kdz32EYWvtFqtmQ/6QEhvxJhaz3MNQaIjBI1LopSLz2nv3Dhl
z6Qg+T6mc/TYhH8M3BNmMGEevflmVcupioM+aw2nj40q/1XEernEB7vFHbPFFQyOSA4e9VJflEdc
oHiNvIA3qPRRi/e1kFleYWwxSmmp4VBxTwG9ydJsL61GCTNhMKZIdvPnQmAr4chUS9n3xlC8nHGU
p87CbzAKp4kbtG8crqOFGaxOO4IPZyM4iuYjFaIZUqILHcxvoJf/2+FTBcDqIyzDyCMszs2bbT0h
VyD30Q/VJpCbGFGOGNBYGC5N3QKI2GHu2o5jndGbPm5JEaYEguzJw22qBy5Er3GQSegxsNfvSbqm
pAr+3NFYWRYuszYkT3onZWDeUFxP4KAYw1ezoU7tNXRxOVsyFyTVDZCd2nbjdzoWLUipFCL3TynR
Uv0QvgtQudLl/bt583HWp+4GbkSdt+2Ronpmb9MjwcWai/CKIj5BcvTFzoFbLX2XXZm0aOn2kYyE
xHuI75ZKlxto8qVk0UyzPKjA2f3w98o52MO4WdnMfMiL7/fsEYa2H2OL2DS/Qcy1U9iiyfcWAYFm
CthX5eOLndV8W7zs1+EfshAANtPaWDF9twI9lp9DaggVu5CZ6ksBj/x5s20xZOdT61RyFXDJcyDm
NwGJSlcv6xqH2+nJxlrjHMdgVwvH4ouJclA6PwaKKpOV8XNJ8hSJoGz45hZy7W07ecBJt86sPDWO
RJKv1yzyNPJUa3cy/c0i7ZA3j9lTTK88v93qRq9wJ2OrFEPpfx7MX9thwGcLiznGfE7rCmMlHYUB
KSIL1kTPeFvcrnQC1N1rKnnJAPRaxpKDXNi194Zx5sRdvH2JSbxBepm/K9OMJM4MW5YgYDqhLGeE
/ha2Z61EIXyIrebI0+K7eebACuKout7zyQSsl6QfOikPJ1uKdYkGu0cXkuehMkoAwgbXMDuo4/5W
T7TTXJR9rRomZTcYSu2zsPnG+iyvpJY9ilr4L284aGRmoO+MLATJbX0zwnyH8KZQzNgDdIUhLK3K
aOgiyLle4FJf7TqK4dcfBkDLX1NlQ9g/HFDLNRRc2ww1ZPjswxmGV38FZ5b6dvkHzVskKzN8Mdt3
wInSrX0g/n3uj9kV8VxWOXSu4bOBGoKmXDRkr6BZjaNlsnXdwRXXHkBTDBssq5l97sqRoepXJlzx
qTl75X2TcIeN5gM8y9qR3VQXNQwrDZx+WiCuKZf44G1rfYhKtvXvoBIykmk64BWL3DyLI/Mlp0B6
++B8Udg16ijgYMYmJDPsYOU81CuE87QQA1WeeXIoEMCbb9GbVvkx3ISOtoWtPf1/cXb3572StU6t
FK6lZUgSYFM++cVOkrj2KobgDYOv3P1kGNB6V4/c1vS/vIb9hkWTvmrWmP4b2CIgYS3JM+dub0Jm
Z2Fgs2tSYO6S/w+IFoE9nvhZ5Rn5pVft284S34rFIGjFEQetShb5rp7r7gvHgJJxjqRSd4tXVqbr
0nP75H4p1XI/oHFNPmQPezELBbIDYYp/HLvgE7zVksbe4byWTv4Hu4qWPbw98W16riKG65zfUcG7
XgO3f7SuV5JpwKP9z3v7Oc8DLJc3SsK09xRgnVBjvVW0hsHJdxNXE9kfYFNz57XLBWumINAjpxLj
EHa1SrIyhMTabVsms6h7oPgJ0jGcO8PXyQNrclJ/MDgt2mw5OiNH2SIDHhGAz4oQeP5iZZ+G16ba
NryHhhEXe3ItLy+RMdWrMtkkV5Dbs5D7/FdRMxpnelHguBTQyZ3s8cd0glQAH4F8+GGzm+fX4Cw3
J80o6svzZ9u8prVnrNSlS/b1TVNkDl/MqfA35hP2ApVpP/XVFle/vNauOeRyO/RwpGbZZKqbgntd
FifJUWlJJRe/4Y6YwET5u8nBVYkxagrPor+OahIYXhTapdy74LkPZu1Zdu/h7TGm2Pb2TTSbsCrc
r2Hhp224wh4xDsaptJn+XsrAx5diNqIOhnBiSkK0fGPG5bDCvezKwZ/b+Kc4lr37elsweNTiDIiq
ETiIMnMHiomES67+ANAWR/6NZfjUxQqSNDrvaLOLLN1BQKUZsC8Xr/s/N6YZxUmzgnEdbVDwLu1J
Js/BsdIavBHalb3SjoAL+QmPYr93Yvcwx9zP6pwZ5ZVE9cs6fPYUdpTunNU8pYJERfQJZAtLSWOm
NiV2iXorVK/VoYzz+0oOP3PvmZ051PnP7rIBEiYMHatD4bVF7qxbB65lE3LelJLFUDgJA7/khvpx
qCYuQDUpC3fsTHF80l+19QVzocqqRPNU8KZPDKy5Xitt+Z3Yf+0BGkHUmkyczYHz3jQK4mya7m/p
elUp7gnmtriafFITbl/TAaBN3gKIyaDoROwDU9tIzVmEHjPKZ52XOSQXmxGdp2ZikWfywZR2YLr1
DNziwKPOAuXe42Ot4mB+f49Z3iYXapdxcB4HoELkq/v5zhpW/7EdhxQxRk8K2sItXHduc7PXMZw9
5QOYTcI35cSk7hCVXo5XRoclRSOpLsjKk8fPO6IyIeh5PUoVMhaXuMXzE6xiVMOPwCYgWeYgiACn
WYKsUdi4vRi22qG9B1JMX3/68BjLtfAe+TCO8aPr1N8VaN9d1zbCyisKBKXx3TmyoGv7Dj3/pOnW
+sCU6ojIbUnp5igrea7RivGxKHp4blMTZjNSGx1yHWwChrk15pOOtuUJPHW9SWz442neHs8xdYSN
XOcWwHg9QUCd+BDvtTmVA0IBbP4M7f2M2wNy7l0NX43dDZGqU04PyqKETB76n/Xbfw6VWkkDvgSa
t4SvFB+4k0VzFteGsHlVnp3nsM35oFzyfhn0djzWLqRl2/6rblKZJXgcb/hMqVJPvlooM4e5A4NI
q8cBres6Jr0FG6wKgukDAM/w+ZrjortDh5UNhmWudPBqPiujUPLQN3BTwubW7NmwYFrjZ98RVAZU
9c5B/m3HZFt42Qe9voGZi1ogbc5s1HvFc0Td2X9WrE7efOI5XnNM4tFEItCBbDHJ9DQkP9tBM/Vd
YHUbzmtl4XbxZZqKHB9AgIB/86uCXhwqMhHiefis2vmC9WlkRrslV6Zg5R+XyDqshXc66lIYJ/Iu
awE83aRB8MNXAo5HMYdptfty5bbp/zct6B7hGLnx1epK0w+E8Gj4NcquXKVl4qfzvGOED2t1hpjH
E50a5bGzLPlTi1SgKZSTXQYBgWXHFAoFdOvsN/njqMTpxgETZLQVjR3rrGx5oMa4xvgAqKs7ewTG
hkizeK7ZIWyg6iFy34JRQkKEFDioM5SKWTwDxq5N1oEVQNS3GMbX53tDfjHLPP50JsqMCGEgmahr
lTEVE+0wd98Z2+tvYbELEbdyPbolOqkWagKCYd0c/1ded6FRvh1/kqezZTBvfqLZcKqu2m/8773V
6B3eV708oaC8Kfs5q9/A6IOQ5VoCoJePVFtIu8fSClAzafcWdML8oLJqhNty5yh/Qln6kcrb/X3n
r0kTm5ENpkO93godg45sXGnoQwn/6xWyAIio1nMjcAA3aRif0YQBf3dh259S5Bl0JLAGyBGhz/64
XwN2pq7IRLbtQdUSMnUfJFmz0zsN+HLCJBOIUxoFIKFF5Vi7DUtpyViF6TIV7j42zOObhyyayHlP
wFVUyKNSiMkU+IPtiz03PJUtg6Bfnqg2WwlhgdrHI3GUqnx/YwjZvrW/+z0EH7QEqv/9mA8IsXKC
s57whssBjLgBcPR49QxYlyf1exdXFOcgh9gQzKjZ/lNgnpDcxgueldkI4Qs1RQvlSnPOcEs2ZK85
veaymHVppzjeG9QSFZ5opbPBbuvcZmfOtZ6x7j5+9aDdgBC5K5Yly4r118fcsqjUvcUR584dHVF4
6eyv0jn35N61w37ruOpiW2sZ/zUEYgETAmm6UCY9uT9UfZcqsReMgh6kolnnLXPnXQ7lzSQrOfJI
np8/q2ixKa1zl7XiGxZc2lG98SVIm0N9/6AgkFgnU+cxnp0c9BCzGV1XseynZ7PsBYjNPYaqK/Ae
ASo3GYGAxvlMeib8bQe00+yFMofzz70XBHEmRgnONGDBDxcqTaZZ6RjpTCCdJKVXU5mP9NlCHhTa
sxTZYNGDS8xu1V45VIDFvtgaGwrvN1fnRQ+1DvmG/m3+4iIieqaImAzaNexoM0HP1teA94FVv4YF
Bmb76IiJvnL7BtamkQLflZBhZ16md30LFfdbID29HNfFtdD4s32IiNYxxyojaBoRgFhXkv93U76u
LgNuk5rQNieTJmZ3+s5NcV6H5Qcx+kJq53/M+4PJf2IyY2gm80JZOYXfHtfqCYOVh/94zA0EDVfJ
OIhM68/EbV97IpFSVUqCXJs0813hSJgi0A7qfnyQQ6/PCslmAXe7JQJhVz4b/7q9nbUZDDLeGpf5
/te9TiXNDnTrIVmVxUcE2BjkXv/DaWxNMbRRG5C2rJ2IG2GLuROmVy5gbprt2K3x0FvJWh3e3pMU
Q4Su1gM25Y+myfPpMGjTzY3UgQyN8LVL7E/BEdss/Rz93AJyF2bnSBJL71EQsPczTQAmjGZIXt1r
CoR+lNjhXj5qyWKUmB79q4Vt/MGM+CopI+9/PSMZO0c65kWPf7gQlUV0HCxf2il1t0rz8OWOZR5q
6H5uhg1/6SwQ1loBdNJ53Casvo6BxS4ODYw6CmDGzpaqVNxkoJlrabBdGxhYDS5vWIlNfTC65/tQ
irga+T0ZBpLDF0rbv8dLkqFSI6ufCYFx8cL02HrWRGJmgREK0dmSA6E5BGCZngTDuL/DdixsrITt
tA3o7fg+VftAlNjyIx0wOiy4C5ZuuATYb6SPSWuyBMYoDTH8qXj1UjPicu+t19rMs0/exFz5dQOF
oJzlG48Ssv8DpJvDFIwpXQClzC+k2IeOxRz5t30js9df0eN4zwgySrscLb5ycYSkTqX3jhRkW51a
XLbkZGhtUnspF2XU36Yjgz+43bESmMzx7qufgt8BwBWsM87z2uviftVmCR9G0v4/EZfjPOKxjuPe
Ivd9cbtPv+lofRRdc8bHY+SITz/h/CazCui7U93aXL5+rzCXt7wzoJLNw/zLHtV3dNzRd+UW7tri
+MuLC02Gm27YWXtwWf3UDkX5OjVZUGiOSR/hkSqukYfubnCzCMk/JlCevs1pWF1QgrCiSBfhwy9a
pJBPJrRkna4fkoLc8j0iAGlRLXi/K50R0V/WmTy97FDrhUDc2i+b3iyeFx+Iofn6LIAg2lJiBUR7
8Kf3kcByMHynLINRt3F7MtwGuwT4ZfdSHwV1SwsHacuaIX6i/YLQMvmkO6mkNulOA31b4hFS1tAG
ZgseOeIj5U1TxvOsB8dkblDEcpYvvc/BQUKdjcL17lo6xw0zMTyvMnpNxyXoCDTTj9UrTOxOnq2W
bcFT+7Wazq8DTNeliv8riqkLytS/0SmO4U3JTOQ8cx0p1bFT8yBD7ruG+wIduFoQqzWwZMHYNcLg
usKZP69s5t8n0T/ReobWNIpstFwHp7cLO0IAvSz7qDgTUiyjrnfhs1J+i6ifc5a4vmdnXdz8JZkD
5HCJLIm+VcUOX2zBvbeCt6tCHm1997rqKDNelAza2atqAd7AI9PCl7obqX52XfAn69SF6m5BmpPw
3i2KFpxbhEfmWUH0QnMP8P9zsYie6lBLqx7aT06FTkvstxEcU7LFOBPn4OkGzSEYgXC2mrlv9wg3
bdaty1jTKu885ERFMtvk1KdipMpCGuy7OAGhs74JU9Ljm/8GpU8FIdKhZxpT3Hc6RrKJYmUbIUFp
cZBqTbX3NKtMOzr5K0807GkbOBEHixehHFQ3TWW+o4jZjDK8CjiyJVrdC5VBq4rTaJDO1lzubVbB
V7dqhd1CcQbC/ScEgWmEKULF3GfUlZsxuxIcTy/ck5UerTEI8kuVLJl8wqOnOa9G0nV6dwn8ZxPI
ufMJLI+mDr3+WyFQtc9QtRsg8SQXngxfymxp5xAoVblHGLZbwNoEM1RFIXSNHrAzxrOzDxPfL3Yp
Mws1mO7XVZTUi0xkfaMopBXLHvOTvXUW+E4I44j8sJW1gZyIJs/cpk/JILQGizz3PpaPTr4NNIH2
XZq7/YJDGjPKIcW7+O7DVO0bf//P9+t4ZajmcnjcPIwwVVn88HNaKUm4asVPKfPN2PkXxxfusfVK
A8cAOBsFmWdhh3xfe7Njw6qWSdLFwDvE1C9TnUAx+X0o1aI7PP9YmfEPDtXqKBZJDaLr77uywOq4
noRB4sSlASV6r2+t+coBywCEcMwzY+tJCF6Lqshw0YmUO+NBJ6HTD+0SZYJtTO3wsmROS2xQyuyv
BHHlpMXIKBALuNPRJ+VZ03o7LAsqNundqxSfQhiF4QaaYO8GXM5IP7y8EURXGfKj8S9Q2MYt/5kp
gdGCWLpRYVtp/A6TcymhF7/iyhX0wqZLGjuqFiSyxO9w7Ourb57D3Jv2mi/JqHBPMnSvCgiDMMi+
TavOk63OWS1hHF6/0n5tpHmlbuGkIkU/2Kq0dt83u2M2rRRx/7dP7L1FMSpgaxrfri6JB0Cghd5y
UjhSgDNu+r250mLKyXOmXqFAe5q7NKBfMaKzy4hdMvuVW6RT2/bzHYPTgwFQR1llryTyJP9/XzFb
exKpRF09qN0f5UsoBt7P6fQ2Y/a/pLuGZvHLIItWJTk0kBZtyVSiRbprHc5yvjSy2g1GclsNp39q
z1wYmEKewvq0zKcKWjnhiNhRX3ieQih+JQqC9XW0J/n8nsjH/iAifpqxIs4wD6weOJoNW/iEj77i
ihCajdyv8Np9EFsXvGbyFfF3wXHHYHm4+EwGs4ftQ/xV9Mp5wH4Ai8xegLtZn3mUA6hN0QBIV5dJ
tugCzTjX9AkAXrMwfBl9EV0r9mCTMaVS+qxa87/oXSid6FFhTkYFIZk3SZHMfImc6zyP6NEUY/77
pa52VbytVggDBfuWwHmJeXrC/G3/W36h9WkyBni0LoTCQhdcoQasnlyoiJP1C2UIL20U5Blhz1Yp
6KDHpi9pYrkmsN5HA9IfVN+7ZY6AO0KqoGmjzY+aOn0IrueCc1viIit6QUYoOTP+q3m2jAeoaKPQ
5HRWqmYOiY6H8jxKX8ogAoKSfSmmBVdPFLjerHDoR18IKjm6vRUveGn0vTo3hFCcbht0DFE0wHhy
ie7jDnBG0gTRc4AJmq9ZWkGqyfRGZ0iCVc1VfyenAB72LnKfondlw7zG8Hes3hmk8KvrcEozCtTk
f8K3FfGFIV3OZwtnWvs9+Cu/BMaa7aTbqsqXptOx59TMXHxr1+ywxGBrC3Cde1kfu43qJBYeBwNy
TVH6k1+Byu+WClTwBpNLtGNxIsaRQQReCMj5GbdkNAOQuoVbPZIlr87yhyvPffrVd5QGYyJuSKd8
FDbfVvvs9rJDeEBWm+0uclwwn+Bt1jQeX6jzL5e16UlxwaryMkCG90/swLdfgdXG83v7fOpemXsJ
VhaD4PyzFoZFSVa6dLQ7h1fb6ptT9z+rRALk6GGavpXZL9mDQHiVgXZb23W4gqUO2+GbON29NC12
JLV5i0Q7t3ECQFHrajTCRLB2rS5Ehk/LDcKawCrrV7F5F2l3fy9PXjcQrBMtsFS4CM0W71hpfCyh
iXj2kRcrVIE95zKyK7AyJQikxVuxqJr5PAfLZCU5w+o5NWxhIv/csjSnPc8gL22N5Mgl5YlUUK92
vbuHTZoFkE7iGMAyLI39XQwTpvq18aPoSIadFn9YEzmK5/fj98bojx41RlyeJp5PmkEW6/1Arqzb
j7pMIiTAOHIOd+q7lN6XdOo2LgIxLeYZIOQ0myh4axOKsaHj9chTWG16tqwfI86sLU1J5CL2fqK9
aUXzPymu8GFSe+OI3ucCp5pfhU8QT6HF0ru+E5ZfQXBLOA0QGz4eUWIEndekXCA+DeO7cVuQtwIo
0It3F/ka/qhL6sPQ2zyfUVJ8MA675U0hV+AFqXeUcUw8wMrQG++Fgtjp4eoUYyUewg11H872x5u1
/MnXctwGLhC9DPXcAlID/ANGI7+g2w8pwLr2udznCmPIkZQ7BmX9MjzAqItlNlMX+E7gsOfvhuPb
3VMlE41VXSY68M6vXameE4ZnFKbxymImrqNfEKlgThi/fSoWloTBiahwa4tXe3zG36AYKedjyUyv
5A+mobMR2ETyfvdW8ZyCftfqtzjqdS/ZbHa1Ihho6lb/ESjVcAcwQw9udbJhqWgfqDdQP0wWPdMU
jhIqQKwgN6oh+kGVAmJp6C8xXjMN9wAAULjGwmwc2byzCGaZJRllpoWF90UsOBUY7Csern5A8CCe
W4bAqLk4IMOoZhuSAUrrzivykHIrJtxhnWy+I/ecv31U1rKsJnGHD2QJMP6P3AfBIGQQoExIosRj
8RIFG0BRHT50jESBHSC91FdSY1+heyg/7zwVpoohftMEtYtouFAiGWFm0fUAqgwwXB98YbMF/BGx
+S6Cs3mI3tQfpCNGFUaZY3sJPT11ZB5rwAg5harym/alyovtukMUU0P6ihh2+bTX3Kn7++ATM39Z
53eE1EQpN24j03JcIeOoT+UjRXfv+nYBcJA5bQS9jwDdZv1c3aGsQCokdviU1vIyLHMVZDRYwO1B
9boIJmgGfJfm0ReXQgOxPv1kPjigKSLO6VNqkcIf0jk/X6jAtINGm3k0DpIOH0KaDHSELzwNHeoP
OUtGlikb6y1f9Q2/rshjec+nayb5oHGgNwnE6tuLWCkpCtfZORRMlMOoH6kqQArPOsN1qzPCJ7eT
1uEwzx3XqPf77caa62UlL8gmeRJoM7cJkoa6bIfroSe1zYofoMJ3A6JtQ3yPP/gYrhNd8MIGDdgH
YVm9/aCBZfgsUv79Oy3pdD1k+zQWLjnyRTSkTE/Kql2qJWzKXdFAku+oLLWJQdR8hI0xt/7x0QbD
oZszzfo5bmfyMPAYQhp/AjV7hTpcHHglnnowJlhquH3r2BlJIkLRkL86VGQdc5+MAWxuEzDWXi40
5v23U0FFcBEQnU9ziqLsBf/zWOO94dCdeykgCFV96Vu6vmdLCZgm41suFatPkhZwrXYUoIKIAYUa
Jnz38y8h2bxsp8MP5HEXhmrkg0SCMu0nsBkK7n2Cq2BAl4Lcn5xaWiwhqmToKuLg0ZhM5l3yG+PL
teVMy/S4bzhTIuvz4Z0Dmn7OD8NJqYF2usux+5+HoeAwsJs+k8P7BnUgDHoI5E/ro26nHc/ELBZR
cpeT0hrED+F2VIwp2ycBKjMAV9pThkVel9Z2C26U7UncAg4Zz+wsD6pMns8wxlp8VbJrxYSkU/y0
TRrhfSdptm52HGjgUGZpmsUfz0SWBMl3pTt4l3ntip4ju0SysV/gREjOzG5CpgcvI3ZxftFuvw/c
d7i+msvWt22xcYcjKD6juGOPvRb6y7WdvsWLRFLjGaviRPsWH9A9CtDxvEEof7/DfS3DZQjB8zKr
wIdccL2+L+HUVNrxnc9OkWd9XwB5hN9Q8jJECIjyRTcaLsjkx6i2jYy0VFlsd8/YWh/cXOMZyDzC
a3xhyHYWdkZaS2HGq5tdVmE+7ryy6GbEE0G9nkdRRN1cV6ZiaPMSa6f5s1od1hvwAlgddsdACjz/
vo0EIxqgN7j4TyaajXqeVel7hqFHkrl2IfQaLC35cW5pbtbskVGRIRo9DpjYeFN4NREmGQwuzs6F
A69UbyU9FixrB6SEM88iUa1UiAq0vJ/wO1nq8TlY/bU5v/6nndDItLXwf20t6dOkp9HcZ8ZkBlxK
khUPcMTBBcUoibW0S0XJUJIHtY9GE0MeVFWbuKH1VScxm6Fu5WjQfezIYgrrVf1aOzRbfTPKUwA4
qgWq/nc9+XLRh7X8yoWFZYLgh4i+VY/TDx/OjN8ID0WaPFUFbe8hkbPThrArT08aXQFIQzwdFyRL
atyCmk/EnG6ktN0xdP6aN8rqN7ZhOBJLvCMeOW7hZDzAZnsLCi+C4/peh+OtwpMku3dVTx+TJFG3
bfwdXDbzg0o9W/v9DnEnu8u7JWKTWnEwYt21B2DlZ5qFJiGNgizm2pfCod0cS1embjzfIyY1jIoI
KkRZ3240EUiUuN2a5x+Do+qZSPGApbxeGooao1IOC0g5M+5Qnsbi1NgVvz7LNXAYVIv5br+SwgG0
LJDPyOia/z0vLJa2BaAXhBARQpgonDYrLVW+NKMELH41nE/zyOSfhP2MofTwAarSKfkH6YqpIzz5
U4grWppJJt8kWwlRMTHYlQby/1pyfrzzwKvKDE35KAwFOsSuVwcb+8hZgcHiR5MiThSQ0//uRp84
jjHtI/eIcvVtDZ7cFNGpTm7EAf+kvvYy2GVI08+Dw0HVtlNtScyet8vyjin6CxsVevwMzO8hXAmQ
SmOwXUsfpX9i1TKRcIv1Y/c2QsmAmC11/o4C0EzrTxGYYjuQ+tI/XOmqV0MSdf+AS9X5pXibxNhb
IOIDeyjj7RBxHvWKtnmxONj21eZ+hCN9bryny1sUc/S901wKtE1WHkyXuVC+hYr8af87F3q4ws3F
w6XqgUTwdQQNYFHJVtF+vpnlN4fQ8CpS/ahsesitsG7zt110/p1c5W758dSuE7r2lG52Ft8E0g4x
baPtS1297n1VxpGsxfU+pXLmiQFdeu7o7tWRrG64DgkhqWfuommAAFMNkj+ldX8z8TDmtKskXfSd
pyoYD1ktAWFOLcBypyGydkZwTya1dMHvJSBiPwDr7wNUicvnUdw6j5KNil8z+QQS8oJqIZiblnAF
6A75wndx2zyVhfWhqsb84C3rOybSCsGSGz1XJpagccD2rzFAws8aOgaU1rFJCIUCrymC17km3Z6P
MYAdBHYqwhZ4mWn3i9dKOKhNmosGZ7nmltZjdqt5XHKJLVCR+8f27Re+2aqHeylvxKtUHmZ8y4Qn
RvX0LWws+hj/UM+RaappzVcZ9zMNxrIDXCjr+EfPcHm5W8hpNeEWEz/4ATHwYFPTPKiX/vztTAn6
Ditk6Cz5nrNobqYgeKzeLmtwo27iWqiSOtYTkjiOg3SLJ08lz+DHA8bbrQogxmwrAqQrvx9KETy2
Z5JFbqN0pgAoTtAfZosEroo9IIofUJztoqezDTM9/xJ5KyDihWC2aEc0j3bEL7njw9dPfrSNOlcB
1pKjPhDJZWa8kT8SbO++qltpugKnxsF5vjnRCKEHnMn45oic/kcFxPS0riy/XxpKaQCLno4IgSqw
M53R2hCUOFwt0gG5ULdfKjQM+QaljqVl/y2GaGaok5tq5XdhRgjti2m2ls/yhUUA1TGhyvhaUsOx
+qAyPrH7824EGXH+5wiTwRjBSKibYabqog3gLVlPufh1drbtfrOaG8eOEW1zCm1qZVnJ/ZaGZCnD
984hYdVEzMWJ+RjTShwoBiMCbJ90rznFcFra4jgbl+r++yI1YtLSCvgg2NqJCajqLuRDwgLQZdlc
E8kWUjhwovAvsrKlYtz/im6CKDkPlse2cGwZDF9siinPPgSfS+S4wNxm9e7JxYycGova+J/SLboI
CoCZuyuMxlUn5oCRXWWImdW4yBzA9wnsvBkSRpwcn+g8xT6peUdi2Zu1L0yaBu9T32VPOJ2ZTCOV
/8mPmFzLXyLmHbYmbYQJRHSgZVc4mvWdilr3GnqFPeC60wlMkN4GmvE/olnXlAkr52Ycjb0JUtR6
GNYf8UhWs5GJ46mPrp2YqAh4hQWjtxqnCvavAfsrQCJRmIDk39J5xA5Bj7HopMvLJjcUctylSahU
+WiO3WmgIsZB4NpmdKSQDRxdaXUbO8SSP+V1oloUCDuG8Ls7gbCBZOpIpY0uHLbdqRdOdoULQ6e2
2tWw8Spa0V0NrodI/VXRZn7e931mtuJtJmVv/H/3Hx1bV9FSVTWiiT1e2vw9D1rSd9CfoEWFK38r
nyREgbq6TvdKMhifBfh0H4VQn9WcLg8YVXohfNaxgJ8xTIkyEuwSo+M3kltdsHCzy11co465ssdV
MDzs4x1qBVx8yNDJSQthD+a3oIX+DKd8i+qPDXkw+QDOwqPVkAbKSXuBR2vrdKkixFz0u7mwKW8V
ebyC65X0gT2ffpb3tW/r6wPunYu0klTDSypzYjRAu5owN1oSFsXmYjIrio/fnppIXwQVpDvS3T7Q
X8NOIyj9g6/dAmhCHuLRLh6ChY061xTCLd4dyG/0+CEjXnNfYvKNngUABPZj6ak59hmlJTpadX+r
9tq6K/XMBlp3M58CK76bXbzdeHOzvR9jMBa29G1jBgcJovngIiESu4SuPX2wtU2A8UVBho6Toqz3
q60Ts4EtATu4F9Ygmx5nEYx16jNhnC0mfSwZtf95BgLY9LdsNRl0XFE0KZ8RToXFa3EHwaHAoNYj
4D0yTDcXhqYWvhY45o5M2C+sugSuOBWXMONBRLiRl9Nty++FvJ/3CqRkkivNtu+0ddWz1lwBwfNS
tJEO9CztjNg9gMXP8wz3OXzJtjToKq4fut6Fk8Dys/e9OhG8Zo2w2kZ5PRnuydeQHAjxfE0Mr62R
MC+Nut5kWN2j09htUQsjLHmDgDnPq5ZksfDIw+JLskPBh9k4JG7aR2OzQqvOBfWXMgV7zw9h2h/0
W1D2UMOjmMw9nBFNHyhwoexEsXpOPnvfxZEDkv4l2LXExpOPppoMtkdtM8IsGkmjNRekfmiFLPN7
T9QhYJkpNGskco2SuAa/C1DCPpYleGqPq+8sHnOouyOfVOYFbHj0CxNmz6Gg/pE+zf5yZ0a1XJZA
+Ku2XH43HsAgVTTCktcJC6WesNow1WfTUrxxZpFM/zL0OzwKx0yzaTk8hxLFCc7Mo6X4hsXX9PTq
F0odHlqYqe+qGsbSU0xS4mtv7JEf44fCkl9GW7rZPehc0dYGM+Y6J6yCues/ZniBiYskB7XDvnxz
P1rdXYfIPNiEU8OftUgVGy3pqObQeeU5yFi497JV+08xhCZex1xGiQiOC3ep4lIqm9ao6LUW8h7w
AoMAcvznNvrUwgiIjjMnx6X64B/mRHXZ1OJqeAyexIdCRwrazkfXSKxThJ0z4WASllNz/wbAPD6r
bxW4FS7W9tFo0sFwqC1dfbtzNKQsdi/jqu70T5L4GNoX304aRxzA5j7F0U+am79FFytkWdomie1M
ILd44r+dfLhkfA/YW1FLVkzYRLEzmgCrY7UeLKp4ByQBPVX4JPu6/bot/5ysyAq1A5FTrAMfFusQ
u/sW6tHbyB7WUO+nsTEaOWRROXY14QK3WlFND6kzCYg5+jCPZCH3tUfO3dh0t7I4d+leSq/9X4My
9RY0x4HcD1iH5N6YgzakIiOw9dMc0p+ZUKIoqaPlShXiQ+ZDbJEy+FIaQMY0Heiq7wJpksuG3uYR
iBm5JwanCI/XWFQ8zvPWGvJSGl93+Z5ilCK0l9C4w4nmBn8ZsR7PAmPrsH2P+d2/aL1HHypGfnqR
hH/Per47hT0UCX3TvX6wmjLnMgnGTuiRKpX14Nv10v46ksZstNSjDV/Hp/8uhEhtPsmXfvwnqy9Z
jU313XwtTFGiY655rNvLE4XkhwWXmRvyJl6nGPBdfoSwNmulYMpkB6SJ159K3phu5YC7FnHn/AzB
x8/9ebWM3nANh2ZyjfCWEQCPxX8wIv0mxGnCbHkYogFrkAQrdYzdvKyff/WE2UkbUSm/l2je5upl
OsV8ZPPFYVaEO9JkB6ySdAu0aJGWnanBJJ7XTNePlcIZQgG/5VTfPWgTHg6JBFTReYgr5DItuJTC
WT/pXYi/QNkh1Y+8yVxTDP7GDylPPCm1uazO1cZUcuf8+Cwe3MovrPkqokk4iNglH4/9W9RkSxxU
IFrSLkpGnWW/6fLgbmyr5D2iAWnPnOgSVNgV1naaqcrN3OOAEOJiLraGDSerXIZlp8K4JP6y1MTm
IenUxUluVoWYn+g/mnBSUk2r5s7D26ml6DiQ1izdSeUU4s92JJJqsy9MBv08El0/YhsaiBhBDBW7
f/2kYVk0RwNDxveCbb+nfPUDGekXWnpGcMkUDmhLS1S0wxmnd2Pc+k1SBrgDoa7Ihu6ZyJZygqo3
tptpOu0c0ZAsibHXab2sBZyfAgfguV42ZX8N/S29JBRHsEiqdaBRkLYgoXEl7mZvM80znGnTOEMd
UJITF9UdQ0iEf6VvNhh5DsI4zDR0vm4vYChEmJ/Dv+mszH4K9dW9jvJPOnxeWC9r5sOuGOplOho1
iGm+VmAg0ND/4vIsOFkxtz6j5fOAAlVI60OSvpGrXbPKXRpjP6u4X/krFL8zfa5V+Ff8Y/YJCZyT
eQr1zdx7sIdGY2HZ/2AbQRHvYp+5TSEfqHaqtxBER9GFC6JZvcoi0a/HOux6vXC8IsR0671b4BkX
OpBbhFVQ0QNVn/8ejiwRG1lu6ze6TvQG5sioYor5ccF8skfwRzZxE7SfiERvU6T39L+XIqDUPuWx
gNSNQc7/LE67WS87Q7PwVfwAH6XZ6TxlbNu2Dsd2kra/b053sfHVSPtcpFWSj5wnxRPxQzMLFg67
1BtCZfEE4jrGymrccOndt37+ZgWMDsuYELiE5x9iTJXkyI+RHK/1cNi3ViZIhmYzRKMA5P5uRH+N
+qSPdD7cfAzLvOfQ7fPFQ3UhTEwhAMXHNMl0cgGH++wAoAtBW+0HFzx+iqFLueJAtx/E/EjpiPxx
Q8KB2qofMtLi4mBJdiVaQVqDLzzNons4GcpIkFdv0n3HJHcdlhAO9Yot8aaQps8bi0sm35N0iW19
5xSOo55fr5I4ZeX+1EOpSqTfagikK1sbJxK05RRS9I4GK2iUmuTj094j0N7ujsB739sSTcxmix2+
3ipy+nXUuByPC0csJbNfH1tkB/p1vW7gMOqb8Gc81F4HC3Dhkms6o6r2Fqp86Tw8AK4uFUYZcQcq
Qt/88XTmEEWXf4jUY9svze5OQMoZfB7nS3SqjWbBIcrZZSoO6Om0QvyjcWkfJ96nSCJsXG98tPK8
N3ClI+Gx8CDrZcgO0l3mnrRo/ewNX1gLOet9p+WUZqKeajk55XWib+V4mr0vtGpM8/twcJwwVIM4
a/b2WpiiiX3SRxEF40Q5mQ0UP1TKVrZMD6tiiB4skbFVfDC2Ddd+gH8Ih00zXLielqpf1u1GOcz2
ww1ThGH+MJaByYQY7GWtlFkayZg9aeGojJtR63EwUKZeIGKflvk64h9QFIAcJzesYWgKFIuDmyH7
xTM3ni5BZHIPh7fBnPhRVP3PYgTzuG4ahVBaBu1/o+dpZSPP4J1FyuNgUFWP3FVkrsO29YLlK1pL
ShPZh+3L3eTdZUnDhK814ROIqGHJdV4SzKkMZlPE5jO0RmBwYVn3dFlfcHw/LJqR6yRoqmw9i6wc
GE/wnaGZyjjt0Vd42dpFA/gN00HTF/2Y3fcOxgB1vZLcQbuhLlgD0Ru5A2k6PY2UMCk1xVriuU7q
EbVzVwuotSx1MBNbkDBiG1r8BEvfP408Rgspgx4nKzSKN2AQUlZy+Y+GtICiJNMFlyfmlB1C+h2m
wPXsimJkdLNy1bwG6rna4QZLO+FZBxXTQStpZ8J8MJyccHAjnu+iSuYq10HteDiw6IChgcKrZRUq
KlS3qaC+zKr+IIHUd3QNFm5Sjdf4obqdW/9z1/5+4NSlflfuMQGdFBU6B1m8+vwJUKjYd4SPG4Ti
n/GcbXb5OrA0Txq2ISP7dLrYSaG5gGmwZGtyh6Iyk5lUEdAav33QTGDK8v+WXxYzU1Aj9Mjz8lgh
7axG2o77COfz8zh8UsGa0DLBEv2MzHpdDZJ34NIFg6SmgcH2VfzrlWSQ3dW27euiIYtsSbQ0+z4V
XF2pmj1+W05MVpouDmckMKyqwBn1ERVNQ35W2LMrg1aju1S2eioWjzz5f2Y95MrynzIkq5+gBY1W
8uUy9MLjPXHLO7x0w/UgAQ6j0WHsaO17uTEC1uu6UXtmz+nqNE9pnXeFKK7ityIyZoRCGC/GhK6C
sf/ZYge+yscq76/BgW44f3D52ZklftoiDybXlqttAQe4e6pFLrPlIwv20FpJH9oijK5WnQajsQl2
8k5jO8HnB1n9wmAHMp+0IZ90v9S4RAyM8+Ii2kRo0Jwwit0qKypRiNpILKwbklgo8kU12dPDJr2X
UXbrQfxwWvErgqBX+hDnm4VVLCS+nZTDxJtc/W021ILEpSyI8FCNPw9AIc2xtthiNb5fwJ9XQ9EM
vv7yeW7u3nKrCx0gtZfZTtzSu1GjoHiPyYX2ZLY8TmyBZFuE1HQiZ2PvgWeeFkok5oS0KKV2zIJx
KQtReQh+qbVB6AID3G8dgtzT+VHYqTQVO7XyeXd92oLy9fY+8BtvkYJqGkApOpajKfLW1qKeAROF
00607W+9KwCRNfcAieLallw6QqCmz5zUrrLGWXH1VQi5kEE0RgDsZAKa0d6fHRoTEG4heVp5HsLX
z6rxHYCOsGl5PIw8OvYFqalj44LF0+5sZSnS8ElyxFcV4Ivwg/ZbX1ZDjpxD7bv/QyorfCFN4uG0
mrax2bIyGgqgPUXgilEvRgxPQuJpzqUlUAOKU73XfXDpuqMRL0b+F2JNJLwI9dZisd8gdzkX19pQ
vqKXMmUZIexF24iWi5aLibizRPZQmPaOwBu5RkGJ+zxmxAtCPXiBtuXqVBEP/KaS6WMaRd3mcxij
975LdGJlZSwI/77E+gsIhzBC1kjuea4+iy/plGeGTmt0WzDxK1vnfidbLdGgbuqbEItBQImsDst0
9VIXogIKnJug1tkE36yiwTPuUm2JOKoUwOJ4kuTcs9tfcua8q2V4AMwIFcd8s0hnLgAHIGTDLtYR
CbL5sYKMXX2GU67pJV9h6kfPIqEcX3hrNJnjZVf1zbxrJFb05q48H3ULPWNvXQvqQKy27jMbaViQ
f/LFq+EqMRTDVgcvp8sxzaO5/zI22tizASVGpzHaK40Tk8IWSMEJsfwdwf2HqkvRs6UoPNPiBqHY
hCEm6gI+ycbBzM0XgU1mUC3kycMPEmk27p9LpFf9BtBdmjTb6DcXqMYOpy16ISfpif2ZsAN9pnIw
fyff9T6k7lhk8HH81WKbnES9ZYdu+wwIUh6zgnuIQLW9W4KxiMVlvb2GUuiAkFdMnE/zq8biSmQq
UGTfkhmqTf98+XpsywrBIRlqv3by2o6FOuzg1QRinVn+m74mZd926teu7wh6olewQBy38yjKi1lz
qiqIqCNbsi0Nra7Hote/+lZLZ+EPeYy1e+qH8GSCQqh25nyDWxoZPfGDWeUz0vPd/veaV10BKzuF
S9zkDJFyG6YLDgJRuAvTg/3YVsGCTBHC4m1yynhGzQTUqxW3NcSRQtG6bRvRkum9kJ5CoVkEQAuN
9Gs6XMjHQ18R3vnKJUL5cmRJg0y2NsGdRHqtt/RersTSIgXi5NO/hACTIqH9BHRGx9P/4cIVSeU8
D2qs+n/Ma0MPcRQK2J+wyGU/IyhYAVt3BGYABvKV8Y4CM7t/Lyp3xp+M72nzQK3YGHKc5v7cInb3
eqXw1CH4gCcrV9U46QMsyvAy3jnooTmNx+A0YQgIdgTRjkFOl4V9n7wHFzbQMVbPwA0Nua1yMjG8
duktT7Xqw+yp6Lvh2HJs252+7FL/UxUneITbR2Zm1KlB36wkTLZWxhleJRoI3uu3ufG7GqqW0XW6
ppak2Wzztu9MxW9vyP2aoTuZjiHqGyiekwNLcEIWSAyCPkiy69a1m5HSOMj53Do2QGaA2uP312ij
pq2Hcq6mirtJSFm2H5Jw7GWKQzuQ164oKI9muG+kYj9dHnJy3+JQVvZGel7Gst4mrbzpFSqfyN2R
xEGTji9pFOW+wZHewTZfcup89pst1lLT4vnZb+WEPo1AQerll3VmB2eHcvMagLE+702Tpy+NEHm2
fy8rWfrTXyf5T9NHZDm8kJQ59pZqX+4Hl3mjAcDrQjoyt80/uucsj7Otr7kdJQjI8Bs1spWbTrrd
/S6xTRD9A2Io7pRCrpSJQ1SoC7n2zc7j0QbvNYVhpaq/6xIFqTcCY04+y90Owd5hH7czEYk/nEwZ
vZZ+l/LQfL/2gdyikN/x1hmhnZC6HApppSWI73SdmwdM1biaZHfrJ7X6l3c9rL2yqyX4/Ujxsvlb
I87OwFytLwC5m3E0nNjD87rm3FrwO9g67DsnW4x6XHtuDkH0QjXXSVDSwSK7a5neUDw2PKhfaLP8
bx8kk6nR5V4tYZYBJ6ooBdF8CQv9GtbU0IX8EuImEnoVeoc3TsxBq/jYP/aPW/ECNyoh8hrh9lpG
+KjZYtNav45Ol5gPn+KrX5eLsyr9PNJ737YDxVJX/x0drNOZi9FkU3FNPZ6FHIzMt39pb8PwHAoD
nIjqb4ix+mZ8QMZi0l7ntN8zhXLc6Ck7ZUJA+kZ3f6DyXqIPdZSyQXPAYEEJQ4+AVkyUAe9owbMV
+lQeUPuxi6nDozs8ZQv6/S0wgKMJWkE37TQpL1Tugp+rh8durvk/Mx3IQvKNV595MPXIwZsGgpNu
/D5+Kh/ywWvMiyhBAf4uklgAdnmgIWohDkqgeI03rgpPq0hS/r/d4ficNtn0rLS212lEgTydCIRM
Vzn3qUwqnDXrXH3mxER/NLc6Q/6ZlGCV/Dp6QKZ2aYEYmpbUPO4OnvXy/m93o6ONf48aMhFvgyyE
FhyZd8pibLAM9Qhymm6XifaBqtXsyjn+Aa1dZ0obo1GJPjCVVP5vvdy6+NJToElvT/MB0pliUQmZ
ALlAxYKQDafrVniCP6A1qo1HN3S+bj+pxIk5ZqCUNvaTLCHxz912AwZ/whnQdRteIEm6fcHKVkAS
kO888V2GkzDrC3QqP2RFqFlMG+nsc7w/BTak5joi3PQLslEvePvgn76M5DpeP3vqVc0cUprhExea
WpTmpbWlczizsuWXT0WE4YVMHO9IbdUxsDXwh6DyZGxX9eVyZOggBTR2n5hp5xE0EB3Z4cynJ+fk
DFZsvbCXbHFkqBLVUWs7fS0oSxx2LxQcmkkIvdE0hp3pq4tgYa/PBRUTzoUWooozmUWaVU5VA3on
GAWkoDihFGvR1VXUe1ZS+SoIOa6T1pvhhGs9niPx80mgN3ZMDwWQ/t3rmQGnKAYfy/wdJsaxkKJ+
+59XY/US881oIgvZ+TrE6D9N0JupHa5o2LYxfwdtoqbO9XzUz4i1vSQsxLoUhYKVajvibq0Loyzt
41X6vXKPmDFVrv3hN61WKkaiHDzxFdl4upqqbVTet20cSsVsYfOtb+WR9nGoYz3GuvLLJonEk9xb
u/fvWO9xTkl0LEX3GGX3r1zVaaW9QP6r0fB7AOviE2/tsvELWnpW+YAZopXpCPHGBsgjdUBw11nm
ChuAd5OSUeG70gRRwlIR5h1522RFshyRvvkZr8lcYbUsRAcO5QT3vxCvTJAf0tD5f1sgCE8Vgu3f
gwAd/K14WWH8oX+KXE0QXiY6Sh082NocgdMdJSVLQkLwIcC2XqFwo6JF8mSOoZk7PTyvqnDKvVGH
UAAy74js3E22AFcMrZew8dcPjEQe8J/9BZ2Fd20/zpx22rBQhLVokr6U8ia+KOP2rFa207NBeAKB
+oXe8HMCUtH6e5q0ZbSNMFk6Y+6ihgP8a51QyFuWZM+EQsqdWoEVIFzE/rGb3pyAygCL7wFm/PaQ
AuYNyOmXc6lO+6BqYdGr3KSxTAPZ+EI9YAumZVyPzjPjKWiz1anEgDmsowKA2WcPSU6UVcOBxzni
26+rLYtFTkPT/lUpgUseg9aG705iSUSYYk721BrPWZN+aKOME3uWqXm22qF9Nr+1tzWpvXM7UKNT
547o1Ch2mqfMssYFZ4p1+SfTIVMhN2wFhyeops7gBmHVQGMGVCQicoUCPYaakPDE4Sn4/b41A+58
jBd/p6AK+is+ZlnQgvp0hWiAlVbTsNrPe1oeXidr1rylfOe7zIqGlNBNJQzEyHiXuWNMm0fM4AB6
5fVLFDEh8JcVYOwWpnvKMHP8t0ODG+D0MRmAjC/d0jiGHGZZVLPus3qFFxAIsAbzSBTl50kMfrDb
uR1XEnYrwocun9+13ib2kijUOUA1FTjEenFdd0ArJVgSQCpk9Ro1nz5S+CMwaM8Y1IsJa0gwsUpP
lFWPrMn7tZ6xR4ZO2Ex3Q0jpkhJ0h0pwns8YMBf8ZCbAqHACPZb6TxklI+dq8DdLWIF5B6n1/932
04Q5amItPVIVI91AzW7KFc4ka5WZkAj8DnuzLQ+v8dApWrLrvNVr3HnHXVSOv9d1tz7Xjx2JwaYP
mtHUERPK7fmXJ5uXcgLjLs0FPFPB8BsZFCf7WgNLXiKmYeFcujR1ttbEwXYXs0ntgW0ZJTCrmyaA
rPb3HmguO3WvZr41OMyBH+sz6Ca4uZEl4IxZmagG5XuoG9r1qyuAKj49MDuBB63LYLGA8N10TyKj
n/HbNn2g/X9DRENB1+o+d9W+7sQGsY0ksSttzqF0WLU/Kzx7w6w6DKEA6ECrlVtqaSpuqCrZ+IhT
DPG0j0XsMECDVn1eEQgRuYXK4pPmTkM+5hXypmYLqHibE3qcexklxyQHf9FtdldKxl0wWLrUh19K
Npz1ErxsL2RZok3VhF1jZHex/fDlC1trEjLwgKQ3jaXazI6/ujdL2zA01UIlOdPcPgI30j/gigkG
uAiVXufbi3RggHXw9L3wdSGh7V7p1/d8wt/F0V6IHpQwch8387F6VvOyJp+/1xKfdAlkoWZB6gpK
IaYLxM4jj23rqmdUJed3ZsjUqB7GoQJjJzhuj3S/RQrSjOGzWBIscGKLmFpnySG8r7am2Z2xUPBY
fjDM6dhztKTPSKdbA4Ms4cnBQ/Ri1EWSacgzTz6zH48JaoJevwbDrfRTGWbdEeWnA4ABZWvw0Bi4
s5sa5YzIUlODkcvb1dU4MX5+g040YO3hqe37zJtQhxKXed+k7LYZF1OxAJ59l8s2ILWGsfAcaLst
v67DgSc6qL6geDUeI2FHruIayqVsrat1eADvLHbbiyV0KjCLzK5q5F1NbmOu8H/sF/tJI/CfT5Rg
ACA60KNztgLQmSdhrzvrGbVYxnAiQr218t523RT0F8sY/ISAIqGLEbiNDv+pzsZkixIz7V5jjvty
1NKy1nwZSKjk+WTr3tkRXmvdwoJcUUozAwG37DTPSU8ipBLxr+YGRacoH0dmyf6wSv3ENYjVsswu
aOHq9vbHh8jODUzXupwpLBVxqUYRDFCq3uhw5qMHBQ6Qz04t8TxEcRPZwR+vc4t4JmkIx6pjQ6Gn
N5MWkmtV64nAP0L4DlI5IkGVEZYnPv8u2mahxsNaiyWMaJoT2T1ZNwl+k8VlH2BZ2r+DsRG0Vm8W
S2zF1xXxHJAwqMMYYmpUu65Tc2dN4w6Am7V5gq51KSkCh6S9M99woS/utGMupD5cIrpoSJPECpBz
+JfSNa7ANpKqe/KyJUUlRqbACTMMj8Ig6ojABeUZUnNjbhYZq3vDGRDvKdxwV6p7AllET5S/k4Cv
Eh9xlsF+o7k6SwBVZA07UPoFmbgg7eemy21mVK1uUF5z1bxdWOTp1ALVBO7XlPgtuwlKdH/fDLe1
zaqXk+LRhZdWEZ8TNrAtS1KIhvBqTCRYklgr7tzeLr+A3r1WutlnA9mehabHhq7oq3Yev9vzz0Sv
2GNC8voksZ4qtjIfYH5UcJ0s1Al+bz7zbzUg0AStuA0Afog/oHm1CeuIMPhF7+ZzWpRRc/7uVzh9
jEEsR8ULqVzg6B1R6tWM7f+TomkWcMIGjKL8Sl++0SKgWh7ZqH61WaxtCKjoJsF8GBg1Oe1VRG4l
jsWebUmWHmDMHgSFrCVDGBDtuXSg1SMa+c9616AuqNj/epTSFuw/+xH4rDWURl7CpxxyIZ2F2HQo
0DTgKU+bCLnxFdMd7G0S3qg+Qw4yIPqHMUVDHjDsPi/6D1t145tMlo0CZ6Yj9eDJgYPGveRq07cw
A2VDXL1soHU9u1AHJIMPoclnmSdaYlofqQ6MaoIL1MvxuajfHl7gAKxQ8UULd6YwsodiDaMmRzg6
eiskD2jLjgESyO1Ovs7fTsZJcy106M217gOyDk+gA4WNm+H8JIxJmGNP1sfLM10NtobA7AOjD5Ee
oJ0jGAqGoZCZoo3rGXkBztWZnxOr+pjGp7701NIg35iSKOPonUUtyUnF7PE+IMeY1nIccUGDndyu
tegrMQUnJovuwKfAk/XjC6zYAqwopdDZlS60UYwuEezmxB7ygoJO1uL2WZ4jARK6azAS7Y/MJm+L
05yamJHgoiG8O5UsCdGsDI9TL6sL1v1ABAZAsN5x1xARVdf/9WgmnPTW3L2fCZcRpMTU423XYETa
NVuPFArNvuUbMb4qjrEeADt+27SGK81H6GGzLMUU4c4AU7lrTUbGwFZci6Yk/2wdCl2WDH5rJvTF
9VVTf2PtuftLL+fYzNjRNGp6nq9ySSPG3ooLl4a4Kdjf57YvsVhDAnCD2TlwV5rZglmiZBzrfh2O
fNOZPWvb4L//PcQ3/m4flMHsJGk2XoqVYnRWyH+/iURIca5QaxWZYN+kAGopN17byd9CNlYLOlNr
wOy6K2x0WnvJLsanJflqnrvaEp4MRgtbEfZUiY8F7nbDTXo9qy0S710Tbre14poWfOeBlLf4AcQp
uIz61WvVflF+2v2JhO+5jzAGyz9YhJltIaB+BVm9Hp5eQOp4UG3VvtM5d0IkWFWs7BAmgsUBri6v
4nsvX+haMg+aQrXxfDQkusow9zIR2z+A10TLKqtX2fQWF1YsjYMrWQz3fPmc7rZVR8g1C5woFEpN
ABls9JSznGGNedZUyrS4HndIaUZAfn3QIWE7ExyRqd5+VagL+NStfzjgw5FpjRob0UKFpyg47KD0
jojjDvGPmqYSZnbjMIKujqBxO+74saKYrogWyg9YJ6xTrnkp+KQR/FRvpoRddjdDRW0xyPc4dO8E
zYuiBRFEGOQ9j9Yzu5Xheewf4Gd9+y8MswzvAbUBiVkcG/+XIYpRa6FStO1MPI2iP2Y8E/RpQpsC
pFT2H9ajKxQbwbYPQfCX9Py0cfdqNokd18wLBvGRbpeH9P8xO6Xxpjmxa49S4T+1Z0aU36K6C18B
DswOGZrThUVcKZoAtCe5ChbyVJ52iWonhSniw9DNBha01PiIAvQZWHfFvTlfue6xiMvJ/Z3QIw5B
V8LuV3Tsh2F0LnGZ8bCodT3meBqgQXpxMrrVNmk8SxgSKn7nxjsSox6Ad2imSU9VJ+/1q0nfh6rW
hwq4pN5VAnaQtxf2VH9hWjGZnjv9DiNxDx39F/5vD92m4AtDHjxOfSqx7Z997nkDrq4IcLtd+AfT
tdVbhUuo9LhuFHTrtp2o81DK6k2TRzCQNk4LmpQHCMgpfGyd3i+vYQcIxNugvi97kILXdymmr/Mb
eGmtmyJdAad9gw3d56R+1v7Ipo1KeW3iJKH/ZTKZhaaAqQrurxmy5KqYfftmEGwDVdiswT5I7MDj
ArCzZsi2YmQ8M203cUP8ZrOvT5DzXHKadQeJ2SYDpaoQbb0AJMw7vtx3ctsOf+GHRg2ToisSrLyI
GNtEsBiaQnnKt/pO1n9HQ1oofyZWSeoakXHoIzqqwGQXicicJOm68swt8VeCIrFgbu0dTzYUudl1
eRlgfIcWDcs89MBLk0t4kJecFfgC/yuEkg/WkBUMH1NQX1Uc1q6hDj2s4D68XzNYByWNj8U33VVV
g3diiJmRtMk/BlKyeLBww7xOPGV9APGCTs1wnPw6o/etiPDf/aAf3mqtEt7L+c9tGfqSex4STwFG
edxSoX+BuJo9ugXQ8lVD7sMFatZVT9XBgub2enMPKL1lQgw0F2eU0jYSXGXOe/ZmADFNxAOrTDSr
eg9wlTr5KOHvD3L+ke5k/+8mNKLT4DUAjKygTBWhQxovRg3dMXkCprErh87CxFSzJNa2MUw5Ys3Q
WQgLY9y5Zi516wMvte853nEpJxe3Xbc0GP38G0s/R+pvN5CUumzg2qvJrD8uwT1L07KrBkAOdT7L
VUZV80URaoOy1Yd9Ocz7CatQrmdyXaLgs38sXRNkuULoc/0dufYf+P/XILnEXMSgixf9mUjewYFH
ogKzaQHyXFPl2YFKhr5SeJnkKdULLRpQJwiY5hVBf4xEPaqYBZg5NhPN5rY6xmD0D/0ifrRKlfvZ
BfAjv5tztD9CAHGmsF6Qd+qfDMKzk+om/YGq7Df1pMIp8sqcahjylPQMqUq9XpEl5QtmOlnrT/4r
sYAnNlhz4gz2UlLrOSk6PyGQWjxFsPN67anKkwCckMX1kXYX86pedTr4t8ihctjwzo3NV5Q+N5uq
nxXTZ3M9yrL58F78Z8dJEJS8j1WBcIfbNtQiRSuwr2lfzjS40tVVW/UpZ4PGaXIIrhzE6+2amITy
FJ3E6V6CT2XVSJ3zkzXpMbKGxSQmQFqHzxA2TPtdKw/xtwLhwvEvcjQJiXPkECaIfn+iKCiFD7Gt
AV7TICFHsLcFWecjMCQA78xOQMzC2iJQbXF/Lon2nEMrddAShNbSiZ7f7App8gogO4Bv0cO1+O63
RFqlSdTy0jvlGrjE0WD/luUFRs0gvwLAunHyXJM/JkxMtGcbRUxAU9kuME4ql0+EJzdQVsqpKV2D
0ZaTgwVElMjfyPvfvg6ZRdvCvnlCOoEtYBam9I3ntGDRq7wLg07YWFz6VdM5eidBWm+15yK5KZd3
U0uLX3mBInLJIOdPFRc3hwaOQ6u/eAqM+IlcRlZIT4a5T1v9PgCiuXq28qYuCsvssgdkzXTTjbIG
0ABnvPF6+0iFSnQcSt3ivgq5QvdqenWpQrJTlowWg+6Lkv5aUbR5bbYACqx4tSsBzJhSakK0IQoW
OOlHpRebzfJ84o3YcKBaVjasU4tmOqZn9tQX5xpveVgPaDjsV3EnkgpGVwwDNpzissANeYaSzm4A
Oj/GxNM5mbET8N5n1MLskhwz6RjxOirWX/lmGWdYeaCcWcadORSwP8buDXCsecgMwr7NFexjJCFq
0SnuMrcy9uX09qp2c//rBhGn6CWTVgMI2U/+J/RD/9Y3bg7ZugiGrRwv1uo83ZjhL5Cuty8cDrPE
Oe7+3xdbXqGVX8DrAhhsfmUs3jOOKHpQHaUnq4Az/RBsA5Cyyp03752W+iSWfRuB27dA7m3qIEXu
BFHUiP+U1R7opVlAt2bBDalpS+m/15USzbgI6rfFyoCmwurDsGb7kpSwfmgBB8oQFRXVquec512j
rRJoafjiR+KYVPDuhjcIdfWTQ5P+O4WEoasJh+BlYAWeNDVU3oOfPImZCcyrbGcyvP2E7c+KwXVO
/RmexaWE09NgJrJRPzrXQ+sf2zf6RbJMp4Tv9TL16npoavjrN/+Gkrb2F9xqgSTLrOUdYbFkwpme
3sCPxwkjin7SR6cMDG8MBY83rtDpO7JkQI8BI2Jv0nixvuZYPQUTRy/8GvOsKCDSh8/QYVfzd2/9
uFo5hqhWkUJMMJz0pt5LRRj/tZxfackEEMJGvYY9vlbyTju2qQhtguZmA96HZ6EpyxPmju2U21Hp
7Y9KNN4QjDh3RkyhkTN2lbjGjyFA+3Z6doqug/9bFN9FAwbnx7f2SWSdUrNCkrnZFGyIdpBimLUc
/q/39PyRWpAzxtvUMTL67WHhwZ1/JxVmo69aoL6qpmqcJhaWi+LKOPL+jyvkRe3Atm0CH0xCCU5o
9sPOb64EbRh0csT4wQuDeUBPEgOlAskBdSfCfed7SGjAve6oxgQUiJ3sHhAyfrAdqBoCJSDqVaDS
moXj0eSX0cfHo1v1+Lvj4mE30+2+ulYlMF59Yg6Y+FL74gwdrfv1DcY7WUG+QQwPhkppXM3T2YVT
NxwmdDbGM+3UuMeZLjLV6tz6w8+JfPTxPUDl5h3gGaGqw2KbaQg0Khv1jsRheToytmlDW/bYZX0A
SFBfsNrtXN3PCeK6wKQuxZ8Ez5bCLs4m/O4I2laAjhe3nakhA55B9p/xo8aleLPA4fqzKiYafN5S
mV3Edo6TW6hAX00Hk4EgAHCuAOU2IhxNPHYHbzDNWXe5EUb/2UdC7d/XivO+RjcCZ9BQbRSwRRj0
GXD+iYUpvjy22n9o5yfIELpgfCgUUIz30LxbkfQBG7klR8cjeZX61NnwIIAPZDAEgBcRcqaCR5O4
TmRShnUGHw0vzXWaplgdr2WI8v7rQFu1y8T+UFkIiEHEz+3vZrMWZ3OMITN6tNjgjiwqYT7uUqsU
MZK0IS+yAYw+NpQXG/XuP56aiCUg+kFa3j0uJs7UN0smd1hJaXONQp697p32b3GboDr8SWfQuHns
GHFZ4Xg6IppOd52YmsgFtTgwFNijhhJDsEq1+wvifI2VSn80dYn6I9nAkpXLh9/xls5OVcpZ8yzP
aN72P8UCZZjLASWmDPpHiZCkn8tIt6MUBOGKN9ZeseSWtjJCDVSBZLsTejSSYarqaAFeX8MbAU64
OjXGR4uLwoWSafrLSQrAAmyGOus+9vAmshZYRFO++QaVg4CeLCzHXffBqWaIN+yhumsl8+QMQzjW
f0QlgXJ7kjxCPwDsjKdctGPfW/Ds1dbcU/bHQEB1Gz/iOjbEMwM0+W4AvC6KWDNZs66hLF59fbrx
b388rNs15JQD2jsK9QEytbVibnN+3pwVV2ivj2XsRwon0hXqRB3SzL1Rq1Ipmb9HJU6XtkM7SdhX
n2KGaHMgpJMDNXg4HGKBS/q0CkfcLdmtvaV9Lm2wFVqlSGQQApJXj0Ij9o0OstX7+uOGf6p3cWNE
Sj3hFcg7aqMyB0xOVp9qWeUDnrXbkS7rneZcGI98dvZ0a0GLC4h/2MSC6/brvUKf00dFAFEGGtnU
dBp8x9Pif28yvfTReyF2HFKMgMcoN2b6xN7TjiKLyLHio9+IW6oHymALJsI6XKO0xusHcaRB6bKF
vg76BF+bYAhPNM4U/iG+J+UVd4FgVIn8UiS+32DzYqlfEvB35CoIqdsl1RW68IyGOrDbMDYAXVcE
ih0nj5hauS/dC0ZpihLpN7Xr0JSO8wXqZJ7faEvgr9mepPQ7dZgGcFKvB6C5mDWJJgiXqTAKrgoz
r21JnMKj3yITDoOKrJ0PdMid9cFQZFUncUUvTTTWrq58Rp0tLNaX5sTKPlOLUSgaopyZVeESjZgv
FbC/OjJEmug2rARPO93c4RwTF2Pt210Dl0i6lV14Irs4LD4hQ1eKI4DoWFojPB33uiBX5bCunX8r
wtO/225tsNArO3UyWjQRUCxsKTjDwKMe8gcKeCnsJnNKmFKzkVVy1DCmmqQ7V0f+esfnnkNQRXgv
mH3+2uGmCfblY5X8c4eDPqukqpI6Lr/lQYQzDkUMIWZYfpGWHjRT4ENXSJFgK8vFd97H6Qyet3A+
cIwmeZhMpxmrR2Wk2dtQhFtFL19a/X+GX5D/QlxiGtioKgEQq4FjC/xNq7tzx2rspVuv7wCypRvA
TbIdTsZm5+BTrtjXi/IcIsjNxMvT20UYlQV/CarnbJtp07q/Mv9gPINHXKYLr63+ZIIGaxnRS2hL
rL6Gq8E2woAi0ejpNAsoLhQQ1WOZwUcSsB/QklyhHgXR6vufqymxWrOzXPspHuPhsJ73s9o6+WkX
pg2olY7ldw9dwG4etLlbYUcOvU+H/Ucq4i7RUzRNlGy3L37+YPVAXiIVxd0ggz2BePJSm9gVsnXA
/4/7tB2OREYbn/9CqHNK2AYlkN9xsRgzBzlpZfpsIUG+im1XNSnz0RxkAfjeqOnxn8Hzv2cDSVjF
IyxUYoAUmsm/Qjyxu8bpfOnHW/hlmx/YCogFglC1e0iO92KkBK9kYamXFrEwrq7+Xp8eV7JnzTLQ
Oce/VvbAY9lnrMLI+ItL0xAdOyypNnQkfdbC/lkiaAzBPKIdjN37lILLDV1FMLTo9x5dFz8KATsF
dJKi+/o/chGEa4IkT6s0CuN8HkwNTH8sGR6EaYtLoVx7VmiC2HHXuNHAUAHIFKAUP5kM+UP9aSwK
3v1rEPvca3xGhNzQendPeleIVcYLt36VW+yhh+tbGFd5PBWhOtnwWpQGzw5PPucewtJ8OTAR66ai
TageMj6fej6+fbdxnRvlEyy8RMMkygsXeQIh4pO147IwYCLrj1Dbkts3LjEg3D7ycMMNy9+W3Tz2
Ykz5HaoOvGXLkEdt2fRp6xJrRFVlQJ5WwUxpZrQz4CkvGnzi/Z6NwMldF3MMyXF6pU7fLItEFWuK
HGmO9+qDUiwE41gM2R1TVWTUBk/qpoRsTYGnFUB0Beix0yIOrPKqN7bsaxmPtW6rzqhQpMNGrcgR
DtDe1WbFMjaNG8A04jIkd773ZvjejagEZ1sLPLMJWocREyFBW/I0FebC4roDpxr71+zZlVq/F1OD
yGR78LH0IBLY7BTZUmTOFSWjh3dhzunHjK1WLm5cH5SrNy5ROkOOe7orHJOeb+A66T5/aPeEtFsy
LSIidvM23lKES2Mo8SRWuJT7deVdCrkHgUGg7YZRhe3pkMFgIXSGvryPYCnlCYCekWpL723RTccv
+tbpMidMI7JwJs5XgrsxUBQIfeiZaID6JTorDZOCz93cEVQnB9C0+Twmj244mw1CHrG9w+npYEYp
Ib9FdCG7s9XGqJPLTETsloXLixvcZ+dTO6Osau+MwS2ATlUk+dUI+jjSDLr3HfafRaiuTjtjSPd+
BX68Pg/R5nsSG62CnqK67H8mFAByBmHZNyJIxzSTvoiiXKY0kYgO8Gyv58sioupbZy+H2ZgdSyCr
KawgFcmCiKdv5R9UMzw5NXS2trDE+vpiQocVnBKQ9BQCyTFUGFwHwvHspRO0k3Vjf0HudeuX7P8Y
s1dIvahfcXOWW2P5aMPTnc8XCXDD8CAvHYEv5ZAU9nDLWZWm/TZErZK6XsmAMDhpeuH1XAQhkwkf
YeFJ5VnPvdZVYANktfifErw5oJMJslmE79KXTfzgxQ1Wj2nLhMXo9IlE7zkvPYXeOmEAFcM1cTVq
yQpgYUGnqpcYc+qu4gjy1C4J+p5q/1wJDI0VYABf5H7TAjMmvDEnIND3b7rtCpclJgnI0RySrAQp
E/nKgXVn3+AYkci4Y46Il8P/5HbH8zu0RpyGycjz7sgYkgpp/VJUMUT4AjLGZnQgucoPZhIlOBFw
SNDjWCfkK86gpyxQ9+puQZ3IPWoCTmUC5h1bMZ5Vc49f2/5deL5VMPtb8/vA8b/ajLujVPQswldt
vrMvACFJA1X+kzGI3AyqC80bXsHnGP3JAxC0lrsa479qwCdenRg/RWfhMCMku0GW8R0wwErWm6lc
2ENoQYYHinnZQEAap1iAyz6wSLe+9qpaVrSzQtHU9V3+DfJDlHniGEm4GoCsIU1Oqz5O3ioGebjw
MnIjv/nZzQpsX+PIBJdSzjOKWR5m2UHJQDahpkXBin7wpROGtp2RbG0Nx+2CzKmrC9U63AzhREAM
Zp6mp4UL4GR7boHcCQu67LEqnybGxyAED3gQydQxVw7qPJrhda6w2WEz3PZRzqAJ4U1SrDraz96v
hpvTFW+zvWmbPWFPgkxvsorfFggotjL8lk60ktkywE/eSgJc3ZcJArNoVomUg96WncKHa+ule7MP
ucgG/MimgDEIZk3+ZaQLeFj+0cDdh0R288mfl1ZtJviXLHaPX1Pb6/pAJpd1fIoleP9jBtOsa9wO
tMR0Yf3gUUWeOjrS+beCwBBhIIpEFFv3xGzMBhi6L1lUkQFGIezYW2mULIylgm5kKZhF3Z+gcnAG
8aW+Wh8wiNLtUOAPTMpEDFB9kNTGCePMyfcmiqBEDeyA62NM+WoaAk6w9iI0xKSTrTt1o95LyEI2
XcZdrKHdaobtOazzVF9mKPRsD7ZBcJeXCvJeEkqO65QKJZt7+dDhotLesVJEc4U/TuW4SOI4gmDt
tuY+psFKakNqZzba03qfvDACVf3B92DS8DxSiW3HXyya9ybKyGK4SMCEhgr0hQ9ibpnv+W4ojJqd
6Ea3l31bUOJdaYCMp2PEkohegweNATt+ikO22NutQ2hdekUofZQ0al7y2GXgQ+RgYWFfOgN+EVYY
RYZ0eLmji5+XhvustBDRek4ql37xVhqXHJEM/uFnmSPYewJpDmbmOOu6p1TUTP1MWABi7IJ8myDH
MEg7SWqCgjgV9fu5eENUKl49ZaESkhR9tMIKUMD6TOe6/CbwSrryF+2ibAxwe6lYtOGUXITdv/8K
DJfrmlC3SHJ9Jx03uxCM8r64pFB+V+5j21POph306ImS1/YSEjshyXHkXGVio8s3I1v+q1i7spz9
fkBGdkS7O+6ng4tzgyzRT5fxu8BhKw1UuVQ002SCFjFC+hGT+mmN/KIqReHQdWs55vhdPtB3vaX8
cQZZgRYpPn4YPixvHI6R0FHcrZpczU6HR4HOVTiqOiJ1HqRKwczaKH1zV5XqSB8S/DB+os9OCU8A
5z880HkE+f1rQ0klAb+aSS17f6wIL44d2bDdNoBXdFftufkWzoqS4UKC9dusJy2MpIF5f+9SJp96
xxaZw97RTC6QhouCYwPkfVnGKXg1aD+Nj984viQxJrD7f5nhk/XIKJNulhXM23Sqj3QIOKMhuYFD
9lyLQy6pemT1XXfpW0UJnikMnOaMvdHOVm6aqazlA88Z9kP8b0qUPyzOmu9P1u8UTtocjJVZCLNK
9FKgHL1dGBL1hH16pp5IO6tfhjRUWHnJBKDVWDb8DI0fjsBYqMN0M/COKqO9aEmLCGAz9WpyilJ4
D0AYsQLoM+M/UCTdaARsb6+7mbdheZA99DBe1JchiwkLY7eNA6P+UgRddBVutLkkmfOSdvvk2NOY
yQ3IXhZrVUcWRSOW8C3XUIvAM9EnNJtb6Y8THdov8C69B+25lNabh7qe6HaWgJnqf1/l1bJOMUVY
OBQAesacN6DjHme3vZTxG40B18KgbPt8rKJJBNFepjaGyCY2l8OMVlXihFx2GrGEyaGdZ1EMpy3a
JEeXEkOzwrE5CnjQP+9zQE9EvHDRMYExBmEbMrwhlTFtuda4ORUoMIn2EJ1GMNi6/lCfXFHlKHc0
ByZrV/MsG8i3pMg3xmi+7ae2E8l6/JcnL/F4LKRzNRO4ZhSGki10HovLIzmHslgVn8mzVjPKHC/V
fupXasQ+5fSOsD34LVVde9j27Vvi8xoEvvfvl38RvNsghMa3xxk3GElTLaqvHfBuHmSX0UsDdTfp
NRqqH3hdwwg73cj/6uwqae/VYd0f2V3teySrAhznZY1YBByFLhEb7crr39r55mq67wXk9RNS2byF
IW8IxtPvnNoRktjnH+dv8yghhs2dHkeAgZEg2B8jfZNh8Q7vi4t2T+aVQkSwxjSSLkJRhmy7Cd5x
EFzHQ4TJh8+BQiBjDtPuQ/W90qSojNnj6wxbJP630dMW3+sI9IpD2jwtNPZYlJbVHrQIQPNiZbmM
r5jzSP0LJxWKFCALAzLDo/eFjAJzxxbw+sGwaDAnSn0nUg1KioZBUEWPHnzkxQerDZ3dbDZaRcI+
h8AEiQpDIML99hgrVec1iIgxxP6b/G1mFctZkBfP7jWWID4O0+6i8K8TQvFAbznJkFjuRpfWv79u
vWrD5ohO856XVlGyfOYU2Y7OCf7lL/P3Mq1nIQakdQufkrI2lWhke4L+749PPMrLiUpVJv9ZYPLg
ODOIvxj4SJWauDWDHO32ToQww4rxwS6SY/4UIeUcp0UXmIcDAwHSl6DK/4LfZWF0VEOcN9bVRGiB
YhcONRbPiMgpPCI+mJ8s+qIpsHrxmz0wjjzeRTDF46sIU2KD8wbUxUXMO1dsfymMjNuubAGRVeJB
NWhamjmRU+B+y/5AxXta/jhw6SRKngPxVQXt0J/9hoayoQCzRTAfFAeoXUXtwQwPip7hyCe4O+fS
N8v7241/jRfj9/03j5zL8g4AfaXypGY3Ev+aJckNQ6qoir1+D+9vb7GhSYuCs53vWCrHFrh5I1uk
Toafwh3Tx4w+MOG9mcB0C6wD9E9JfkXm86nQTLtMkBnR9jgIghvgCAohax8kM4DTKVnZDF01uQVh
6nt/p7LX0BSNovk33WHw0qRWIXWaJpptOE/WyEFea+4v6WuE0pwvTFqaAOAp1KNEFbOrq/1k8a9A
cUsBWU+uy1GVFEcUHEKp19QzV1df+d1MD2y5FTBTQvjLgtejXTEaf0yzk1r6Gsa+ssrFIyD4C8Se
/oom1zXoIL+k1+Iec5C0OkLalort2ten29tmfM1U43JaOZCRO92rQHB0nzMV3K6gjYqRp4nlJvLg
+LwBagkzMrvuvNfG8seeNlrUFfq7YGTCkcFBLlpaMyGIz+0u7XgBEO4x/6EUq32pO1uWbUS5ohl0
iz3Mrr1SPPRuUk6a2F7wVLWv4f7YBcnrNBwdeT9qnLZN90I60n10PfGdt3JDIbltFlZMkGQTpQ1Y
8mAX75fcdl699DSFISbs6NC74hhLNwSRqldVAjEcfIDgVClR0rY40K4d0hl40xJFHgio800f/vq0
5P79zIBh+2QMmaEqF/GwhznNSVASGFW6eZkoK0jke9rVv56prlwfa7MpZEScRNR7ptcU/QxpuaJ+
VBpmVPEjrR3jJxIK7W7dO49CuGz94oELPm/sNZ45QUZM5zrI/8egulFbSrqu6rDSHhjiCLHdUP6e
1VJ4w6YJfOyTPNXm63kHhQGLBrpAW++IjCLtVFYzgowuJl7jdCbJ42Bk8xPUcnTPApjl3dE/QmnZ
IdfsDYl1izURGpPUdsZmCsBXXbH7M/vkzgOA7prBKd/GKx0OlArrFjg1NxU6B++hNbWwYT58JeRg
ODEkh2XJpU97L/9rJgGf9bauG0oPeJlu/D9yd9FhgyyL7Ac8M/ZWCk3jRqdn1Guy7hvcvefZv0aP
Hq7lUjpin/oc9DUCzQoOxHcpdqVnr3qYkccatSBTbK/RtnOYepQzWs1Tm4WV/ENGqpD3G1nDCX5v
NlKgrRiLZdRI9+6y7dokgXXp5wQwOkg8P+/E4jT2vEHvAT/h2NkT4l8MDEa/rNos+1bWcwphH+Tu
JN+2HBeTX6dXV3CiviQRTlUPY+t5qE0wDcU/vxh5M0ZO4toT5QD9DohlwQgKvRVrXMebmCDL/jz0
5zB1J+w7cgxeWmztjRpZrfFQzGTvlHvecYAQWJgc8qjOPeFsiokYoGw0g5Ls9A29pVQv9Ho9gYhF
4KoUb50ZDUhw7wi8ko5CcajGR96/yj8gCtfDlAm30nOQnvJo3pZwhyR23S0P/ll3etNiVWkT3k2I
sZo1ONpZvWEC3Xku7BNH4EgDhhwRiFIpTzBXzndO+CWxmqpnMS9wEgU1ted+WnlLCFnLZGSFhAgE
8c1pOSKPMQh5tIAVagC6HRa2Od3cI8J5/e58uAM67MlLuzE+sxbXMxSeNCbqOpaSFY8SoNjF2KPB
+ZoOHW7Vp76VGRq26jkYyuhtv9SO0TlclGcrFXae0GNl1RNjfG6pISnP8YzqDit6AIctWrXTzJU2
5hE8bfvFgsSBIbTvkvGHaf9c69IutS6cU1o5bg9nB/RnN/Jk3Iabf6V1lVf8ulbn8l58ajJeHnQU
Y2JnkNdwgucpZY8xOKTReMkzGB+Ay+aZIiVS2MbV+Mpzg7CZPaJpADEfgzmBsXtT+XKTliR1MVfP
IAYKCBbZ8W3UF3ah/zyYYIdPzQeHqFSxycY9SBG2nFkw8HlB7Ur49NythX50LwACnXua8p//OcgB
u7nw7HxsuebzQ88BQDp/ZynlaCvWlOVb2QBspFncE1pZd/Y7zzU7npQzbZBWLYbkpDq5PuWmnRE/
IImmJhSqWz4OTSV8zfjBbRPZ1pIpEhsT5h6Zum82xhhts82y6y6M6GMwYrOzyNhWCyVg+dCkjiun
FPmPs2apg8vbTtPY0OKIuIUh4C7Z6hf1E9rH7GChU44IOTpRMpd9/e8HYTpgiavvjjtpnzpcyf8L
35pufbq2W9XS9AAvmeggtBGOekv/KFJYhnW+9hAkThDYqh7fyqtI49PTyimodxJqhXYUmTjgJIB7
JpyqIqEguFh27M76sdN8vxz0GXrw8cmUdFf2Hbb+hUJn7YK5PjjDbJTJVw16htiy2yoEFsUg2KqO
42KLkwgqtqIJ28wKz02fJZmtaELBVC2mYMWpPFTrGAqBoWaiLqga+OhnBCENObGSSqRrdl72MP6D
yttLOIgHxCGcZX+Y07sAG+s1ZiTSegCfZgnsbZwO75/IVV2a6kJ+6jj8j5CQq53C1yaBfHmASjWI
MJV4wa0Kzqdn7lZwuALS2n0tjVD14lmVziQ/y/cAoJ5iL/gQdIDJpq7VdQGVLNzq4Pb5G+JCdE+P
BO0gBDt6r4gI/FbYN7SLECIQ+B5Gwz9jHrNu8I00J+lRKSK9PJpMsmhtGyt+/WF4XKvWmcMWsxaA
Sbo+duTn+FsrDOy7+n7gkLfoVHXP4/C0hAqYKKZAW4/06D9LtcpGl9T6HqV8q+gkFup1aJuyw9B3
kKmGPQjua8h5P58G/fy+NMGOpufA2yxngFBeCrCc3Oqi7QtZ1VulbUDWHMWiIMLPao3nTnDbKr8u
JeM41OwCI2W/2gLB11s3G0NwH38F1ot0RalI8YxRxUHqFF5AJG5gbpSe6D/UIgvbMB086CCALa2w
LCHOUNViMlRbfmUCc9/HqzmAZjyK75yO/KDwUPivcRPPbpIHNJMqWCQ/9DtT1Hk2B1PGWkC8AarA
46qQ5ILaKFQEYcyNiILyV/9nAufqRsS9LpD5pkUSjSWZNqMel7KtuSXxGPKUEKN7Vf144YbZYG1f
uiX1sJYFWD7IoE1x4anlrNn8B4PhYInCa/NMrVBJEpeUG2UHp4HfxogUeKyLDy6LDRz3sF4DVBcd
WxuohmcK5C88wbaD5rtE6h/UQ0A3Mze7ngOwmIEx/S7B4F0OZkwqFs4ONQx9IBU/JIxopZhFDqwk
BaBodV8ejAVFfWqe+HnMxZHEpcD4mFG15cMThFMMsfEbRBFk+fiXcWdw3po10IwA5N8godE1gYS1
gUo5d6WQ19P1ICX0EGZoQa/pFMwhGu00u3LleKV7Y67C5wmGquBPg5UwWO/lr8FDfZ5qExMvSFmt
KXlYtruQL9ngMQ1eiUTU/3/AgdpKpT9hkhpogU7tVDmsa3eNuyO1fcL5YOE7sOTpyxpDleRT+nx2
08ovo2kIuTCRY4A+DRbylqXdxFZkJYQevuqrliG3sDCVeZj/IdillEEcl2zhmIpPxrlJbLfzzeza
yqogtDTrKJl27aiZnjoPasoIJlOnYPNOmiKEp4IOeuKTwTUBkoYDGH4g5BkR/x6xCafLfUvJbxwS
Czx/mf3Ta2TxGC6GkVN2fR0U7YIVlosVYvGHCdBQ58gmYSMRSH/h0F/LZPbP543jJfoi50UQHAXm
u6FXhMrxMI5sKp+HUkoPvn0KTtlAU3Mt+yUyETuxUsweacjumdnG6lSyhW5940DC4QW6VZhO8r4j
VU/GAvKACBFHs3XOGzRoAKfPNFbpE7eQE6BvUKGMPnI8C/rULOZS9YFy+hknW2/3SbvIxRPKaFvP
PFLL2O7Sxvje1+lKjGLDKbVyy3E+HwELlMcji6IV24foG3Im2JHwGiwI2x6cqBH7vfEDuH0dVUd+
mRFTQl8CgbTTRXIOu4qc7BqCCHXO/+uh2WCG/Bg/VAUh/qL8UGBGRGb6a2diQqNdo/Y9xJcJU6DU
OK+k58qx0wFZ3VogTUJ77wrzJ5o5Hqb6dO19qZDzYyhul/usUCRR4P92CLdigg4fQf+ooRuA22D+
6q7e9g9zB98TYY5i8Cji1Y8u6HLCedwyAwe8CJ4n9pbZP/aUQzhVZxQIm7byLQp0RjShNcfIV/yo
cjIoSNeW+mLRFIef750ksJIkYMSNV3Wntq7/J+349sKZedl9beZMY2YUsbRzAlBx8//DgN21j3uA
6E0LFbugHN63Vz+oKlM6ns+x8yaq6A4c54C3ciCpsIDSvejr+xuuH2ZaHdtjW280pwF1PZ85dCuI
uOyrWZJoUxhJNzxvNgEAZl+LU6puVx5fI1dyrqKZkKKZSSwVcmQyn65Ff9fZ5XhcvF+DXUOAqB8w
ZDHLgvjcx0JCS1ykesSRd6EbDyxiWdOKzA1wljN7v2ewNNAmsP2dm0BsAObqpiiAcZWsmslZG+OO
S6nMLWhHjkcfNSKPH0JxsNOUQwzlFuns7UFV23MYY73lwythdV+cXWLxPdXi+dqA4O0zAzjqAvgv
B5lCItHC2ZInN0LSGf/zQ94CvGC7476zSv4d5JOY7WXv0IGT5ajhSNetA8uJsHscJNQF3X0ahvQd
Umy5fi3g9NaRrmXYyznmoW9WJOAjVTEbubKKqXOCxcomp7AfgOD/v5MwBgMsEyY87NCda3N0mS7C
2YZZShqaBUGinmXjAxbWnCkMbOZsmMqEXCtVPvjDOer1HzyxYoLAuNYkxi30SVe34aI0E49jkXIJ
N/lxaQ4V55eh91F67c38KUD6dPGe/bqBoyU70CD0WfMifADCLw9JuadCqbtQ96YgrKmECVArBtaV
B+ornZVqjSxD0wXGMDFlqI07Jje8bRnAbdOtKoVMtkR56C6hlKkv41qf/IvAG5FvQ0Q3AmvFzXVM
zw8XwDkgmJPHUWIW8VYeDSOyxwmAcSSTOTQo9ysj1B2vH50QRAGWtkY7FjBB7jwhXnm8Lg0mo3hM
DKdZIiYBkjIbxspYMfViywa9TItYaE21YjWf4Xg/EZZnXAi820GujvYgCTBoSS6QkuFV2UL0RaV/
mmnKhaX1klEgbkH7ycLEm8Dk4tplCT0l0UZF9MaLT4MuGZ1B4tIq/JK4zLZQU073YIkQORTAnn3d
/pS3cvFtJ6s9PVyOE34e9HR1VIxq38OyEflItWpEoYMI/PB2ghbn/OkjQ8szolZCItuRwP/kqnOx
tVPEsWhKe8+YNNlKmptSPniEVpKzEmWicY6TlCm3SdBsOPr3cm+GTuQTVIqLUn9OleGtRK6yOi5s
Lx+Dg9QqbbnOK4Xdl/tJ06v3q4Vnh7a8D1icwOZ3/baEAUa5aXHoT2vxTeCfEB0TXvN5swbSuVR0
AvDi9ohCvy+ezboh6HAD38/AEB+Y6ZsSZs3yrCjQuM/z/n2cfZgBt2tn4wnzfufvKzq70tlRBVdf
FBdrG5MUesrUtSlcZ0vDYJ2S/8IAAnSBftSobVFfUimcL+OFFhaMzsd8JTMIXPUECGYymPm13sis
+hN+UtuNa3X/hwDytl1ukuIbrKZRvsmLggOEYA6GaxQIlaA3FiaqwgJ/uX7rsduKMLr1r7jFv4Ze
z/KEByJbPKp9jksIDh52532ZDIgRBKJmBwukQS65t/PhqmoANPbpI+7RbQEW/X4moaGY+tEiCVVH
Jcb0V/gxYqwdj32tyXfeXSocy8mtk1ogPKkThTa0KPLA/45/h2QJeSyByn6wmrxlOpqzR339JeEX
FzZdzi3OCPKsNQoBHgRvITfvCoyKkV+ePHwPOG5/uBpMhwaEBsYfXD3vOevwitc/YZkMLA3MXIBS
CwE41eEIqigPSu51A+P5OjKoYNjbTRBIxYuB1Ht/QiWgqYRaiOHHji7Ktca6gsD+Vcjp8PonOm6f
nh/shOU7RKkrAphctGGL4x9vDkmBSXZx5DYekVf93511FWi8bQghMCjpM9b3CZAvQrQ0iw8xHkDz
hbwKGCepOXzJlXsNzl3m7Utqz446/bFN/S8lU4x96HhDW6KALzGPeo85I5RbAeP2PHQu1hDAn+9G
7LgrhCg96s5A+Llby3XOSuZN5OtJkuj2lASZtI9DYLDRd8Lv410X25rtPn0oY5ckO7VqsuBpNpaQ
PQJZD6jEbEPwdlj1Bag98vOkD/X5SehFp7dXhc7Qtoh44QQ3MVcCtrCbEQrIlSFWQSs5ot2lOr87
TokoRJxDJfgjkZZbU8i490uba2JomJYOg1JTf95Kcy4aacUq6t1g0GdOSlCBkr/xWRwO29oRrggp
gGK8U1VjVsGgOYBZfv2iHmmozJYnGYq71mCOY45Eb2u9KSyz8XxEJob70mIT43ZqSCQWMfwXDaov
OGk543zWvm6DC9idBjYYJJSVPAk/V+CvLQgyF5LWM8a4v2LOdcT2yNPaev7A76o+qfBAKW8E8xdO
sYqPn3RjZEdfxWGk+PQVLG03TCyPUXAbCcEquks50qpYzONiKYesZCriGpcpY+HTgS2zc3IEDfgn
EQz9b8c96D9I4YgLbVAiGWMYL5fCB9Hq4oRks+9DQPvbh/DqVWOolpU4RJxbbAuY/DVr0b4wmMp6
f/FutCiWB2NV2rtU3b8+K6xXKE+8h2DG9F6gq0RMfy4eIASXWhVMjjMMC8m98oak4nybG6kvx6P/
iNsHqH/GcO1l67UNAVtXB1KOMaIOiQfo4KxnS3XUvfLEExzyakKf0H2wrDQXNO3gX1lln6KiS5h+
imhtRIk82wsbSxlkMYbsyqVgLOj6QKOyPNedMhYzImYuhoLK0F5ergtf7IWRfgOZOkfCR9HlDXw4
oRKYhGkzvlN+weP+G8va4l2ymy+vSU9rQRiQxbwIB61vuDgLECTsys/cGmpTzopRN1sdQEwKwpI3
OvizB+8ITR/udxRCm0aHI05eXcm0a5ixtg7+YL8pDUSPo+GGiSZEp+fvKgRRy4QMbNnjbHUUqG4h
oOosAtsL+TrXvAdrgMgztNhyIsYpaLMJrj5NJI6X7wrbeMYrVnwEWrUt+SkH+qYxCV6Mgcr6oT7F
hfUlyVy8EejUbx8bBU71YP3XckF8S9MTZrBFJEwfn8SMg9duoVGSayewuqVaVZ6154bd2ljihcd3
isKSzJtBpFWIV44zTjoaID9OtacnQjslRleV95XQ/CZW903g/mn3O0CjnhUS+3S8vNJTMKhcqlyE
tV9U0op8suDjlgbQY6vaT0q1ztb6yXBbmQhoSf8MrttrF0Mm32tRVw8CYMkAvLtoodT5iorcgP0/
/a612aplHrLi7rXikcOyStsYVYFHDOKv0hgYxzkCQUmBeXSTuN83qU1sx2IMlCE5k/uEA6TX/o5J
JpIZirK82snE7eOaqcDSqAsS0UglY3SkhRySIllCkSTSVuVZzbf2yItLW2CtnkocwZPoWjJs5a85
G9JCqK9W/hb9w7URvoTybusgH1JTRTAAqHX4AI4516PzDGSxqyJzeN+4TRbixXi1LuuCbcfSkYyL
L2WGnBRioQ/UEocYGYRdCWVUtGBPhIZMnBHYAT+sVVjwxZO6S6ddAYAt8zn5sNJ1vNcDm6Xwo6rn
Qgw7zYy8MvGPUVGpe5TivcVg21tkuBw66q2COoQr+4ToOwwvWyUfdXFvOA2v8KPjOjz+GzjoKzh+
b71YF2WZwSucZVgVi18rDfNbWgAw3yLAYv3VwCpeD0CFLrmdiuNHvrquenAr1XJWqjgAeqAF7VTW
jSh9GqrJdAGbK22IfOp1MdVHujsikwo5Epf0bdF2W0G3cqUKXJsPNSCbatwnhqRNksC/RYq9EMgA
U7MZ/gaSglX4nErvPps6WxFoNjpInNvKtnClu1riP4ZbIaHjcTHA5ln/YbjYJ7C7NMwdCrwPT77w
wY86B0ppzcgHWZ4v4g2tmwy940A7OAbCuqSQitlav7f9tb8QTRaA/Ycffl9q+VqvyPOE7xpgtu5l
NnTP9eb49A/6EEMJFx+9C6ufYmpLIM8KcnLezcI1UvLm/9PWJa1GP6tGgBAcUq/xstcREE4iWoo5
6ttZ1eeLTOdQJ3ATdeC9/ZMq8rU2YFmG075SmIhUO6GLPkLY1VdQq+5NyvYKVv9Tg4JwwcVnKGGR
y9TQZrCbO2wx9JPp5HRnfD6EPMZzRXjo6/n3M/DxtO/yWDDmpuoiXDBYlOzIMXKZ9OGrkslhc8sx
e72TmbElajQuHEayCsXsQaVB7PsCRN0ckwsB+E3eVMx80a44aQxQAAtgz67gO5hIO3QfR+ZFn4jX
pO6HaHDeysf/743p67u9dbrf5ydTZgoNnYOzgMocv05G3lLnlGvi+MEUtxk9CUm8/4IIsy4DKQpa
xQbMXkZmuC3aN8wmqj1NLTkGWcSr8XGDLVV2mZaYIlNl+xxg4FvrsA22uvuNpd4EZpQGGQl5+E1m
L+c4GiCTmWRxEh2ZxUmkfgWArBFIh0Xb6nPc04P6bCan64wfQWel4n4q1fNtguJvHXwQ0WRNxeoU
0X8a846SG1SyHDXRVe7B+sK2Ci7jaXMER0dHVt10zZsMNCzSfne/gVl6vIVBaNPcG1eD+EdqkiZP
a0GgY4c966y/GynNCJyVkHlQZejMTtgB0QIauoLaV9MRspvPbiAKLV4L/ce42vLLRPJ4Ajrywj62
ij4xGTc+HVTE6HIOsA/xmm5+nByHLS1LSJQtOcsNScRqOUPZmPXZAxsyFTM5raeMjMFuvetCAJRh
0L0YvIM6RLe/yqaXnhxVFCiVedI4s385TtKvLksaJFbMF1YdOdP68J9OI1FqzgR4OBYVfQV6BMfG
aorxGwzbHOoYHEqwR665vnQHw0aGKmpBoYul/wHSR/A/99Wuyko7UkwszFWWTb0wlBXlxAOyfOiB
k2wPwYa70P/1lHgiekTFqEd8z0bccUa5iIxN80w+gDI5e9o5asZU9eJRbK0uAmcx6ataeRDDyRsU
iDV3RfoKy2cpqTONnIPeYKW7g9i3rGvJ3cVoZ5IUMVVU7FQD5QXkDVlOlJbuDZk8jUnXIUNyQIYW
e17HcQ1RHarwN3RpWNmB6gh1SjGbZkQ6aRbYbY4GhxmOLOWHg+WLJlFQSrWXHCCmJM0wFBndxw20
HpDkEPxgozcDDgn2vhykRGYcYwipk9Cu3hqbFEyH3wvYK/13Y0tuww8VfxL6MVg8WGp+eQspmpAG
8dghhPFUOZczb93TVnMfqF0tyU1scETmnXDg86l+5MaglUQIbTC076iA7TDDaKdNngrcvj78RNmH
+RTjvU3KXtJ6EGaMjaIdauXofYnt2iK30H+6mKqpo4ybi4otmF9tegP6LNvKX3bvyA6rrdEBkuI9
2U6o7OfN22F+/IFGbGrnKNHutHZV+VO4B179QOeEp1PvOB4ixPbFzi6+rLT/QOLb4R32P+b22JSH
fNjcQCw9Vj+yq+Hjbp/uyBKs7AFLHRRymVjO7SfO1+AgjhVONOrEAtmAw4zRIAV3CAld4XAK51Mr
7lHZtxjUb1/cVYydrDhfe5JC0wm70HUmLTFEcIEIrkCAH2kxuDBSnPZ6MhN7gBiksMFEiNqhZpvy
FZRTN4P9MQL//KuQaaaLrSFLa/ydbaETcRmcIfTmc9XrM9eNoW11tPURw6eEvBfHFD20Tz/vTnPX
puY2skikLvPgSVcZ4IiW6gxOqLLRm+mTV+WKc8ojIUPKKvVhCT/yfy7TcFa3Hc847xBuwW0V9DeN
OqwjnxalU92d5Qkm/+4UAlxTrrkX685aR2Jwn4MuVMnfFWInZD9c9E1j4/B9oQCaHNvilbjcxEg7
XNBZPIeBW+nHSqxiwPFoyM8ZQNXA3xuKSSTUdK6cmBLXHm1CqB9nSzmzIyHZ+M+3qmm00knxxBts
s1BBeRhQZfGdS/1XPf37B+zBox6hZqNLhs6iBNzv0EmZJlYhCWpK9k8nSLBgxni6YlqKpAf1fzdN
5CoyEKkolNUf2RMKiDnG8SVnhHVn0LM9fRlxhpKtl3R71JBtL2Ku5+2e98rnk4AAr/P1u/bxKtS8
7G3gEpcg4gFlmLwA+nqKHf81FvOkda48VUEzBG9aUi9jYyltqIlISXLuOer5dqoxfG3zAPsEVv5u
qhWWvdm42BjdnN7/zihp73mdg3o3aL5wGZAeW6jkTuwoaNk/IasmpLDCFCfpgYnnaJ+fwgvrHtNR
Eu3k0IBeXFbxUl19rYKZBUtK43srHhtIioZp1UHlbDfGQwChOZNr6R8AI91QLBEC7Q+iflHb5Csf
1rGdzOKtDU/PiQ1aEM1+Jd152VrjU+c5A4jdzxSqT2sgvbuUf+vwowyP22/pjlt9r1x3kfPDt6ax
PkgMXCZ0GqgZZtbFSnGcQ4I0jY8IQRKmRRRa2y7jLZVkRJg6gbVhzxtrg/Yd6vtCmWNgLZ1ph0zR
vy/17nbe6j0DIVH5fPNBaYw8Fnc/hkwKf9wa2tBolvqjeliTeP+Ev9XXC7HNDHEVJksjLpo1mkYY
zmG8m2OdmgGR+4aK7bpZa81If3S98QYsPHi/rDQsFbu9yk7FQJXaYm0MnQe/3aznw28ek1CWFpHW
I+4ZdxBRmrILZc6p9DNLpJz5fwSoUmVvkM8ZbwdOSd0hPAUpOqvW4YqCXp7Ncw1PA3rzvkTrvsVm
ribIt/BuqPpDq0x7pHMZtKYppeIp4WNiInTlHt1eEZGWJjUp1QeFSR9LPS3kMeJ8n71jJtMtzQxd
G83o/qnoS9MVjQmgqrOOfBsndGgv+9enx4n150lxuWFrKyT0FzMz/Zdc20PMxbecsmDvaglpjDjm
f+4mFPwapeB9KFjxD0CFVchePobQbrzflWjm3xjp4mwv5TKb5DDIvSvYXuCtIfjaM7Stm7ncFTly
+QXfGZIzP4wijJNgSE7eA8P2nEplxx3jETvY76e0MKMZt54AHIHRoRdPbUfD3QnyS/nS/zgNrz70
EQeFqAAbdQ9YxFHjdKc2gvp+tynJE2sRGR6bmzWVOdAhdio0Q8KZBfBYhb4CBT3eOiWve9YYCGxM
1z0nH58ePrSPSwAB/SQrGakbRpKImzOEbAmEe5IFkyRKruYvdcZEWDsUok8RtBN5jE1h5OjMepiC
vC+ZuPadWf/9o6HtGbJIYqjBBKQSib6CIz8m+PsKOOvQl9nWmCvo+hH5LD847SoZX7Xiy6oniLWT
qgU5qGWTVT9wT833zQbXP91utAKwbSWff0uGIGrTHUAiiASUkNu8FVt3lLtC/tZ+I+rjXftgvREj
9OjF29RkqXO7rkRgOSz+PGEEK0FGUnDqL3j1aQvZ5/DtEQKhCfhHlGT6cWiM411HfHEXmlAlsMOx
J7AFZRiJZczELgqBtp032Q3qKQBNP4riGps2GTiRSSOd/66eZkn5RsfniFshnYNUiYdAZn+zf0LC
ffIRBz0uGhROnMLsEm3vNVDcGZ5MkYNF+/55slHfETUYvTNo7QchBp7LsoWwTFXF0yvnX1LnNNDz
4+sAJHQjcvhiNrjOuK5kgJpA3pK2Gg42dYani+k515Iqcapka3I3bsw0kgWuDY8GhyEcBM9/9cJO
TVHbiZoa6/lgkOku7XVSzxPuYUE+LZNOojotlouuzb0yuRcmsDuA4U5ft5QAlCP6rS8j+6219boP
3x9N2tQJ2FO/rhcXtQ8IF60CVOH/E587jA5Fa8zQY/RqLxlrbXcLVYwNkOj2oA+28UzbmDE6FqvR
ZpyKjQ851LncwLCnw4blyfkpN6fSPlmJnn2pWJr2/SmaG3nUsWQEfJzO+IzjmdjFgSUM1+FybQlI
D8egnzexEG9IWMaMHZ0eP9r4I4AIh5F8lmNt94pPZzWOS0UtranDGrCXVeQmzdrdq+myrvaoZmWI
clA3oAhU9/QgdoXznmp45HKksmMCMM3Z+D0cE1/ZSiHpsU0F5HJu9YpzZ/zw1wV1cAmOqedMTu+C
gmP1MqXq2IHCwHv9KBWrg1XFMvw++/7k/WWPxOjpSCZr6kSh2YsNsXETvWb4hE5+oYXLlNMGTwWw
ROYkWoL8YiK/490aCHPT3/qA7pmE47IrXFoAnKuhsdm0YeN/+qHDr86eTPl6uQ5LwZhaDIUmQ3Wq
YCbo4GovD7jhtZca1hVceqvlXIpLgvULoWa88glQx81JG+oup3FJOfAeLO0oqg11JUe2md0hPtJH
txi/LCQwvnA7gaF6ZqMC2fMroEdagmPc06/i0cfVlLa7oUEua7T4xiwp1HdXv+3HskuAYjzAg4R4
/c53kS5co9D3G+LAFnR9trNvG5RRsC8CK3CUBWa6H75CBqC3IjL0zqIU+LchMKka3X+LcVzC96GZ
IW/hSBE5CK0HGdaEa0Q+ZZTHO9SCKW7ltE/M6SoeFtoYd3mjgyOWKD49ahU8nNdXePNzPJOp5XQ9
3kL3JBfUtH1VOfD/PLUN8mC9Zj2wmMuR+YRkzmiJPDukfO7LI1rkdB3bOjQxYf1J+s8oqtriP7KV
BNgdD72FNARz2KseK+lh0IC15QTkxGybJ8ojYzlHjO3C8y8MPcpLSk0PVEmYflk6Yuj+iV0oORrG
m7Qan3tNSdHhhdoJ8FGxutEOzuqwUGKvlVXEIc7CjI9iXwvmKLD8i03V5PruqdCuMe9Aybb2CcYs
NqJz2KELjLb2NJoHX5garMWZDLEyuLMwlKpazKH0ZRYYHnt00yqqWO9KQy2RrwZ2CJtRp/fLzvkv
iSyxTW8vD5TCxhsbNLglXa0rAZlCMf5wZ/VDqScsyJ+4WyN5MIRAJKu0Vt8cYIjPymZuvvp0N1MK
x6tfAHqj0ABcUjxJCWYbpp54PGpnI7Z/I2MefNY+3MG99HCmDbXsl2+Bh90IfigzTkxIKP9x4ZK7
snvH2LH363UzbjG3ysAz79s2inqRZo3jLnOb4Y9x6SazY6QbMHizT4JnpWUDpj4bfmfqu3d7txq5
NJUt1EzrlED47gHJLC8oAK7kXD5FDX8It8KOYFZiXdxIvqTVsQ+mt5Gucryjldzi3c6bdy527Kx8
SU0d+t8J0Sk0eKkVpi25zC5ZAnYadvoChTXGQOEn1T7spf05Q3Pu17lZmiTq9i5zS0SltgS9w9W8
od7gxKy6HnBzqn87sodtx+2lgwCX05sakPG0Ifoh32o8h0SF89o9HUPQj9WtvbxLxpgOntrBsY+Z
nUR6ZEPCnRVsxFyAaSPlWw3SuQpP8coHbVy5m1muNcBkCHNv1fjzjSAQTLlqvJOqh6ozNyVq3KNg
bslQP4TnxWsaw5J9eFE1tSIUSc4mY5XjodtXNBOlpYniZ5JwcCZp/d4FworOS7LQhLKaCCVH8YAo
jKh7fHL4xPRSpK4cMunO7ryjVvab8dMqp7yY+8syhGB2tH3LB3lPSKkGNgwLTd26BxllCbMRSrq1
sgoNHc4neFN6dqbHOwOxFIDcHAYoU8PX2GIsI6a/7TLSCpCXJIuvRPnVUAwL+k+OKBvxpnK1DxSk
LJBkYXxpvqLug2Am0RjufbSnQ6SUL9gAUQnf/NuAGjWwVr5LMBXeDFRE+MnHnVygCeVAFSuwrH/s
mCcGbS9+Kqj5whQJal8SxpCnzEHjbIMyGJ53osBaxhAKj4nCwKd1vFYtbXRO8XeFLpwNBYzFyYrs
QIVoPQ6M4LtDb/gla8KTfgbBPM5yp2cUTOXynxdTbwUgiTJIZ/ZGroeQCt8paJO8Jw5fyLuuDJlk
YQp0zVGgWuiLTRTP+pky01lJU9E7d1rmbwYSZg/cy2stNHejdRlhPLn3Pd3tUVt478gjGfhy4Cj4
w09qwl2tN967jd2p8J7okQAaoxcXXtqhnWz9C3QD/7s9N4G56VYshod1YDlst5184Of/8sja+AIf
ndoqpXcIzDGKHnddrZk+YB0Jc2Koa6DYPULVdFIim61YwIF5K1AHj3Q/fkU0my/MIMucTNobwjvD
BF3aGcJkzM1UdXQjQ/qU9WHkUBiDN5gm9AVv/ES1gvBR2GMPMznO6QSHTHP+90xnOLfp7uPhM3Ht
u8pBPwPPyqcCMCJ1XbsRn9ugTaccHq9zNlEsGPxasEg+23p07JV2U8A0HDix0L+LqYsEBAnOfbdt
DymvMRst3pQ7a2guHF8RNYUi4kQyG07FyCKfQQcGnn8tsw94X8yhYXa1GNq6CgA1oL0WyFzS2XTU
Efm0DuUr6hma8mm2vb5qPYWIkjeikYHQqfr/RFX6n07gVWSb4gAHk8FrX29pxuJBxwW/N4G1aRgz
/BvP1wpgzcr8WV90tFziTQGWE0d11migvvjtfv8zDZfR4/vxu2Z3SJaE2pjwL6akHX5/ZFP5mEJI
JZ3+f6ShurQ0frfChB2lryyBCMdjfoezhH9WI8oLbxB9QZebDtCMFo353gvu16bkpna54aaOBzwS
yJQSz0EICmThBVt5TgxSym8FziJMNTzkP1AkXapjp57RxdPtw57Rp0tO2V15c7vjjGSxv0He3YHH
x/xg68JkPnoVl4GjpULgE4bnd6XClvv1hab5np7UlARFask9+aRte+1XhuG4L0oRGkfcNDY8WKWh
xcAukb3+f3fkRBivgzJ3Mi04dFu+U7kLUOQWfYgcweQnlgvM9pgXj0xO1tYNxcC9Z2y80J3H+Xll
UIeEQXRFTR4awqYj0bnueXo9GCr/3GnJbet9asRDLzwL+v/XinoizC9woEaX0kuYeqEdyL2FY/aR
1UvGBnivyjV+OO7PkcDVYInKHSxXvuEfQ8hD+1GoAxxZQ/gwVOp1cwnNhzc5RGIufbD6oG7WdrGC
ypQv6LXXC1JEq4SoEn0biUtNmdU6LhglDdIDS726CCVMq7Tt4FIH09nnL159YfZ7lQgPk6o1PP2f
mrq2IvUyDXf/+1HkK4mfBMNbYaK+YcG7LZqfI9ID+1vffzdHDw8KzVrVCKlGIJAm6suAlPm4j1ms
dDNkVVZ1RstiHBAYVIIU2NkVizCLhlY32lRaZDZashkS9x6Sf2GDSKtbOCzyDKGHSASr7EzUFeSC
snUMKdQURWdRBHEZtJhgW4MWwwhwWszJAZw9iTco9j8sCSlIrMNbGMTgunEE50D3qzBEia8f8p6R
9bBX0GAdRzEEDnQRPFcoaJU7qDKFXMHC3oe6BsRXDWp/KxHAnpLI1voAMj7hnl7WzsN7SaEH7I0e
FCKp/Ocrx9ePNRupjg6UdxMC7fUbLwnLqgPd9CiCQNDDgsigJuquBfZVmmqH3fbc0XDS2ybLynnl
//ZbYw6kJvN244D1iknL5lkemR3ulI5u1EwFbYac89EAPrxExhoBTCg79UZyv5qed7hhSUrfLkAs
h6DFUCRi0epVg2EdEbqlHrR9ZKiLMR3AW4jMFzZWvEFztra4MkMlVhnaF0ne3tejgZI1pJV88B07
PHDZD0Q29hmCk9aoZ+gdjJ927xOdIA/7x/x4y0GOCiQBU+4LR7FKVKEeZoPjDvIvFLCZ7L98Rm4n
qK2icEteheFwN+sdR/GrRWGcJS8296kJcjyQYIXBIa5pNx/X9NKhFJUW6FDtoOsI7DZXthuxbnCb
wiBSOjB7yeHfKC/oS/MPMeLaC+2+SkE4wdYh1Gjs5l7lZPo1UGCWvoNk+iDlQEGkX8+Xj2Nkmefu
16SENjMYi3PeTEs5JnmTwGn/F5Ani/ll2zWKJ8ugvXTASovMUc3FXNSEk91buS7VFOdu4c4IdaTZ
JiO4PiwC8f2d8PgB8OAxYAjMdpeoQvnnjYBDB6VSj5WQdCfKoDS1oCa/UDpA9PVwBfW7vLDmLJK8
r4VKvxSK9m+2JEAx3lV92layHJ4tMdC8hO98V2GhYN1rU2u+mr2vpEJ3st2hxIKCOOATiRbHPEmP
242GSv0kqqpGAFOH+KQc6iBDQUOjBM/FK/EFVFJEc2wu8Jw5l+OQSlGKj3kZasyfQuH7NF49FLc9
Ui2BJR/DHKSaYukniL7jmP1+s+RX2L3Ag88jClY0CcgsCTUADy5l/aaogUpb2DGYS2mzAaTuKvSa
8toOVe1lxwUFE32inslAkKzB11S5zNdPDQZSinggKwUmacNPvVcMlN4dNQKhkR2sN+xyUpMdEJ5I
Tqj+UpSB6i1+mcv71EGMfNWP796QPROhtkANmNcs2QO9m/nm3OOFjxX03YB0Ge846PkMX6DZfxIT
KdqegyYiZtt8JJfgSU3FSrUWe3sZzgw5mypH7fN9ZvmrfReVjlN4q7/axgjg+m5hnDRX3BOMOZY2
2HFmAvIfB0lCFvTYcy4/FwCaHCHhct1KPVNXZ8MTpbVDnxI/O0tWAgZnQ4frlJWYu/lUt1iy9maO
uTGdk8MyZJYQ7S2759lQCeuca+8Z0dkk0iDh0LRrEg7aFLEv+0npnsbLPPN6/KM+B/FJvzcuLAjI
NxNq0S26IWqjEQnuRHxygxDngtlqqdMFn3wMwbSPhhkcrVByuSwr1V5ljY5et2/aqW2nlo5mSRR7
443ay26uYkkg8bEYau2eq7cAw6TNwF0HjQZEgh7io4lvLXa38wbMVNdSOVRh3kslwLVIQ2Iy4wYz
XmpvdQfdDwAE+XykyaTUHEhqwSeUa0n0p8gPnnRHMau2VEV8s1qaQ9cbQZr8QQkbQ5ZG+P67WYlp
d5vfBNZ9LfQeh8OYaKVYoPGayaSsIdIxX1vnFV+LdOmyUYTA2twbRNnS0IdWUN/ArvCatJTKSF90
rSrtCQahfQZ5iW+C4lj5fnCWIs4uBrpzoaMsiVWnty1OcqGKzqwz41nLT7PKWLP96Gg4yKJpAoi6
X6O1eTE0SzTQ6AyI8PxmVJvP1vJt56nyf1B7frCjKZebeAe38dx/lQx+o1/6OMM7by1H1mQsKruo
TpqT93VqxomtllK6yj0iMDdsLcMckMdnrf1ZPwFr3U9eWZRPUOaJUC2RJRebwAfj8NgRU762cmxK
iXribcrxjhqVcQ7QLC/Ej3wdNcxyj3s/fkWEubO3UTIPu0PirlJ1DGHucDqZmPwTMjood7+9q4le
oEUAfneAQy54qIWmwB/o6atJQo2DSJj4VySCgcUI9ZQpoLtx2FuhIJRqwAq5X2wULcrNk6EoYHpM
37tqmxGs52XWOPVJpcnsGwbPXnl8zQmmw1PDB9Lmbyza3ftJQoPv5B5h3PZgVef7KWem/xBX86yd
z1isjGagx58I39thoGEVB+CpZgiPSAqRMmZld1+7FI0TQ895Mt1EnEbxbCDsTyHFDVXPajKmgZfV
9urt8tfmC0rASXJmgNm23/POrqxzBPjJyJK7ci79zQjCthmrXrkr70a4+Ai1gzVqYcFf18f+HsJ2
bo1i+DenNSapf/upIflJ6uwg5UI9+b1qK2jr1UIiFJIvpp+apD0VQD5f9QaBfBL+53VLGRfkQWLt
Hy6R3Hp2BFJkNbvtOH40t20xNSm7Yo/Za1lXsbNMY6KV2XhPb79bPB2lksDH2gk9DZ+/BS+yeFmh
Ti9l3dXbrI0ZiYy6ZhvrIG9lUL5fJ6hQVchZonDuGJcq+tOY6AufTllURdKJEUSbGm+8GK1sOZxC
jIm+48L/Pt6LlErk8Q7FzaZ7buBVAmC+2AD3Hk28ullIFJIBqoLgwKkHQnn5V6gIHJwHU3xxLP7l
aQTFE+0zsPGYVKLEJjJk6sLhUTMgdBgbUes/a080uT6hp+Eeaw9MRieJVUJaIrg2z9Afbk3jPMDQ
8toAN1ONbbvhkiTfDskVk6MwQJlYLW1o/w0XCaJBQY0PbncTXZr/T/MXNug2vmVVn9OV/5BEazfw
bwNxlEBTF8lDVqNT7Gz434afQ4g2Yb4c2ksaYtUMZihzrOXe+IvGycVX1EYl6eClPHd+NHwwu7aN
91XomuBk5D5Mww+0S3PnscvRhuQ08daWuSjPVBHQXVwfeMyzbGV0x8V+Hfv73falfCkMWtIZdrKM
MHDX9+st+cBI9cb0t3oe7+cMNOtS0DJshlQwx9KMmu8XQ6h0TCb9MYHnc4RdJ16+BdWHhorHIm3t
yg8FGFJEgbHI9bc3pnR141NoduNcbYnYSzn98NxCtYTT0ytE1zCYmDVtlJgCm6OEgLq2Me0YwZQ2
//xZ36hbYnFEPM0CaY9d5VCM5unG3heA+4pmZHRQFqXsu34z7W8wuo+vAnzuJvPAl64r9e5vbVNP
/dz0z7hpZtt18P5+xx0XkJ8vLFlvBqEKaB3Y75qQ/tvfi7AcPlJYN9Ai9kC64kYxRdxS22bJixWB
/AFvUmlWspWpUtEywMzdxoApThBp0V6GI1AhTm8VQ8eFxTfiOHYjvfOTEGsFjDNK/mzHMdVcIwjv
maI1fkfblc1BNnshzzDVBTYueLZNHVkcH7bQR7YH+krLR3H0MBoHH4q72pxFb21hXKjDlAcuX1xo
AJJfrLxQpxd9f75Pec9qegAqg6K7OKgd1gr8G+HgwqvLV5H58rdizt7JdguNyi3bINQ8t3I9dZw7
4abG95zPN34N3ZDrYFLSJxuyjFA8nJ3LjdVkbE7JZFjPMhiiczhJ+NoVBoY1lJQJGHDMouwTAqfi
6P0nT7yGjiewd+Zv1OjVGCW+F1xcxDGZjeGspeBmykavlQtCc5VnPEKaSNAN1qhtfuyIh0PjjFU9
p05P96F9YQZP5LXubXtlQvFpV6wpxYQZPyayW5slKz1fkYPnWJraS6of8FoHUmCZEXlsckH4TEyq
GT3sbP2lvJYG2bFbzL/m4jtpFn4t1Vs+6bQygSrSKaE0X2RCWy0mWxzs4+CmJdMW4nWEalyyqEbg
u2aUNO18UI0drsrChkKs47/S1t3K8rdCofp3PFeIpDUumlvaLhnGtWR+weF5ughJ7c4/Unx4mFMh
Js1AjYcOni0SVEvQuzmDLOcwU72EzBRRNm4VrI6rpa8SB/uJnbvOn8oZ5RQHOIaDnQ954pwmc8CF
U0a7H7ifGmvRTIMb58C3fUfrEefhOapMKXE6eyAr4hOQn05blRzautuyCPxkPRuzlSf0JWnJAeQO
czvsdek4SIGst6fa6HdUqRMiqJCF0paaztPJZO9x9a2d9PzFieKavkDjDcaQH59w6arlFrPA4cEB
iN+zigK67tN9dTqXPS7vVnpE6KN8E71qWnHW2ayqBwp+ShiwPeFgp+E3Tc+F742Igfb9JKqeqLDu
98r9WK7zzSk1WGCt5znluM46Qc99gAf8f1PNlLbDAVPmdWfOx2ZiImEYjkpHHbQ861Sc9ksIkwOW
VqGlLylFNzR/ISkJOcbeFPsxQl7NGH+kLO9at3FZ50v7vogFhs/4BFN0YeRR50gs2I5YGPogTpi5
0PZHfYLk215TcKNOJPc0xgJYzOgU+e/48bgwFah4WssNglsv3LJ6qKryoKKK3C/MzbEMUkCbhp53
ljAhfGJm7HoU2UJBrJsNVHMfNgjpwPNELxUaxsvLz9vHNhqCOxBth7xuKFZhnWrTuJHbfGIJfIEK
O9JryAVDiLPmSpFZ7Uk2BPsAdQKZIJHk5A026NER06XcHuK4dCptoBhC4f4wPXGgxgaP7aDh1r0s
iGoSOUTrYAJVh6ulFctAN2iNXbFx5nS9SErvhHAUF4U0yGUqA2MwKubIVNzwzmavfzGWBvJ1z1ow
s46UVKPWsMMH+2+50GYIl8syDHjBII0R8QEZBoIQAGS/BJjRgCqdGacgew6HvglZtrqlgm38YdIV
Vc6424eEExHeUsgDWpYdjG63vPGQdl2Q+wohkbWYUjYY/d9NtdPoXx3sS5aWX8/TIJKBrObvRZH1
KD/PaoqNLRIT7q+b1SkQHfE4b6nch53olI4pf6toHcElMQ7ngaiH7pLiL1BQ7tVnTa8TYhAWz0X7
jHdjHD5cCbIEizFNhPtEDWfQqDStk6vB5KIKb1g70H6h56xUkSkHZNXCNM3ymbLwHyT8NqDKKxOz
CzF7gwI8UYlY3pUqyk/A/cCLsiQYEM8OgjW9uhJm8Bf/cWxs0J4ZYB9XWY0Avi+FO9g2u8kUcqW7
8LK5WSEJNj5fzSX0JzVu4uF8yeb0F4Zd223YxOitKrG4PaANsNeyqewZGORGSpumT0AplU2e0hG9
YDU7ZSjA+FcfCJVDYZBoiu4U1zHniQvZd7+MgTNjxt4A09f87gwmenfrdjJD+bm4gFE77Sy5PfQs
iBGmGFgYt5tB355vnnUFHz25YOTIcXOVM75glhEyYdXCl8i69m+WIsjIo3e84fMlDnJMx6y+d4ZC
l+p8zmFD5fw1OM2T6Z8c/YMwbByusgok0ko/Cgh/yE/Q27JjAjfmfR6zK+r5F3vQctU2vWEXYoeV
hR6YoWPaCl5xXdHREHfYVw7XpooczeAzxF4koKIVm9mOieHlpFQ8mqQjdd4cEe2OUsKcjLpFigbk
GKsL6JTkuqs5lwNQ+1dQ7xzB4vRCF+WXeDn6aF0KwrFt7CnZSwugG6xFJLbNXaPoLM6e4Dg30/l6
Zpo5ZykE/uiGsNP2/9oASKrIa/jUWP5mB366q+tTZiN5d/xAqDAxG22a33jagCDnWx/5LvSlw2en
36APEIGfkdYGMDDAS3rCkUXs8hoItxkcmuMk0B7TCwo/wALpTnswetkoPnjw4i6D1Ccd3FyssKD3
W7yT+DQb4AufeKKZAZxGWDiY0JvKRMTwSUZzevln1eEAb7QeQRENSXwExfs/5AhnJ1l8MCxgolf4
2r/Jc9Jbuj26aXjzDuWrdFqaSU1YsTDyGEujj3Jum7BnVF7+85eQSD0pa1l9bPXigtLFT17pc4q9
KqfSp6+ual7gdPMKE4SxpO9WDFPEJK6kiIJjwAYCewH1FpsT+cZKoYJ9HsUgfrIT1aVn4Li5R/s8
68whUQuDw/g/1CPA0p7vSFFn9zzcHY3akPI6eBnvQIdv60XdYiiyU4Idfr5vnGKTFnoWHrGLXPow
jnO7oBJKMcYrtGFGJ0eWAoses1F0l3bNqZAJyEuFmVbWscC6oPQrJfEQDwa4heg7DKFerwLwgg60
8AUcYVE7gQE4IPxAb20WndfTY3EJS3YGC8eoQQpRQf79m0A7NZw1b9JxHimzxlanNoz7L1Lg/pzj
h0mzBH67QDENyuvjYruGwG+pE/bglncAb/H7Zj6gok5RVdLuH3j7owtR+VafRuxQZkr6aXQ/3mPX
FdV22iSPIRQEbOIcLM70i3Uj85avKqKH+zsASN/j9Miy97amw3DGCVVvhNLdVSCJrSoIijfuHNnq
qtlhxJEO+GaIbaHX9Ttr2eEvr8pgR0f9vLGBeUtdTJKbfkSTxcn3eOqlBqZ+WiricwA32UFGuol5
Fv7KQ5HLB36FAMrTjqJvS8L+1BIHHV7jpV8NPy4Zj6Tugh4vtKNw0n2vkGLWbWyu17trdfx+oKm4
XNibc0+S5UM9eSNGh6iVL7Ipa31e44A38tvzQTBczFY4DMa0Hau5H4pPYvRAOyG/lflJEMdkyFFq
eHnQonIDLbSdkdRAd6VQe0rGMZmpwY61mu2amqqnwYDSNDi57oO6zzfFVMkZnbvXUoCzvM0N9cFE
e1wffFarxTPos1/db3rNmggj6qXEmZBwR0F/fRbUgqhpn4VRFAKbX8an93QuUxJgmWFMgjlSoecS
0nBjBfibikPfdSDRF9KnN9wSD36qeSTGKTd3HonyEi17ZP/aaoovnaWtgdTr/eNd1Pm9E9l29hYN
VHmxyMbTUOLiyeoWVv7pkvd3WQJyyiPv3N/2PGn0m/ZtRCql/aM6A1KzABdl1dI71B/qq3q/fRdp
LPWl/Hy/v394J6M4siD8Tv+4tgXIRc7R72TYSv6ixmAgOAzN3AobvjH6ef0+RDcPptLI+DQzUXq7
LUINwmBW/ojGYBq/Igt2EuuMjr4h98EGGV8oi3JQ36ugwDWXRGvaxEgK8vOmE+QntBtx+AAqNx9v
wOScemd+qFFMqWvWOVFdxJA7mq6+37uWNvsdvy4N9MxYBAOrp/smDjJte9MiPfZSYL2zXHMhGAkW
jkhy12cpCweIgLtvEn15Z4KEmSNApwYjk6HDdH7XeO68oGW5ytvsvrnvkaPUkIyKn+KmGNXF1Suy
QTTqCboDuRRXUUQ5bBdmdII/2SiS+IXEumF02XNHRc+xr29gkqIcDm2Mh8jGICsdSjkJMAapTPx4
Epu1aHiQslmC522b4rflwHyNA73vamBCyJzGNR971orReimJCT/6qHJc5o6fMZLzperA9I3KyT5G
2nURTrDvCZLeQkqNCZ2ZVb7xdopUhyITz5pfD/cWLpFO2xzSuMIgKABTREjdJZPS+Zgb/Bivj627
rAJ81buX0Qwp6Hn5NLcmDOpqcq1XFtbX/4k7044jwblBdn8sUPb++oxbBjUO/81xhiVl/SFbfd/t
0aMdXtWeMJ22ol/L5ebh4oaAYn69JPJwMWDoCL5SaSNHLD92lzv2kiWzV0oMEzRkG376UzIYs9//
XqJTx/siEPiU/b/a+r97BpPN6rbaRvNQj2qFtDMgGjdjwZS31iVBLvy3t9PBNOBa9dpxETuFczeW
QkD4tNSnB17lD/LL/L34jxe3/Aj2gYVDGUfoiXaSCXxqy76h5C43NFWQd7KCcEPgh+BOlKbp3c1Z
s9v0smXtibtrB4rhryxGKFdiCR19VqROwlAtP0NRQtdF4tD9kxhZFrkjV9Ds8K84lrG7qAGdHRq6
vhiHyk7GE64oIvN3jDkgudmsk0j9Pmx6k7CiYfcSWa3oyPRnf1I/g7XjNABORwruKKSX+MOoObSH
ZxX7opkiJylGOrNB9ccxinVybHyawHkNLKXc55NCSo1qL6EXG5Iz9i9j6nNNWGJQNIT7zHkNG335
daI9UxbQjOpxau2zC+p8TTyKRL/svouOSkoodFnDOCTmCLcd/fJMhY6pit8hv540Y/pkQunh4Gym
kcgiX6DF/4qO1rd+ss1wTuHVXthkLZK5Ddj1vjCccueS1ZDJyeF3lElKGTMLzEW+AvK+upnt+84t
biGOYxZbSvBWE3TpsdrC2S7HCOgxthbsX+49WGbt3J5XcEjX+4nxg1llX+c+bUvYxQUkK0/O8HYD
Q1m9TlEU1pPp2ZfOUiIKrjsVzUQGOsOk7yszIXD94d0D7HUhpHTr1gdC1jUo7jcmvuuMHexjtmeG
dSL3YaRUcq1279CSA0VaCs+vO+Y36F05IS1mo4TsdddufO30I49Lri0oqqXpS62D7B3mZ2tHLe+V
JwnnphpRJdEVgJflkVfIhXeczhjY/93CUkbatDmTV7BM2Kplo7vaP7HAzkRv3/JffMJ53yzDoN+Q
cjSYKLOAuAFnPMxwxz6/NKm7OgqdoMynfjXg+O7nMIOVM2GTUp2y8xQR2/FIETEVQcsBpZI+JePd
antiMgYE0MgJrGOV7CxyWP54+JxUXmltbiVvzVfFtceW6u53ygD4NCP04cZ/bn/CCxd+miJbB3dy
QEqcjfa7q5/9m6cZJYy8hpmCSjmMz54G0qITcY+zVfOt9ayI8SEaHvuyF56DECSKeo2myh5+C878
dR1LEMF85IEubUAovVvP62pWbaeUdTjEgClBspp9Ls4+NQnW86+9I9HXh6F2dRd/gkCE/tx003Z0
07r/7HGtxViQ21pAzbjfhZdL5sacwEJeknZv2HtrGqO3RV1c54eqr2UgzUUBXo+OAQyfIhMjuThP
ul4EVmfHVP+yIBajXV8PeQO00pmahouWACZ8V04q9S/bGkYvHs4rGxHJYu2iolB3Ui5vmgRuoX0K
NelSfftsx8dlzrJx3jZquA/12yyYa5C3dw7gvPpC2YW2CH9oSWWE9bGhl9DxK+q6XB37k2lkD+gX
siUj9u7A5rRAlvx/hCmmyBFcT5RwXotZWjnwLd3/r/k+VMkPNA+Y0XfCSnsi9YfF0RpFGx4hnnV9
+KV+AozMDVgmZ/cH7whu+5KiuCE7Xqr+SZnhK15L810LpsPVxcZmCev5L4PEQ2tb3ARmvl0/lXZb
3WRitvjXP93zxY9X/ibrml+LgpCmIwzk7R35ws+BN8cdRu1X3SJy+WfSrll2JCewCPJapowdspYY
yIp2gTGYdOa16IuzFGZQwDWaOHCCZkxpwPyAI+BUUfkcmnNErKw0vdgTZ+4xHTUrgupWxzAyAJkw
Oe7/p0kuU1NhLYuMYZJFmqCnX6pqKEdi13nYvJ9g+vfBLpFSrSWGTPf1irwe/Ffe1BdW8eWKVNQp
SbeMct/zHMJnhn6KoxzCxlXIoY2Iwvo54fNBOD12VGakEgY64xushHxvLiCHLlfpjkEp8qg5vjY0
yuqZdG2/hrlIHU8m88YE6a6Q5FDDUXdAjnmVrUVo9N77P8FSoh2buJ8IGTKZcVqJ3SJn4R60RaRl
zqZYnae18yysadfSdsloDwXwwvxMjSEI8bhf2XVglPaUpR6zCQxwVDGjwGd92sxucBKiyLEY+NQI
PtMZ8N6NXN67OCDa+0H5V+NBCepXnFRnnPbFT475SkhFcxM2QroVhkAnxAw9vUe9kKoLO+aO9Lon
E9J+sDkgbyApxTatWHlVJ3IjEgDlT5a98bLM/qUJWo/NFUelVlVltxLnQFRTU2FWHNtRMRM0lYXA
vXGww8ExYKTWEoAdeHUDbsR7EDOc3sjVNy9DZYW0ZM0cxByS2zG66YvglpJnsSibzNMIcVi+NN/n
ghd9mq0GnBP5JiU687UWNsWmVkpJPEMocbLBGpZ401/881ci+WODZblWpcJ83MbF/GBMDw7W/SHG
LrBGawBXfAQWx/6CgA/W2oJe6ylOfQ4tlabJjAeWvdx6ROmLcZW4BqlUpIdKKElaXSnNRIqtFT1E
C9gPM+GVgYoh6SV7YKAIUN8WKb81MC6nxn3uVB5yEsmJW1QRwi0v9syJLSi0gQZjMAOhGGlhZBA6
ugJhd96bGzIgDDaQRl7bI2CqozdJCCpelogfBwQ8C25o3F+nYO8Y1Ns8Mgj0wpZ76Joc0J12ax4k
tXb7xKtg1Mw5WVOZKAAl+CxS9FY0xvAYyb5r1IIcUIEytWkTRzuPceb59nIL/VWwQ3/qZEU+vpMl
pVmK9L1Jqm5gL9YYFIEerL9nE2CwlrZICfcPFv14hHN0WdIhYTMJ9O5hwe6IC4MFzdoq9XLCcQqh
A8ioZQdBwB3++Z8oJxKafD3GZFBokYp1LBruyJdPhwpQVg63mNrtaCl4P1F84uk+oqKS0pBZ6+6N
ukF7X87eG0MOWiZT/A7h2qEYqWKM0Cm8sn59uiR8P621KSX5ml0abruuwOr10MidqlM7tmK1nQ6j
zwp0UO6dcfoYKHvPusACw+SVA8M4z/kIVEpmkUfYBrHQesJIC0HNoXCZ/YQ5k+WJTdm+Sco6mixl
9ApopqZnm1gQWtbraFzZrAkURaMYqxt8m9/FwIkbT8dewHEPp2VmrbS82VMgvanqtgUB4XxIj0Gi
cjQwT3MCiPbePmiC0yFkAg9iMMYlLoTA97rN8MssU5NPxu9zNlnyo5o9nOqzWp+s5r9mc0UnR9wy
pDpY5gOMDy5sFOBg4xxTnYynBsOW1VgHhE4tV9xY+6b5kD0RtfUhzFoJtsbLFktCfvLYSR5bz9cA
3l/tbnvlsyZhlyLh4WdjsOwcqELXek4Du/Khp2talHzGSm0qBsfi3Ymu3gls5kIZxuKP2NsOVnCn
IGhPde0u0qd74PXV+0PfdQmT3iHLKW6xgfVvwFWPNBwPXaRl4lbHBcmhBKVawfZgH5mKRai0t/HM
aumQa6rrDKIovc4IizA9dABb7rjNHGPzJcl5x11b4UIQa7FU7exTZsi4bi+Eo6vUaJra33YRRpxr
BDtXW7ptGHG339XMaQQrN6incBTrioHfXos61UoZmLlqKKRlJwMpMq0HwymxkGiTolUZgtPtzTyG
KxC4FeGSSJuOKCu9ARf8XV+CFP9Id/2vy6hGyHoAN1yI8Q8LAdHN+bfb7Xd1wlO7kHN1VTuAhfzJ
aJeFeEdeRzzF9+d5UfyBKXA4o2czPrOTc43hMkW/kHPqyoGe8g0sJMJOjgfG8f78vbPP8lP5cJBF
QXNDvQR/NAXu247n0bCKNxk2JM4z1z1H13aOAmHU4sFXgYIT2TynG5w95dxqVtseHdhJZjIgOnMO
0dqM3tl44xa8BXT9oNO+KjfCHUF05ZEKO+Fvh/gzC+/iHrOsRruv2uKrhwkEOSZLABhjPCEiSIRb
T3eEOD8mplt4++tHNIEdyIBd1Xk1ani18L43luHZn1sD7iMz+WcuwRylAuiHcoRw4yYZwjuZRLkr
IZAz33m7g7IzF0leYKopDQoFlKXdzi0DqIPTxcECFiimEMycUw7+RuZTAG/EDPKAoH+0jh9Cp46s
v6ZcFCdWPb5+KCyzs46Z23V0kTp17zUiP1Cm2UP8HXriNu9pYQ92yhGWn3rcm47tkNHHLydqg49D
L8KDX+5UzZ9U6YiTHYiLG3O3G8lSxHx8XzxxKBAb2nMcGp2LHlW8fMKsDJ7sGkRD8MH1DofdZywP
FymfzhcvcoSlRhukWnBbcft7KsiknV0EBdodQl74cDNOa7CiaNyhkrYZgvgbN3w/ECW/1yfuvcNt
D+WZX85YuIaGxpwSyaT0xeYAJsUUDuCh6Fm8dbgUGgNCgHxFSIFFBPoIcQzQP9Cgd7ymj0lG9HFq
ObS4Ufma7zcnbksVSpyefd7oZyZFpPbEA4NCnRqsYdJ6xu1q8mRs/+o3bZdZSl3sXMGrXREAKuka
bCw3ksQHrm0UJO4JAeQqr/IRrsdORFZgE7BDNyLniKL6jI2PQdWXTFQJT3g97RCGWNjz++7rFpA5
W7gd8Qj7p2QGIjSN0Rdw/2K4fMlQxKqmtz/EuVyUB5dmoHLSEV5N8Z8pTJ1v8v5stpc//i9A93w0
GEVoEwrMmQL70cHvl2/FhvzihbpLINnDY3cNqrCBFfLqyJmrUy7wadx2XpopcGBbt2Imkh2xJPMk
WG/0Z98Hl/r6rM6oZXtaO87ramKEOkTqBNVBNXFeFHFHpoGNLxjfA92cR2UtfTprWZgfQAC5ivMz
IZD/pXtXOpjxh5z0i4OwMjBc37jS8rkplCpMCZ/Mln0h1XMmhlhELBDfPV3MhNb7tzUGyjucTJPs
d5wcp0m+wBAFcRJCXqx0/BoCYaYN9QOIRnc+3dCMEIlfCpxJN787pKgOLoXZtchBO+tXbmyWjN5x
RFPrE/Acgq0lw2utY/Qwj0n/ndyIwSYZr1cXoa+RKqJlF849VAxItLhU749nGaT4gkEGuAAddWcY
TC84R5yjNspUM3G+uHvn1Fq/rBV3eBE0166xKyCK887tbo57sxaN1KxRMIn+SRtYBjMUc0xl7JIJ
Pj4DKtIvy69OLHWExd2hEFSl98wN+OEParJ/2NeVOQQVxcLQAWfPSEhN/roHpDcBMqHTyzeipFzY
AwAxnUdc59WZAj7CoYWLz0cw+xg3oVKBGORa6Pth6i+P0GCw2lHCJf5g4+T+85qzJvBd0mcJfcC1
+c7ZZnfppiiZsM/l58JnfGoBYDudFZrO4W7Ydu0unqI3ASbCOuXKsEquoRs59QpPk0XARelAJnm+
t/09fXSudqoioUauef/VQmcVJaEqc0v8pGV9E5wnODU9Qh0240E06wO2B3pSJswqul/B3GygJlC8
WA06z3V/udoAK5JuCDfjDeYKGJlWvyCIsCIHy9Zbmooa+5mFeX8WqFiDvDogVreTENTRQPWzlhTQ
FiFGWz1t4KvSbmqVHLueoH0xIZHtbdEvMVl0RwyHoQx5YAQMjlgdpYjDZlinnoaHjhZT/iNyuL04
pqYdAWIqq74qG0mv7SxwX8wkMu93bNFWpjI3MHh6zrAqkxhz562+25IQoOLlKrmteeirNNEhpvJh
JKifBPurpMDAR+uvdOD7txaOcrc7d/oDPw6V4MWvK5+uA42M6r956m26L8AYa+qmj1dJr5sT44dK
gssOG6B+wnfQbdtLFmngU9F4Y7f6nCANBugFGzyiVL9FfVIMAB6N1ILstFSuJYxHMk0DOVYmwupL
hC0NLQZnDT9odpVnQCbabZNRa7txPWZRKzW/2k0IT2Z4rmMNWTHGYnth0s/NHeenVLje52+SLiZZ
M3e0ffsEhAuqWq9PpAXcP4cBNjkPkEXF059eGTogac4W3qTw5SP5Kg2G5eMiM7FlzxTHx9gNJR8/
e09yi4QPjFpoh6hKfFMXTauaEUsTaj66K/XczE8Gh8qskjtUiWUy3RGGUML9g3mI1KSktqykkgOw
EkW6pyG1EmChiVUvTguHSYc7WzpNxcoT2nPUIqOYwykwQnOQ8tK0hiH1x+90TKPbE9vUjYffa1kn
p0uk/erDKzHuiHq2FVslIAJneysbN7XTlKV0zHPCHH4LCguBD2BNvHG1TCd/VEF7W8y/n/s/DAro
ZGYEAGcIIF+uw3DU+2RL0n1MPbH2TGB+U4f1eyXip7cXWZ4qo7QAeSwlAl5zIEw1hKXcS7es5eEe
NPZF9XFZ7r7phoaHwc3pVaUgaSMS7zjR2DkcRcUJ9MXwauyxqsRMMMt/C7gxQXKStGcoCNUs+PSt
Y/mW6cNUwYvUT4jwgqWD6u17yfIVLTqv1PTBHvc2a7zldq8UOnRetm3yq3MOpO3rqB9YQIEti8Ru
tXOlZ/tNYvHczAWLDEVGGFMxq4KPsgPHmP11c4SEQ1kpBAMwq40gDQAsGlxSGCD8JK3ykNYGix5Z
CDb757ZB870EbmQkTlhKjSpuTeSZypme51boO+45muhpXDOBS7d3qTJlwdB1QEfCd2bFFdH50MR+
D/+mkY25xrsxVO/O34udbzG+ZZl4IS6Cur3bglOMflcyRxfdQ43jf92Xoa4fv5Zbb/BKZMkubD4L
gpJ8pDQDUmL828UKfbhSy8EmdFQkAmRT1VIN+4ENeIbUL5UY03gMnskSKZISLwIGscs851asG8fP
U7ikaeDyOrMXvYcB7LIHiiCM7EHhjOQx9UeQTqJjtcQaaPZAcpgv7PCqGBrRWaq0kkTIiqt7CKCt
imjmgKQNs0f5KMtbbpTarckfc18uKuTVQkIQaQMmlofWumy9vquwMiFJSFey4n1YnPOAFcu5+gHQ
FWtd8mZMkfYJiEremUXUIKaNM4GtPUyBLDmZ9h5P+MCtj5fHqDd89oVxl+NyjpRQ5/gDgbkr0XkI
/jj1tVgOI9raHk1E1VrxVO8pxFNIusqHNGBQ73BQdYtMJM5U3vt+ungWrGCxeaQYpHTS++sPp/HE
ebLsULP/0TB4eOPZiVVSSvW3AVKYzD36N5Yd4Sh+Rcl0ImuXN7jEpRjrbSCXeOLP7QufPBHQ+br6
LJF6E69tX1NjiNQA591rDte3z7For1SF7eqr1vcI38JfVh6PoiV2j5gSaSdOc9CD+BWVihq3Tam/
atpZV/iPdTBKDAOiZoPKeYUQ+Hqw30cS62i2pufcjvElRX9n/63Jh7nDCPX+wTA44d08OAjYUqY2
5Vk24w6ajWRcyH/6W+rDf+mj2NQlfFiT1qTy/XHvvZn8tQdWWNnrMa9FtJ9YalMEV0b1BduAQ868
R2ovUMvV74npgQlYrA9n17v5W0isrWGB3AV9DBqrolqy0ICI7zfGFLuiqAAv7s1VZJTNhwVwCyDp
sLFGw8uxHAbHAQlO8Czrgm+KlL2L5PM32Mvvg5qndbM2JPnEOy7KZEC4S0Mwja4A960mSIBg8qdh
QyWSSKYMGlJ3CR/C2RALwQoWSxhWZlG1qgoYJcBszQ+K/cwd58LLSNlFFC6JWQKiYCJhubuYPGNO
pK5Qz5RGIfnrOhF8s18mJcHV6fJVlQqiLpz60ioFOGnW0Omfvt7Dh/gNZrBkt1NEJq0ME2Ir6TQq
5JriWAVR1ctiGrOo4psqzIzEjUnyo9iZqfDS4qeS1I5XvT3zeLvgMAftQ0+mB4nN4fuVENfoeEVD
94440A6b1xNdApaohh/BwOBolJsxT8/sTmtGM3odF+pHpS+J5S5pHHFFcWVuZu+P6CCZQY6zLSvr
d1kpypDDVdsivj5j9Yk8uFCnNcNmv5zgzkVYBTM0PmiYp8CFgZGITPvjTw5U5ngFb8K+sYDCftXO
vO6NaXSdHY8IzKBniBI0xz/llGb/EkVP4SJutJXwIGlDibWtHMyiHIi69Zz5vhRVCdi1IWyIFeUQ
r865SUmA6GR6ftQqI3RqRl9JQ6UJDxmPEo9XidjpblmzAkt09BtlDv40XcEwY1mIlkiAZd+448XI
4G+5RPdPbq2lYApiA+0hgv1tt/6kQo09YFpFtzNbb2ovRsrZRgYIraFQoPYpb8DZvWOnfZzQ/H6h
Okm56h+BvTyoHtSjOHAjoXvjyxtte1bLBjiYz8dNh7/rzMcjhr8QGf59x7w1L9TfJXMNbsmeUq0l
FexoxZH/C27ZHkpahjMd1+U1tCC35zMo4TDHWKHwCM3JzpLVo2ZRTSm4CgvkCanbtvJ9oejiDt3l
vPi8LuhzF/5gSGTHyopiceC2PZ1Oy6pOsnFyjW6X09HCiPegos8tD/KSDa0J/UV0OIJLKyLJsmNY
qZydaLTaDUyE8LloZCVjbEVc2krVJCpfHU/YRZKbu2Lla/AQTcZIkuTcgZhHL+1CjQW0boLGkmSO
t7cJr+hSMJGmML8yUQWRYDM9cenIUQYIe2q9lmgWHzFIAqBgFJjBkZN5Ls/y/z9U/Lutq9SDbZXN
xYtrW1GzVQUK28MKq4u2TZsBzOVXeDgZRQnVe6xepHHpqwGOHyoC45MP3SwPZUsqX9TiNEeNXLOd
Dwyc2UUhXMNLelSxJ56d6EpiVPjPZG0GBRQi5ROp8aL1aksEf65u7djB/ptU6STLHwkuU4+RM8Es
3uFHxnxm0CTNZmwv1yX/KGJROSssBnEuhCyb2/zY//JWYJ8Y13+VG9la6R/SxJJM5fJpEZxxJa8Q
auVDLm+snvOpUOJSa2AHk+QPQQBzcvjKGKe+JIBs8bW8yqw0vVzfSNiwBMGp4KJ1SU8V/7R+u64O
x0m+qhS2xMifABsKVE3kuLeCdFmpSNsl3qp1UdmrOCAXEQLVRZotavZexOVTYA7/FkZ2YeAT9WzR
ae4r/f4+4Im2dxLuyW7ry+j6Dl2kXc/nRr97C1RV1DH/ymuAn/ksOoOBGYIx/1fWUYLEBuiB23Wd
FGK1Z0jZbtCDO1qba8URJyPLLoAYh9TaVK08JtsPIhtFb+320mPb+rX9Ox5MU59PKWi9HIIvjlgQ
Ghx7cQVbwlyEJ3JWSOZuxJG6qNvofg198dNw1wgYKpeb+fE6a3+Wf0MgKp4uHdAtvFJSLKRIHREy
tGK4EAspMKVOnhxg0yeXISU8eJB+c4eZWmcZ+VE1oBKBXQ0RUpuYHBQ45nO498XIWgUNjclTH+o3
KGS511UbqbPqee+O/vEknSbgRnSbK78kUph4ngqs93u/s20Cl7DjY2/gW32Tbba3BpjaoDkJyACv
767XCUzWuctzxZIBy8b//8dSQbm33+ZLsA16srI5K1BInIJJiB9/ZpevYcQ1HGpOs55YwjtsrC3Y
Vbsip2db+M00D5GBc1S2A8ANXaT8t22xGAVvUYI46dZQqdieQ43qLBqQcOiHSQpc3R90ohLqwlzy
a8i8c7/jTqboZl5GSiVSPEaDN7gVJhBysE3KFODInK6LLOBU87nRMx0C2b+Au2MIxu12/L6++fGt
H7dw4iJkzuj2F77vlFngqe9TEjEmYRutA4IoSJCnVUyr8PHcqvg19jCQH4ytTiZ1/rGo0MjOTsLh
xkbkkSqpzt1HX5vcAWmgyEMUlz3zfAxBAF/yuuTQhmHF5MecDGh6bjEBa+i4nP1lfFCofQ/qIIJT
6ruTV4DzZd8jLkg/+wQv60VhicE8CZSHwYHlpfeGzcLkzs8mlk9d5rDDU2xv+zl5J+Ym2draFeA1
u438U0jXTswoAoKKDrJmGVkStTvTHs2vzdSRSVXcehEs6iuZKIXDOGYF8OksMzcwjO68yNAW6HAJ
bkyd/REInz8CnNd0dGcEHWUyhXRlEMAoiNXVyZQHxM15qA0KsoI+GWI1ViegqCunS6kX4CnuS38g
PvwEhKI/h2py1piZAgHi7jMAReMper6jBLK/NcvJBUOIGHShE2uQ3JBJp77amr0KuRoc6FTXh7p6
uwW0wf6tDTCOmjlIAgBgIIRW7gth22eXLSZce2qBRrODyzYXN5yFtMOXZS/3+bCt7GE+CDWas4To
trHxP5COOUFSYQR9Puey3jVm36ZV1Y4VDpJd+MTHedYHrsHIvLmLGzDuhsMetANBCGbtNI07Ycte
sF4bZMllpTXMMRssEQeY9TCREiY2huKLMg78RDWqJEhBU73trtBGoE8bEK/v8Qj6snlagvcJ85dC
c9VqPLPK6rs1+y2pJAKLZWhOb3f3ZVD+faYIhchdhFymoICpMIkPJweHuwBv+OFOW4Hshe91Tam0
z8TqPqugK8khyt2InnAOZglA/w3t9TnCUGZxaqFHVSouBsx6XaFXM7DUbOJt8Vr3pg4U4v1p5Y1Q
ky+xf1WDQSgMZ9mkYUs/leuOGVhPsAyUnv8FWMQcQrhDwnn6/jozAw+27udTTwbL00ChI8P5JFx1
0O1hx4NawSj5gOvkypu7ocSfY2alFwnEIKo35pfuWE7AxDmo5Ijci4/LW2JxRU6MfV3EWFTESjYc
gXwvpzKJuKo2CKDgQL/l1wIlR9kx77KVcqlzD/9d+Y2asIbh/66UXzBmZTe+44R4O2BKEWVhESVv
UAyFYFumcnuGj+uHukWZWRn4sw3RpbA9qXKERA0GVBjPUPsQkmRAhF7JYN5w8PbOMfAO1Z0pFq29
TwtbbaxmCj74nM1G2blNgqz0G2o3EJ8hlNWKqzWGFywNgmSING3zkZQlex/PWVN1Kn5J6vxOxXQ4
mjW1qmNzRHJC7oLpc4xeJZfmrsn17jpdyitUKkhY0RBzsPpiKfDa6xIPFfWexThUSCLdlqegfaTh
nk5lZMYQdp64WjcB0coCeQdfn5Q+/sxOuknlTwunqX4eY4bAG+CRj52hxGfiiA0i491d4QwdRlct
8kMFa92ypwGnkXnfQ1a5PAs/KvBF8GKgHLLEIbEtxIslocBb82/BNgTCPs5Glrbb0dpQMlVZ+6jm
BUDFnDf7xdYCJow5ofiqUdglHUxrFqvvveUBc49mhXmO/JNJvpjWoBwfkKjhlzxJsQ9f4tTKgG+G
tmDxFce62u1URH8fpN9d0WV+6mBxvpktxZgiZP4FUjFCcy/Mf+swiQOxsphXoZDMQNbzu3zd9NR+
cAyrav3KsE7TzZmx3a+E4/cYY9MAGngZHIQ7KewcI4mArenvNMYPf13pjiA73aYmk/GCyO8+wncq
6Hr+5Stx0DuLknLf+SuOrBLHey2Vf6hBPQvdkpM6Uv2bOHFmelBQSDN8Qg/wLLyBvYGCXsMzSBBb
EcuoBZTqsNaWQcnMZeS6Z9IFPGLEwABK2X9CoccW1pgroTWvsUUL6ciGDDXxyJIR/AGkEYr3adND
1aPDpuO9a4M7gjqsC0IceUsUdkZZ9W2wahp8YC5ITM36WHnOMN1bA7frywCsIZD1pcRs/dW+Rj9u
wB4WPrFutsRaEzY5O9NMZbD3usexl6lWLLov59O83EDcQKnSCeOTl5eANGBc7kWucWCtb3uMHNOa
xbkpveB38PuYBUC+bov8DxxBQJGDmv8wcTdwD8qkftHNGb634AkMj89zuTVGZiRi2m/UNY9Jcvmh
Bl/Bkl7lt8mC/vrdxPhlmGdXIQjI+ynlZuUzVBn33gGbg04gmRoUU5FpPhOe9sSRyANgxCDZ79W3
59Zhdozor6tDrVeI6OpvpaMMaIJL5qEDM4AE8fpnNL3xyLh4YiY7Gbao1m6aM9+rA3GrIEYQuAJs
proxeVV4SKgK2n/QiPAt8l8XOe4cL/pIOH7w+hHhkgjGJLJLD0KMiNBsrH5tKpn9yNdP+y9fJny1
VMPY/nFu/obXHswz63VYTrQAMo9p3KQL4Rrvh2Xijf8Qw55bzOuY4joD3/7blTp3vZIB+peN3C8h
K3+DLBXWHiCY2hkR9ecBnj0lsqA5s+UJidX+Pjim2leqiK6i/wRPNosdag2wWjBm6Wr/6I7M/Efr
2Xk3p5MeuyuacBxN74M7qmqBEI1bWyXYJeal9h+dCDx0FNqMmLclZWRtYt7+kF69sX3DarldEnd/
nj5zIW8QPFCkly7R6Up772nLLmvrMMTk2hqYZtw5ui0GRdFQHU1wjZpQFHTNJdc+pMIqmEdpUF8g
Ru903m7IT/S1yqm1fEDe5SVcrvj03KKOfxSfE0iX7425VONMnGyWIs3I6lISoSE5JYPgJVAVkxV7
c9W6hnlkYm+L2xv9/HZ5IqGBdn+84KurWG+bKZvvvkNm/c+/anAS+fNNYr6XXoiChKptJIoMXLvg
OoHMHDucw/Yx77oYWkP0wrTG9aGOQmCRm6zl4Hqe6Dc0zM3bTdsW8R8rK5WDPymn97aBgJk+aw00
uRuoONYBdnlPqTBslAzGv0w0icY3TSNJeCLSKtpAt0d8JqcBYjSn7IN5O/4xRYLte/kFPj05uZqe
A+CpZ5YoR4hIcRZvPOoVKgelU282cxaa5X1z1MnLefnYIvXjxrG3qcjPEK1mQi6NFsAEaPanq83N
Hsvv+Ar1Gv81M9io9vfGWxp0vSuzEh/5JoUuKwFP6Y48HVOxuQLrYeDZ4tO4hT9GWqQvlurB5vLC
DIhsI0Azv/X1XXrBoiTIBICsMybRhWeMFE8DJBk92Zx5gaZkpAMjGWgZ7ZNbhjcMmHJ1qZptyvrU
7I474hngH+v/s4OV93/uSL/KC0f6+jhqX9qkYgWA4JqQqXLsBmlRFN79JMHybCpVYrWiaqZ+EuR0
rVT5fDlXZfKAbYihoiqlNB+xQUeCSIs4zz3t8WrpvSlKqiKie3w/326hbc19Zc551br0o2sB6tEb
e6ctDRq+wglt7qLTeaMtI+pp5SgKIFxT57NgPi1hDbHqFe9OEM4jKmIy32Y4EMPclnba6il3tjOV
BYr+vSgY01b6gbKASgYh/42KKR7Z6PCPUtT4B2Tr+Cb8FwoCuz04UWRUhfe8ZfPAHxHSP9XAS1d0
fFBNiVGhqGiNspsqB18RouGNdJYiuRqUKe5nRPsYjzhnWge/OW/cI5sB48b6Zaow0V02WvqFZ0oP
HQTQZs9WDRVUPBSuTPCeTx+RkJs0V1O14XhiB6PEB1zn5NJkuXB+pQo3WnvC3iEUEGle0MPtcDZi
d5bJ6CYmMH8GCCBHkRSU/5v1Ixh5pKsAErW10/KZBh8ycq/Y2kP1toixHmcwiaWy6ZridMAklkSE
mFsR/BoWGQ4CIsw0aEwYNZ3WzEPp0plIPh7YKxEVYPV4VcaR71u9RNPfL3tMLgnn6T/Cqt5bEpdq
5i731YuS45EMd0raMunqhzauDlD+fNHiPfi7UgC9k/Nccc140SPgdflZzP3ir46i/eiaM79qKUWd
6T3Cx5rdEkwYCRYTbG/BquhnRfFTNyZS5YpsAnQAYNwdXGs0KIjIsOn6uFTRYNniYHu+obeft4rX
8z8l4XP3H1Mv8h5r4pQC7b0CWM5oNndrLBwZb584/qiPXqT5l2fXWjLm6upvygOXHIm6i6m3HI0C
Vlr45NsCyfKDbLGjKZ31kmUq9davlskuTLePpX+LWOvEfzzvNUWxVBczBQFOfg7+BC7KXhhv1WUQ
VMrZgl/XLfxgjIcfUADoyhV1+xXqvVAlAKHYra8YCrUDNk6Dl/UHK4oY3HUV+tQ+BIxRAnpIxSu/
kZzY/yni139WJFzOd7PAfJ3jiP2W1d/JZq6VT7E/Z+pdHG7dbWnDLCgxZ3dUJNGcPErdP8VR4pV5
FL4VAdZRjjmKhhYdN5j+vRGFDb6/Kd8QwfwsFAxqJkaWhFD5AwxPwWfQj/25+nHeR+0zSK5CpUuA
rLNvLeBviBslLG5BK4Q3YAeu11QZVCOVCfjApi52Qg+WPd7ILwozAZc65+5DH2kVETIli9y8lsFU
7A5e8ZehTCTr4lDn/wypEVbyDuF/1c6CQR8Ugvm5V/PdOnsMd5t2Ha9N+q229wheYGuq6ejFVeFS
oDRszIDiJkJw9vvfqZiH73LHEYK/P5+cQIwt52e3y0mIeCeoX4VoFW49p7FlyEvZzicVl4ZB7t3Y
iJk80VFmkRdVS3fteRX18n2b4uNtMzyU1CxNTjeeMdijaDlBG4h9jAUX6HoayEIjE9+IkD4eH2Q8
kNh795/H8qNPm6M4VsMeezT/Z0wuz+W9SHGhr7+uzQrxdMeW+hl7Q/qu++YcAskAQac0OPvJwGnN
SU7iLub1e9gEAwppfqsXMMbzZGSjxgbUBJPKDRF8iewurpMlnVKrbct5NqaDl72kX0GLIaItNhhO
YXv0+uQScn/to/zcKAj5n086yMaQ74bF1vbbiOz6ylXFSDRBwcwYzmxiD43yGS6Jt3qALGmi0igq
rxpsGm/Ni7//KstGQJR3J/5aTC82DXH0YvqHuHNpz1B8KT8xTG5BtvgyOPHXxUMVJ9LmGl7edXJ9
eObgHTO9N2ZW7XdrT6ersiMTIvjvP7V7+zcd8MmNcEyktIscw3t+1eU7N1K9qkMvNpF/g6uXDstJ
HnF6ENUxDRP7ik5NNcZE/2G4iXeFMxQ5nkf2ZU0ZnOfRITSHzxwd928tOJBp7oFxX8yOk9l2bQfJ
aiWFysaiTMkghIGdtuIA+sGh7UlSoCDw8ecNxPlzmhrieb0ZXORrAwdfqNpYNvc0DLIhNP1D7QHg
xrX1qZ8lMycBMYE7aTie78uzUkrbqiQxtRPi7itIERuTL61JMQkC7znC8KK8cvtSwjG8MhdmOWDI
QVKhB7K18fzEZ+roiB4PhGmvO0QtTihk8kYJfZBKxzOwTtrCgjh1Ztg05DyVIo69HIlIjWrut8TU
D2etn0UCEHH0UvJsNQGL+MXjjf3Mq5MFXqKCckv+0AbI7xvtKZeBzRKl8y/QOe9vcdrLzoYrKdKx
/8sezPNAYaQeKFHDcjSgyT6YlCFL0s0V/mFhL3qJcqZ/sloKBFjSeJeKnraQP0YPrU2JAbMGY9EW
UUUxwDZdWqaNzVf0Q6Qy7xRWgiOu8oyo/IS6ynqul1jPZxGg+N4QP/E5TYBTNBVcI7ZenG5HSiWO
UHE1ingHXXAyxOqpICHzHqg1QdgrZIZO9Y0GsS9OrpEf+Cir1otq0LNTY0ZtIcGnZplsr2KIfK9a
23xVlg50WNwx/UEWe/mMbNLsZWeUUtmEbLbERgI9EV8zAcK7L0Xmh7c3AuXZidMxaG56UXpFzv17
TaiqvQMAq0bkrN4FGhdDo7imiW7en/DHRUz1f0cbyu/O7XRPnTmqiWkjzLwaCFLqSOGmC8TMu76/
Hf58k0srgoKT+JcECwZG9PDcqrVWQQ3WF+GbvUJx+tkPQXFD8ASLRDP59qD7+sejL8thcohcgf9O
1QhU14pnEB4xrjx5kTyKCIFefofY9VIrbn5eJq9pXbqsKk3jN6oSPoRwni6vUeleVgXuvhLqoB5M
MlWwGk+lTuUY5Cez/5WIi9cD8mHjdoIWhg653/Prp6+TOlK4FUS/Aj9kyyCEkJVL3Gf/GGsLeHB8
wKJ0/Glf/MyEhtZsmQS+GPgCix8Q87OUzLE3dCEL6owJP7JErFHrnBZ8EMafLuc3RWb8aTeYIhT8
Aom6nSANycYJ+m/oP+FoSiyBtFaaPbhe3hr1P4FXPOs9iE4PEDaK42bI00xbSaFK4yHg9+pw8OzX
t2fdBsHQ0iASW5+08nv/Wz9WqMXKgQOCsL+B7oYGCPM4XD1Zco3SCNd/U8tEgpOH3VYELy5O9CiJ
noHknYgGy81tJrtI7ljZHG4Ph8VpiPOy81kV4yzTdUI7bHj/+tDs4Drd3MQY3HVzcgIpTQMYPyKK
UMTPNOq8LjifbWiWkJgYvnPdr45cnx7DwvEETJwu7nzI4LwljQQqXIFldQANe0bcAq/Xukteltjo
y+fCUkUwJXzaFYfH9fSHcD/7x4xl6V6FNUPlblYsdqwJ7OvVL05NZO/KwwkHxvJUCiGoCI9T7PkY
I6fLYlIqZZlv4Ap90Zo0wIzhlYWLrNHZDTT/jFFmNZxEsF9zs8yd5/dUVmeRXgkgbgYJvS0u4lG7
6GFnhONShe1fZBmEhBhdfxk0DYRA9NoHcmK1keveLJTXeLDhduDxEsVVs+5dIyco53Vz8QGdRLjR
730YM59flm12FHnsnEbmBrGBWr9A3xGvamYJkHrwZ/8K+R3XbVsfI1H3lM9ckjbXftULK6gTE9Hx
gkdFS8h1EJysfcf4nua2X/d0ZQwbifOUrQaxShRbeBBo2eAarnQ1M0y+JtE3A5nlx8ukjv1jNM/h
TPFabPMwGHXjQk/USKAOdmLls1xhhkf0pf5+6O72cw7dtx3Vwr+H6tqgonCBNjxM/84mFyqS+sBF
R3G4QReesUxfy4VlEMv6AW6oVdSGqlSfTuZ8gF/no3K3R0ISt0SSeB7SVxuQq+fDgc8SskFpR0tu
JzOy+gy+DUMW1D3Xt80Q8r3Qr0LZ4Lu/I0IaxGlPoJbY0zWhdfgtJnAnd/yAXw4QUtBMJQUoEUfQ
SxjO2i3nc+iv3zHaCpMFkbNzZOOaG6u9QGq1+4ffXU4hpemW1wGdwz247KsV60iwgSEBNSCzAFr+
ZloNT/gltX6pQCKP0cCth1o/H4Wgt/hilKk26d4QH58Fw2XeuEw/7DJAI4HO1eV9uGfF4UmsvKLO
KtW8q8P3EDrhKIxBeYFSv4G2KLY1xSM+NdEdRdgSk4rNUlk2X1MlEFnujzaJbBYsizDmBy5D/qAb
GLzf640qMMZw3nKR/jZ/Xs1Yeuf0ljIyTbL3Xoi4g58NOyTJemPTaG/FzYrBGYLDuuHlozbpMDSS
YQWtReZai0GqqhP3xRj9KsiCnylrkIs6xSrCkuEuPFdacVZCib5SzMnpT6Z+F93cCi0sf5is1cV1
X0YEwz/92K6Wkb6PJxUIVK3y4qocGJQF3B3oxEfK2jDOGfasvzNNd9OveCD+L2KF1WxBk28BROWd
SeujplXejknMaUFuifcWP0rkK+NtdvnUxeUsUoqfR9F2oT5iDNFu7f7tNDK3oNFEDYKONV57QyoA
eb+4u/QcBTbf/Oc01Bvu+WDjl1FfFpzM30lo4zUKug0Or9eJ34qRoAaTREfVP/qjYfXT0eV4QkBo
OR+Lkr8HpU5MLPWv6uc9qWuMXhTi6FY+VLVp+L7z6V7FMuu/RA591pOq6Az1v3YQijpkzBYqRvF+
lscuPWF1fuP/2qawirmhdD/dtTgI2Hyts7eTwSSFTl7qq5iwt7I0mkdWj7Vx9S7Sq5hjTkgtr5tx
E471b8X0MOWwa48VBTnCx2nWVugkWbdwEE+Oobi3BJWtM6NgAiyTc0c+hE9IofLymrZ7fmLUOR1F
fcIYkn7+D1gfMOEJN3Lv1IRMBBSsnGwaf8WfVVQLFJw5wZS9rT7AwPMOozxRasO04x6/vzBxSPxV
X8fiC0KEj2wx0dxkMyiV6aGvvpdKAv4NOGkLALAomicDc5UGKzvzXU6jitcYk9eENO+UiHz5lFa6
jWcCPwrIvPoEya9WckEITzlF7DTRWbrvsffhup3HYctIdls2eak30g9tgiQRlM4yeOxyaEnGGkRp
p/ji1V72gv0I+1Ywcnj2w27q2uP48KYAeneHv06x1PgFPzJYDiHO91qNrlX2yT+5VabDpDLuxwrP
6Ej3UuBnmDm//u85uQjfaeBwtefc8klU6Lp7w06wV7exMSDyoH6ZZhFmYlo3ossII/fIVZXBuuFR
0ogI5HYwpsLKN1rWIF5F4z8ERfAHjlwbydkSxB0i192qHehs/AWadn9WoEeqik3Ji4d3+OOxi6v4
SVLr6JGznaYE607SigDvkxxTouS9cIsmRW+tsESFbsb9v7vObneBwUWPNecHtlxpqeYPSPUOv90T
STANtTMLs7pPTDbUULY85B6oAMttADEy72Apv6M016XgHTC8rKItblp8iGQGbnHFGRIGF0jfImeV
8rlyIxkHKK4iGVwRkaCPU72muRUxfG90oUfLA6yefufz2brOJ2dvYYle2u5wgXSNLtNQIZ1DumXb
JTfr0+oa33HycQArI5qaqpk2v25rZAorB3pBWvQ0GAPdkJpzNUtTzfWf6xWCmOLLLjreTGUNnBsf
i+/Y1i5WanxMwY9pLDQyCoPDnSYhETZ8Qft4QKo6731olwfqKi62WtxqVORhzDc1zwu6Vs7vc9YZ
PdpjS635Fkh0ND6OSGoyU79l/skgYrfl1njq2E3tIpimc3P7CCyrRxUVxDpv1YQeiX9DCSyPrIFj
ad83jrnQ+2C3GY9GI6s0kjO+oRtXbZcKDH5RcCPrkv00Kmy2w31Nt9XwJnVWUXbrrtLrDVobTzn4
mEIqLYh/BIO0PiOcX/u9ESXfpZHJP4U5TEOha56CKUlZMp+5hc5msxU6N/vc0H0PmWNJFfN3s0Pp
3aEFBQxvcWHww68UtACK6cSCsCWMsr8owwQc6Ne31831+90B86axzuJmdNnpMJuZoD7amnLxTiUu
QrcbsnOWmIjaKPimp4wYYC8ffMxNws+F4jD1azYxjGj+xxJA1HTgzw8wvj0ctXZlVDuaUbBxopIR
aPweIwcOrqAe1dErowRraerYXHPB+5jIi3GM2KjUJIuxTNXTg74kjslHLDdmMjC+q5fdC33HzV8r
Ei1BtJjkcHPCBysJotGB37YXhCDkXxFioDHC3dWcp1WxOMK256L38+w1QZ/6wCLgc3p3m0+mbfhZ
nlGfIpomfMyzcNsOJ8MUsp0TTDhMucp+pxXClXTELjDTsgtbaBcYSJMEBxY9cP3lKDEPzNeYanMR
YdzTSWs6GmAjBdJtnv/S4N/j5rrYw9TNL6lv7qrDzqg4RJfocYqazuSYmjkOIZmbt4GPxI7tkGsV
syyCW8d5ZXN0x315cCFYgvKQZ+LenpNsKk87GKFmDchwZMO/b6WrivGKNIbGIT+pPeMW5BMQ81zT
x3IDJ6pWUIRvQPIM304MbNx3xkGEa3OYA9p9ooIxrj8nb7ZSdj3FpwEUjMv2SCqLevuK8gVPCZIT
CDssrd4nzzi4sxYdmxZl1zNu0lyVirQADVz18fbJ3y4QucSt4UanEvhsCy1c/su4vEpA3gT+ehjD
XBUmxV7sn9j4B+EZQ0+/+aRmZxW6hgS5JbWNyf+3P9KayKjzvIqY5gVFx70FHqJ4uf2dTbB78zsL
prkY9VkGLkXs5mkSicIW5zaF4GOmG8XLvHlZcUs7i9efUYlHVwDeX/WCm7fEkuQNwUVypvr+Q5vG
sYrQxP8w2XzsjC1et2MBFy5FBIuPgSxQeh8G7v64iw++qeFNEBWAPdlpB+tjVjxDNVKHxsrzcBnc
cbGiPIc8+3QyM7MXLHqqeI/6y1DstoWAOUOkK96cc9/MuDAHrW2zs+ibYZp2GMIwMnStD+/L99AD
joy0EjNP4hFgWDjruzU8CLf98wrPWphyQnFxLiBYrHSC/taoHgPjmSezN7GpJlAMxXy1y7tbIEMH
+cl/6ftSxmqVx3u4NVAHFD9yAa+de1V/GLDlyxXVPJV9fe0SGLdW/kNVPgdd5v8blKnaCTt8XMl2
JC+Tvq7AaiOWVUTJsE4yX0CPnn70gBSZ9yIxH/rVbZyuVUMUA/dD3rXE3BKz7tXtDCzb2GFfYYWJ
DpvbUGdZo67Bs+nx03sm0i5tNEuGyvKnytze/qEbsg5tZLmMptt7s4LRJcVYPZXqqQs0fuczdzZB
JkECwaAaUb35lfAo2TGBG1Eit/I6Viykou83vx5LXnuF3U5Gi+kPbuCIjDMV3Od/oy87UiT/xf+G
8mPV6/GSxlwg8HOSlyUqgKC9nXfTIO4PIftngsWo2Tf+apHDvDQAu0WkVmq/+kQCEXvpMJEhhGAV
GZSKVhuTHT185HCHXKbHjQYPXiIcD21nUPp7tXIg+wkNYrpCgTExjLJ1Xvdp1r0ftB2wDUTl58ln
PCc2bEPg1W7O05yW78V7B7Pk9EDNqlt6GIeMmPxeR01ZMVMqV8u05X8NNyWV2FIGRO2eNxUPaavx
grihp62PxrKnyLOb6NpQoqS3acMOo06XCbtGXLzMKOsicYugWr2klFmaSeKx2y8PD1sKmfjI7hH+
obIjvtKb7DhIClQT+Es9abSaHEiXjD/8S7P2M+ymS/fIpF4bdWM6nmkEWBr14DE6OrCJ9kQagy3r
ei70llHYOfjLWinq6kB72o+Ry/WMbfye9VtL5Bi9+L/L20XXY2VYzM9fWRqMgOBKU9KcTtsEZQXj
PiBdiQt0qEqpuQ5wreIYFInAr0G6B5Ogihi87q5lsEdSuPQ/ZZkqxLL/HoGAwgYXc4xaloXcq4hU
hL5rEanvvVE5+YI+1HM0DM7+YadgwKGJX07fTjCLaolgoemSWi1o2NLFSCz2eaUZre81WhPDfAq0
QOzirq80Ov55VD0kntD7b7IThr43sAtcADnsCFcfRg3e3K1oV21werygv+8WLbPnpj0a/xmFZtWt
68vHRgD2tYt4mu5i5zK6O2Ia5xVbOmmOoDfepSShutZuyK40BZV2XtkxFyK2ExgY43c44TaVBi0C
rifYv/FQXnSbTEfiumvzVp6R33vtGQREC/PLMXP7ij2zQqun3p0DgBiiEftQvnZTBmGBiyLmXXPm
3oHa/IkRgYB/caeWAQ2ZUD7Oa2DMZoLoDTEAGfC+uBQBcX6Ks0Jh+gb8gZw1WKt19aVUxOE9k65f
r+HtVIUJJvASOtmFonr5DDwZHLA9e1aP3M+Jkj9yiL6b4QF0lBK/PVMb+5QfHVmpxiwAPwnigNAT
h6INs8ytS+iABSv27pF7L/mxjBHzo1L3g07IZtCvX48VZDjojgrowwHVhrBYcoTVcziThnGt7wuP
L1ZyEhdt3oYN6upmFlVcUY+FjmSbuCZ4FAEPIQ5YB9juO92Fm7vISYYN/Jae1D1mojDg7Ga4XxHL
PCQAkAzXTrHzydIcMlYC/HHJ+Z3LqRTjXNP4lwUyaR9jkUE3C6fUsnzjpkQaFEONV/xGWQCtZ3OI
d49c/B23Os597tzh/13NjgR32KasV3tMiziZVMh3nFVOArDNNZcLbGzF0T8SsR0YVNe/X19VhU70
UsOoNTvlkmt3iXtXkXkWZUs7PGTxmc7p2h9l2E7KN+MoCROgJ1r+ZmQqCqow+TpRxMVt4CxE1lOy
G1QE5sYdKXb4N/H3s4YYbf6NATCwFyV3hV9muN9585UBYLiXwXrA5406Vlg1Ck9OCwwktfvVykQr
tT+kp0025U58HDDcO/MYIqNNwzNEi+BT9wB/yMO3A2kDC/6qCVyI3IqMlKD4zDzFko3KIusyGm8C
dYwRja7WwL7506ZpJ9FsWln2lDxF3ini5AQ9qKee02Uep5oDgLCkGyQkieNaKBBynn/+vWoxgSqG
zCAMpe+N8qfRjjllTOQe2fByTQr85uegIwIwHeHq/8dhJrqSVQcM312E+/n0JCnQTLu35G+0zfzS
C2uO6z+taE92/QbaVctIHMkzc4FR1QdytYpST41j6aIFxmAPm9XZgku81hqr4HqHtcHiMHe4nh2k
aSHKIx2BPQ1AtGQJOEUDOZIZGYW/ie6aY/xQ5ShyALX7v/vxpiK3qEPLfwXM7/qQDnN3NmY4wVnk
zomybq4n5rCo22Il4iCRaokJ4mLez/MyT0TsqOHovxB3DJYnawNXwVlZHh20vcbjT9wFsXNnrimB
V4b8iKQ04Z8pBwqQK1Z5TV56rX/iFf19ApgZ5AhaS3ccRE24XXJwbJzY6RI0g9KB9zZwvouhJONQ
nuitR7fG3vSHPmZElotePJcB9YCyYV9+TnZpKFV2LHzcY+N0hUnla1xtGREVIV9hn7nuqxdM2z6E
J1KBjZLwAJZhcZLVFokgvKwm0RcUccjaEzdKnaAvHlVnuM82j0aWXOc5anjbcLQsM7RwZJd/ewLi
oQR2Jo/ai2D8Vvp8O2U7iB7hUX0M7+8KFMQEa2QD6ev+NPgvcFlX7PCMML3IZbrdbuxifbj3F4FQ
Gn3ypbdciFeJoTdBJZ/y4ZYGNFzAel6GOP4BWp3oDmw1begfRqInbcQ4K66zNFm8H6zo08etDmjR
23zu3gUvjjIB3ZKvFJ4p8BeAXMWKjy+axfgXBRM+149TQL8pjN+R+UEyj30/zH50rF4UYucuYUwF
+xUHf++CUbwMQkKyzBI0ytvaxFhLhxE8UtogS8yZhUKYWbBTzuelK5DSmJ8oCTk1Z04jmGoFpWaJ
Hos7iaDbTtk3yDCZo6Pk7PQ90duGlENFlbfH42+m301xqjleBGEDIZM4qVGdVvKeVW805V7HhF80
GbFuqfgsN6SyINQApNoB3weLCEo9Wl4EdS+/t9pYbu2AQ6yFeS+rLR/QF+JGI3brq9V+bF4oaqVY
0etJTGPiiJi372qQm+wJ+yYrGFmC6pP+XJJqbvzlGAmvSjNNoSEW4Q398AECt1DxPQHZ6mQi7EGw
gRoWsxbffXgrLaqjZ61ZQ6SLFD3I1Yh/XLlyH/Eol1Wf62FD+0Y6kz+LvLhNLg22aBV06CL7vYbi
KzzX7xzvWlv4YXBzCUkEMO99xnMqD0JqYrt67IStHDFRTcyWucy9Vd9ZttfzzVAA/DLBQ/2k5r9H
Nc6DEmbQcgrivzD0bFJqlb2eFl7NyLFiAMbPjhab51Vlq/UWmFDWI++98rzXyg+E6wVmB+7DPvdG
LZg1c9R6zGuHQj794uMV6JWkTl6HQDeatB+zGrDXq4DeMkpNzRtzPZbDYQEXkozD4YT5sa17t25N
Ca4NSRk3JLgutbUxW3TDgKXtrKgyjouj7JFjvNY+7NHI99L6heR49i8Ob4MSfT1Z2ZSTxUokiFsV
OdNnf5hDb65YXc60Y8P1RrW4YZEz1yCndOqP0tWn3Nce0nA6E9ZGdR1S3phOYZs3TqjEbbaxOWdx
0es3wMJ9Mu/cBHZtcShCE1YJxXwphGR0g5IXrPUUgb209+ejBlgu6btewwQlLb3IrLvhE2D7KDCW
wNqdXdiujOL+RwtwuHCBcYRXP0VMLNOBCUserPH5PyOb3Kv7s+pyDIuD7VAZTTOf6a+kusyXOd8N
u5/isVE5dOXQAguAtZD0OWFX/tOo+KTlYpyDTIww8fxpSyAsxHXnkTjWvwQtn8OEQdtSFeUlVSG6
vloyN/ouxzNP6AYZdBd5LUJFTI2a6tVEI49Q4ybkSKCv8FEj6orv8D+01BPNXWaWQGawiTkIGTDD
H51lVcntEmB0YHshTfuRBjZfSBKVk26DcsI8HL6mu4eBV+/XHl5C/3eLwtfPY+ZQrqa8wnmlq+0a
/s6tL44ivMpsOorx18k8RbcJhq5T3/iKlmbLEyNiBHQ435PMSm3Or8Hv9uVGf4R1RgZ7dSd9WRgd
AGB5MMmqGq9brVPeGalNICxaVO4avTohJ+9BA5IInw+qvEYMTeoOadf6nS9kyAbGjwsxViud2GGj
FUhGF4+uQeTWdXtgIeD0+9SXMUqX8WPx3xXc5s/Jr58uz+KVsjV33DqfrwssEGvsVucsEoLyd1WU
sAGyA47pVN0sA9lyH2eUpHS9SP9KjPV5SiVYbOmI1urmJatXd8hdwAokaU5hTptfTffmjgQMuhRl
zMLrsXS2C2nZc+QA2EJuF9cUyyzP44jZfgKSyfYKvdbAZCizqOLKeuPaAd6skibwp0BmH1nrJ4Z0
rNV+9C5QUxI6ljWv6roULkbsOpxEzZxFXezJmfSoG652Iw2NxKsFzbK4A3vbkcIdMKnzNC6eGngk
EslU+Eb3TYybFEc7XwD00rjNOt0MKFp1rig2Kl7MN2vDS/W+iungjKOGnWi6ZAHI+2gmKCCT2uBb
OrfDkjBPFMdWqA18r5VctPX00wBo3S0l6mXvTV8xz1skblJ9Oj0RRYefeCl5/QWUL1NMN1H0B2nO
3JhY+eeT2uAwyWBa5jUV5vP0yS1o/MVlIvv5B5oKk4DNPrhGV53rGA9rEWn1NnCRidJFc+HIb+5Q
DfU9Rydu2Qsq1wpv9ynCRSh+AZzIRvkFigpqYhuXKgXbzHHOHTin4msVSYr3xwBxxAM5cHfFuawS
DowUxyTxeubXnlXrz/yiI3ROHCPHh2+ugUwSINotexuHvcx/cBfY2PX4RBnbvt9WIIssvouC0qpD
WLkf9ON/RPYqY7JKXdp01rzpmmIqycyixtCbvR7Py8z9dv+1lmHZ2KjHXY509htV8NZKqNJyOxTn
ncEonX+39d8PEFDny2KuK+VmKR5sMZWP12fe3WO2g80gXu/VCc0PLV3PM7tvQDA8fqWu6nHIK53c
H9eTmAbyvN197IQCM+YJx5WapdvilLLlnFi7kv160comkKp1kakOtpEWzz9Jef9bJKnOjUBSCb4U
ATigBuGJoiEod5UZUWKxwNjFEOal+MJKKYxwiD+9QbGOEFkumze8JcVSuCpp2OiNGmB2PEJXvk8D
dgEC91ZI+Z58Gp6J1ywVebDJtVj5XmLjsd025ATkNBp//Gft96DqEe+BEAtFUUkc2Jt5d776Oqc/
jRSuS3kIWp6/ghrFn3vtTdVIlbtuWE3P+QiUKzLTAMRtmw7Go9d8cX09Ced1Ii4Fhhm20Bj4No0o
kwbdUG/RbR6Puo5ay4WG7iA3J/yOIzImkcTnOH5H7yZ//Nk2M2domvmUaBkOvoIRh9VGNp5TxjKc
yEx1Jx9H6i2UtLsLKQWVC5u6GoLQV7m/7u/RzkvdWrNY6k2nrdp6at3U4wANh36Y+MEm5gIyG5xB
ncnOpUwrhjO1ak88m+K+p+w1HKYUhK2F4aXTtZ/8lo+Cn9+NuMZDHhvUm978JMso6Jl9HZj+WVJV
KAE9EiJdlFKuo+zRi3/OEOe5PUYcAvYivdod31/lPwtdgM4EJKCVQx4KlLQ9YkLRYDDpcfXbw+Pl
0geV0b5Yj9xVYABkW3fdlncGYI7iVWHL+Ms5RkrAtZvPtm0GMs4OM/J159gVZ/qkK9xQfh1I3M4X
Qi16xGX6f3JaWc/AFhjQKp6xwa1YFMaj5eO1+/lXliTURL+YmW7OGYv7tL7mMAsH0vjkinwr51HI
1EwJ2kEFYniXXBAhtrctjCPopR7zX/g/aUTOhkPy/5kruoRMbb3+i7oA4ydbTjhse+f2hil9NUrP
/lTcZxZ1a83ZmAobcn7bJ2smuJt+SNg139LAgrglguW4vvo2saqS8LD7jjGLdR+kJxi0Txu5D1BZ
oyEXZEiZy7+YJ2W/Qp8/yAqOjoDZ7VxDuUyTDi7CrAxv4dafX730aVA+9iQe85X9JmN49mmqxk8g
vU/oEU0pZ8+EIshTP5H6OMkgJdVq2ZgT5Gr6K0k+26Os0CvaRFcjgY/plptxN4S2PNWhB5rIsFmv
rnuCiNbGdFElEH9InVrQQtfc81MFQueHwoJKv0GbMpS2VR3QzRc4/sIBZCUFyNZL+35gYROV40RM
4MO8Xk+Ma6QVCmZUK2Ru8o/9XOlIVwcdUKfiQKvvx51K0LAoSq/X5tf3WEXG1ZYhy7wd1AtYHT2X
I1jnCYIeBX4Tz8dCBkPUKKv9wKfVSP9AHTyDjtOcPnfHzDsUuSH9aN8v7juE/K1s+lYEIRx8kERj
C1aj3ENp9OGl4OLy5dsxguox/XDnaGisUNlvUU/Bf0zWLSpj4IpwApdhBoZUiC4ybEtkFhr+8yHl
dylP+Aipb9qkFs8FIyEhHGxDwI8SuKxX65Xfd9qtiKebglPOjdenkG5zJ3wV0cYJVlDdDer3FI4X
WO0+klyOrt6Mh5/U1dwkGrEJt+yZazw2F6UG2lcBxoC98fM40pcmLiajaTcSKjiRlhZEmW32THXe
FvzKiXMtyAdlqdDQMXq6ihb2wBHAsBn6ZI/eeZqExUuLllqGDdwiXTrwXRLSyacQQe3Kawwo7000
50dg2Ig42mlU4wz3VGuE6Tb5jyoKJsWpWDLTwXGg53hSlYsGVS25G3n794rV3IGrjead8NOc0bSm
oKYKDU+Wh2vfWUt1zdc+1cExg6MqtO+Tx+0kyX8Hm0owTyM/KP+3Q2Kqr2xOdb1HRKd7W9f8ZhY0
5DqLDnFS7aBxHp4KtaKQUFMt4Rvi+IT5ahoURDzJwqetWwSs0FtbL5g3Wh2X1565QxGNKPwU4aXt
aTAIWb3BiZtMEwG2dHT0l03Tc+v8WaLbaCkVKB/obVk0DVCwP+q7e7ycHaGB1NVEtCSNDVT01I1V
Oi9r+eqUyo2hbP6zLbvTaCLd3Err1iq22DpW10lObblWLUOY4IQ07LpZPUy2JYYqvpnUa1b+7IkZ
k+yowZRH5VFDIRO6LOZSQnT8EXlz9y0+gQWJIVxs0vL8BYHseD15hPVC+yiHhrHUfeltllb7w1Ko
yuH/MNnGxultQxFil3wgH1MedNGf5f1n0adZmfCwTJH9kaBRXtbxFGbrV1Y4OFWxypbMwGizjX5O
JOHsg9t6BmgRawKigj6qxGddEzUgZmF4SPzUDja5iIgYqN/6YtVdK4hFQDqA+2cNPut4U6rsR7vK
zhpWMg7yqx4X6PX1a0nF7Vk507Hy9ng0VRX9AxJex+etodsz136QjiWROHIq7WvvoBfLb3Fby0p1
0lPef+VzKm7klxojKqwPhLUR6kFpojURWlwLVt1urlyb/Zo+g9hCTFQI9BLZP9VcIi0StQ4MF1rw
YvMUYrAxAe/3lWLh3Sp6Acv9CtBGdg0vuaew8XjAEpKzItsFngm4R7LpU6yjJBLspfeRRWmaNDfk
LUb0dTRSiDo+PGN9FLmXAvM8fJ6I45iHxfrgLxUlGTmarFbBAqWq85wqB5pX0zOfTZjNJwdFt6cV
F0GHiYBquhU4TKBFXEWc0/UIjgnUJnHFLFwUWR1vnaTii9Q1pCy00VUEZxiHNIiMAUmYVzOI/f9N
U05jWnOJ8KJdedSpGkrDa8UWGyVEbVyNCpvbgQgVT2VYo2so96zFOHmlSi8LLn8IxjOjoBIOONYw
stOb2tVOln8BcZFT0Z+WfUr+gMMZ0ggN1fxIutJWFm3i4uSjUKe0pXXJs2VYKHLyMxhsZnruY1Gd
IzIHTSx1tdQ8PTPVWsyMGiPoD9a8HXeLTZiXvw2NnLjaA60QRQ2vDtus4VRd3xAD9WthwwVKjdMH
EnIY6tJiWFW6wYi4uLUDQJ7qxBSliRmn1K6tiHkkAJ59yLJUdRSd8nixVnz/2ZgxmICKCn9RDxCY
eLYdtdTRcuDwsG0clRPV8i++hMs3nYF6/5DHRS9h60KxkQeoTEEQWOi1ZHT5i7nIgxqj2IM1qZxe
1BdZv85UQtYOznJplOnw7yyiMqKtvUJJJSCQo+uVsBbeQN2WGaV58OVx2VIMjn/LXhWYjnqqxgFv
vfF9wajporQHLXthnG5ywmxKhyg9NyHcONSyzWrMWctc8HrKmDWAuNqfOBnJ+XtD/15/T3Qqqnp+
og0wj+IAiPgvB8FFN6m5+j5egHV+gAAiMD0p923wDPvzpV1Pp7fsKlcHHNvNBo92c1cQaBAG5Mze
kCWA7p8vNAcApc7jlaM224G/TxY0n+oaSkiJnAXI0/qqUpB0jqi7F+fLTm+0umgCPGfho3uNTSlX
J8JlyeSjxvY1rHwaXeQyCfYKw4UCiC2TYHF+zs61FJBAOiwaENxpKx/2SbMX0nZ8l7Zl3jldyqHH
vIHl9MDuI7y6U/cARJ1p075kfBVP0EtGgniIIqQwVeWkos+mHW4a9y/Tbebf6tc2aNX/tZLvz+RZ
1Kx6BJtRJZ5FEqUgLOhyHB167KZnltlza+Z6oRFuU2+8u0ZR1gdDvWsTNEnsrD+c2ub9X1kVJvE6
qEXxykOnhmfkvt4rZU7HGbmDuxiFunKeR/58GzrF+V+VilJ4XqzMPA90OIZd5Qnf5V2e/TjuE+Mo
NQ62WGl3rp2AUNdg/tFrvSgr1Nz/GhI84k9flg7Q/BMIDqTag0G4volI6tJBY0yJ26b2oX/9H8rz
tqiy1Z7o1qdJFBSUoPYXmGIDrI0srv5WBcbYv+MjEYZd7BLWhWtPe4ocpIeV/JqXLaIhqflaGqg/
OyGhpsvMIea1XF1Fhde0hh0NweGZTGJ2MX0zaRMu6+ZFMz16JH6fa1DZ/KSrmK6OUKFUysK+/yGQ
Fx4YANK7fQlM112NY9RkV5xA0QaqQCuvC7voQnJKh9pvmy04+Hy0sqMLEEaEKL5MSHDPKcTgUy30
LAO3hlm9sficbbHZ9yvaHZmFYNj5Kpfb4+AtlzI5nQiwQ7ioRyVLNumK503mvH1IJykJPQsWbuRo
HI3Y626VjZQ00jnqvPS8PSPEzjOpABYgykjfhfCOmqPXzsubPysTnEYGkQnJpHx2hjl30m+ropjH
BnwVDVcAjvqsEtwtotUX1onW4cwI/K0yiL0dbHXRSwmotB/W9dfT4iZZ+Ve8acat5knnEv7tg6n6
B960iJrJhMNW4dEQKGKQ1QJU44b7OiK7aOI7vbeNsiyPFxtYujYgPEp2fmgk+XZNrtPIC+pYeQcN
toiw9fECupR7GgCdFYerynD36GHayFsHUFZJyROOmXr7rPzKuuIfIrG9oGPMk4g9lX5LZMM0119Q
8VEW4mreMgnktDVpOWBfQqS2D3UjoD/qB4Wsxw11WAoFNqT+MlqGH0SUPW8baETLP3lZ1LU7DR4L
HfmQ+Wy1QcwBJTZlIibiDoI/bj6WpiSk/mz6QKRyNI7Dg0+xAaqygTaADsrntvE9VrUSRaG3DyRv
WyzG9JZkd61ktej4QSEoeLfHoNftvNp4XhSB2L9qTusuGMLqLjMVk7i5ujnMwQ0+WyNfkzlXznjM
BOGqZbbav3DLE85x8ZVntNkSkCHiEGIBNXUonyobLVCO94CxBEG9q+VRvM2HHuVi9J2RkVH32Tio
9pborzflkGK8ACvbZn6xrWNI2U7QKOfqNU3O8Uuh32dKIH/eN+jz4aUUfZZO8miZn1WZthUBAPql
Mx0t8XJ6hZVtAB7VCVg4bQno716ySp5Nd9ObPW3RxAuXfGKwuVMb492mQYCbbh6JTdvUEYsrfJUa
X7HONZ88UJLj0A2XNa/9Y1eOb52EiD2khXTFWEkg4XJbYP4e91ClGrEuwrmwWAhsWjNjPulgAoNf
IAqD2g8Jf6XAeUXlWS0B1bw860aAD1MSbkg0Kfow/KR88l2eGVK4KftkjOzRav+fPgg+HDD4dX2X
AGnhmHb/aCFxQplcQBnrxPl2ydQ6yja7jL0/KUqsMWgTfJDSzGByecAi9vthCW5dWMSXOgxmsPsD
njmsaFMaQBcgAuakdM5AvJRMasm5qIF940uWfNfpnktfEhROBUp/E7VJOZDS5pDiXsTWUL6x4KvU
mf4LbLi92yRIUkeFZ/NZWaDAI0nAPvgmFQICnwIlgs4lGlX9k5HugysI2KAKJfbXG/rkcPBn6z7P
tHBaEjYrbh4VAx0k9CK6BDrbqzp74xAvO8Cc/Jnn5deU3mmbEDQcrOwVlxejH34+AuLfQondgQb+
7fKWWWIxZMulMtkLc2kmBTDcaXpz5F91MFcONYiDp4esZkbYMFQfLGHCcv5/m3wJlzffA/JB5xxF
aRieyro1IIVX5XL2NHp0nJ/h6l9P9Q3zOu7Vub8obwYMoK42V5QTIQ3VWl2DFIYbN9YnRmztTeS2
YPS0PvaICMb6g8soZjd5XuByHKE+xIxMTmDGIIuMWJ8y5ENLZX9IyHinKqZRjOV7l2MWEa1xsHVK
kswXIaIvQE253dehVb9O6x2mvAlr+c7TEf0hELcZfAqjLRzmQRo61063NC6xuvovi0yZ2bpEGujZ
eoHU/NBgg+EDyetSTs2WBGnXSFNtwRL8yUOTstBmBUrG0A2p20m/VN3A2PtFmBJJAzvDVT1zKqw8
tpr1crlsF5qgw+5G/uYIXh5oxmP5ParnDQJmX+Go1YyJNSyINWnM9uPDzmholGg//IqTDGhnajz5
U0Tf9zzsfZwOx9ZPqWHNIlUjuxslEdGf+Y3Vb0ynp7u4Hfv3jeCoh1dkYhbgtKCznn4kWOqX/Y2e
KEWWv7j0rDd3tC1fC6d3X4DKx9KDgUGdHeLyWlF0gkj7Kqo22SROKuP/GgHf6kTM1TntNkILiG99
Aw408Dbb1drShPlyDI4yVjuJZ+C9LzaId9K7ixxQUXzCmQp3+8/UzFs4Cc0dh/JcX5Zuqs8r/JAK
hEe0VdQBB8uJ5kQBUz2z9YgZgl+PftCCzO+/s3znukSZPXbk7nJRxZ9+agnjjhp0lmwvrAIFVHHs
eiv9OFijkMgkZk6SYKoVqRQ33EjvkO2+1Z6fJ9luvSij+6q+PJbRyMEArLvF+xEACRaL/VqNhxj0
YbWiWkwAc1AioKQqiINtwtftrFLo8NolS6Fgu1tudfwQ1VQGGW345lXbu0alvty/6SC4TXM9odoi
Oc7u6qq7jhTAjFVgJAJvPTIx/32PtcqsQgh5JQvlGmY/e4d7w55FOoLnOLYlJLxRH8W8v7ZpYCwq
JT7I1+2Ruw2rWO7weiY32oLNQJnO5n9F6GL+5+lciAldA37Flben41O+OIbwhtXlnXGs5VdQjZhQ
ONYXh1RlTCD0mlqdi/uUCcE4DGQRfoCaYY5vl9ZBZpWYpVi1pHMelvP/u8w39EzDjRdoI0lVp54H
8MNKgYt0iWoRjH4BB9miHGraKsMulJdfL9rVFdnjXDmqbf7gYH6W16g2IU1VP1rE315VdvRBHHBJ
d2dHnAmmORoBWR8pkoi2PU4njrkaWuNqOkV12pY0yftnFeDDps8H18u4YeI2I4AZBIhbbEl0TTx3
odNxP5+s+z97EQfQVD4OzcxInhB5XXaqJqbFRfpENvyWIi+vx5HKaWxJTav6TWQyTgF6T+8NZaBg
2wZD2tTX/wAP0aCHaT+g9SfFsCP6crtb3EohYXtQxIKEs29yQCJOuFVfQwjPID2Eedapk53qdJaY
iPT3wr6TfDMoSEgW1KTon/CFSOZWu8Ec9CwYjYbVQBpjpP+0SXlGvkcnMtKXLBFRHCMqn1BtlP+e
MeaBvKdudrbZXNgiZGsNTSnhrYyTgDme/yvdC9Yeb5+cKjQge5ypNiR93FauWnOv4BvzfyWwvYIK
cv//FfuXGjYYai7TvYxGV37wp+zmD+iWgoVWxZSKqCnTbhCML/wxKyHUaBRntQPSiVit2b0uKjLM
8rWEDNzgmtAZs2kPOGJzpxCjd1W7i59Yt8bsm9T7JwxE0btCDb+nnGsAm1Gzq/bEQprN1UodmmPn
ahIjnrEDo5UmeA3m/lWbd97JGrZUrDIMxO13V18I9ZbDcH0BdtBq9XyNlxbmtBoa4Gv8gL80Dfxg
88fu3a3N4wQdN74S5sMcDPA/8UzH6QE7jt6bZFcr2yjuDRo22riGI2Cx4PC2LGocFm23xaRb0SHH
gdi5MmfHq1Eg5CRVUD5KivQmCMtelaWJekKNCENU+H94TkF/46uzF+mD7NlKcYnuLIgLGZwC+G3K
ZPY+QGcN95VYTEMTmuK9fid1SU4arsm/qxR24oZaa6OGB3c37X5Y2SK+Kgh1vQRh2+aLI0HY3liM
hjVdqVkPPIAuJA30us5HKK5Yi3gthe1AMqc95KHhjgmCOXF34BwagGC5nOxFd1YGSRaoLdDKG1JO
ozNQiceCkIt2wUxcWIoXgZwIQ292D2dUhEt7daNrQFQMeSZltBG56P1GOc19pcPt+d7NQgxOZtC7
KRfULzYqdWElMgDuxtNA9oGSPxpWvhfxreiOvJS9JITmZ0MfhrgzUf70FeJwS+57TnOBiPh0wAUJ
OwwvGBcHACiJKWcgxjl5B+E8dJpla3E16eI1z80030mq5AQS1KxKK9yJSx1MwIaFBryMAiIiAhC6
tE4/dTCIsCnDbpSB5F5CY2vm4M9pLfnEzSgFjE53nhZ+XrJBNGQjMSL4/ps6N7LuRw+Xryh1dJXP
wGjBBKAwBw5aiTyghZwBuw1wcOrwIn/EaJorOvja390bp+sk5JGASSWdI00t6tDu88mF+uniukyu
DuQ9AxHJTWPlktBKDMev3tVm9RUzx+/LeT/YQfmS4Lx7j6KXrTuL/9fPU9+Mw8z1sFg3567oE+9h
+NYrljxmDAiCeOjaBlbDZusXcQKADf8uIe+7Iooisdp/YzJSlQ22SUW8Wrg4Q/kwtEA7bkVihFL5
s+1l0tpaM75JIMti/iIJgTR6O/wdWL8vADM9lYy9/YWR8DFknzYGRT5suX3EdnPFTqCqcD5/QMcb
4avKiSskDmu28IbDiSh9mOvcm0VmFl2NAc0keeG6ENvO3kGdgt99JYp3D4VfX2AbAVffhFJQ335y
fPt3FaBzofNITesqDwFVPmoZPdXbI9Rs7Pp/eLKhkCz/M2khKJoQ0EIqgzosYEC2v4IjXMr8+Puz
6TUqvVLnTdMWoKZQOtiPd39Or3vQqsBZQpT4fO6mkwPjG1r/rlqTcpZbh4PKl2GU6RYlvZsRTuYx
musRwG6YaWZqCSueN+vLIj9lPRlt1SOhVPtzKujPXgbO8rIHGcwtbTN1bseRXQ7hJsyNTOHIi3Ee
NUTssvl5HWyDkkaGOb5PA567jAlgx+mgoGiwEUmnm22mcC5rpjqlFI7ukCy64a2e+Z0BFCHe1HBv
naAfh7GM81nImBT7s1fBHH7Agx1I1jgsEfhvp2e7lPzaw3sQHykWuKxPx4EUmJuk94aUr/GbsS1G
F6t3hCfkJU2ef+mrKDiFG80FeGDdAnVeQtPXVBBagDBNTy9giKMv2AGmw2r3CoBH2/Ug4ePDZnWv
6TohLZgdBijwDgrPT/h57FUJrNXux5o7YhQA8COWeQEaHu8iOs3/LMOjhGr+RmMnjjs4B9CYEeWX
SlMl++INxkM4cwcHBFhsYYKSHgT1LQVxJy+tApNPDT1fTLCS2s0PyK4r+l2KCw2rJPZVXGPA0rqM
4xuwAyUnPulmmvKooQYd0q5Ha4Njw5CCOtouXONuR0EpIJbl4kapE7K9W9qtROV5MA6UkC4AR1WQ
3Xoei1WXXG/pVWQzn9ROhpxo01kNPC4Rc+V9UaSd1mtaLAKVTnsnEO4fcCj6v2yebJoA2QaDiNzP
6/QPucv/d7Wf7Y3Sj+4LHzFl+99jIAnZJpkZimPNiOE0fuaDnZPCgovvGphlnqCyWi0n5StqqY4k
Z1gU2zirNylE8Y6g2CYvEgmzCZZNqFA5aAbwkqvoj81cMZpgf79hSuoI0acQ8e3JtJOj1UrXt9oQ
QhHSqKt2gNt2MVouemU6B3Lbp5KKXazpUsdsPe/oDf4VBZ2rrSGpG1rg8+1wZ0XhFE+TYwZOacCN
gOEdKCgmoz0e1irE87dVsBeXnPQOHE6af07hGaHw4SJmb87NKDuHhIbvnuPA98r6JWCUgDG1A0ye
8wFXh1SVg0z5OKCO3xJ7egkU96ff6Yt76iOn963e+fJcJsUBCrwVdGme3ds5S7zsLns7VWHhbb7v
EiF9nzh4fbpzcTLQ6E4lxQ6oyS1cdwGenZHw8p0AYXupP0RLWvT5sI1t0SPpK2al0JFSl760UqYx
7cH685vvGgSGFQMNh2SMulhIBvDROxhR94ddkbv6YTEXnJjMKgDB6Wj2mOAPaV7ULTiNBXU0WB5p
lwPvEua1hyhjQqRz2tLhORIJv9d7MX25WnQfRoUnQaP7QvKkufvp9KrYqS+lKsln1a5EA4B4k8FM
zTbQS334MYcCvZT3csiq3c4tDJJQqCSbTz7ZugfOIGlUtBt5SKdb6v2GpCZX3KHAKfoLsvO0NNN2
t+aP25qc39r6b+AJd2Yg2DF6vdkJxXEERp6hqDSPL6USrZWEvLx2FIYSa3Y7PqaLrnRYs0rbKHQt
uIW5d2Db4XiDPAXtrXAA24ssSlezlhcD67kiIEXXcBv/nCxzYa+aZCXsQp9rvsEbHBi2sJzArhuZ
084/oKPpE6AzLRMid6A15ZGSXeajRvdVtJrMB9bvY0BBd1yUYu8ztmavOWyntoKiHTPK8JhbV/Ua
MpUk90nFQsindNhQDFU7uz1KM4EJKQUhoGt82vp1Jxqj6mqv8ND4Tx2O6XH8kQLMhkmM4s4elikd
4DPUxLQgitVKsaVgJDj7awCTQmBM/xNr65yOzwdHyoWdeyKkddVhTtp3wb5fDTGxrCwgZQb79UHi
pt4QzDBW0RcOgRGuXMMTPj9neiC9rsfuilxffmYsspk8WB3tNblyHCTR5hfNh1MHh8fU1Zz4Wmsu
0gVRbwJLvVb7aoOYNbf/pSDnc1+6/ivrTu/CpXB/g3vF43Oy3Ph5vQmLZla9xo9L/8kiZJ4G/E44
OPfRFJRLrKXYuvTiedudRKpWMLZgc70GHZt8sbDSVvnJCBYRYbb9ob477MWsLTHFyYNiyBQ4EbP7
9yl39dGX01dmQK4DAEy6YV6AWIcm8byTFYJxGKjrqxtCSnr0wmElIYOJL38lzEZ0uZGwwoh6+7ze
hpXrjpcA6RuBQiE0/J/TvWMlK3b5/xq8TfvVGKwC4jBpgDbgja3CEbx56KYIvkQe719+P72utnmK
ze2vsAWxkONRoCOWCWziXNmx6bOXEiMoWWq0wNCYq5BBOxDSIJwgQeqlwA5fKNw2Eaa9Gv3g8YKv
FDwFkeepJXZHXnshHhv+5xDe0x+tAB0GeIttNoiTPpLaCXjOdI8gHiSfhvTRuYIt/rJeb32EbD/r
vICtDhOuR7AV4yJTObcA1TwILQ8K8l70O/861rGsNeX/PH8esh+EaShwKPqy+PCIKJu8YgZ6Cn+f
9MPAxJixWwrxr3nefhsQpdaXVIR81uuQveZ0QoARzewA7GLx7y26Ul7cyFT19x3ZwCEeUKCNkm9j
ZcnhmrzSx5gcvfLXbpaNRHD4eoSBomqoMosvTriuxsXTXwIrt/s6q3c4vj8BWPc/yjbdeYxLHgW/
aMcY9Ps3mh8tRXPtqVn/s1dHD5e64TLZwD7VEn3UpJ2Yr58w7AdwMHIo6RVly+lMjVGVAjibbQmt
NfJUlxOXQ5JPRHZrnyd5C8YQ96yuNvLQ4lD+Ip+wEpizl51VP1xARgIAM8DfV9Bv6oTI0Pkf531Z
Cal2nf/FbhhYYw1qXOncrIargC9yoNXgAsax9zxEuDlm7rJ05BThxehKx3pKvxwpUKAuEH5T0EY3
CwU9P1RtscYiMX8MApp9E91BNqfnpYym22kuEw76kezeBf4CF+4ODbuglCs8uPuv5r2Ei8kwb40p
1xrDWTfQAiQ2J3u6BzrRYkPjYcPbxUkKccxT71G+IRyDDHY+HvJ9lSP3jvatZntbg6bszU6Bdcp3
xa6KvOrcnE+OaH5QI2fyiQubwtgbzJ5MdxTY/APjWcLWiUgunSLDo1kkTtQKGXYHUT2wJ8BaHLwn
VfS93X0zCeqoc1W7GumpvUCIoxfLS5trazuKZQiWTMp3snLcHrAFWpJuzc2mNp+OQl4Lbbl9wDpn
1RZtusNy9Jn+yip139EWw3gkZsKzim11lWtXP1SkTro43Kl1RjuHH/TT36jnpp3YDuqxxS1+WT/5
mep09NfXyEwCSLbaET/mrCOUz3klBqzscOX1irqAExSVrgNrl/O9WcLglY9BNSn/NQzbNt9f6btk
fOj9tsCi0W00wpnvjjHB51uX4jo1nLe/YTlHj3KNi8VGOuGuzRgxTWUhQlVk/PIMXFNw3LgU+EmN
LkEG0uogzJMl7V+fnXuTGa9Ju6zdO0F9XpY3gqQgi/jtAAMKuwz+OEiFpq+7PkthqqM4dNo4E8s3
PRI2jLMT+uTsH1f4FWJlagiTSmj3NPLSytrGdEttxYzPrrn+S/SVU9yXlYgSlt4kgz+OHofD6J9m
hAjFYLPEla4n0SF/Bev61RKmLwAyrdE79BMuLN5ynrDEH55gDj4soce9ryzQBuvJ9fcfp/H3bpPC
rQOmkB+ngS109xsAEu++tLioWGxLTFVCBHlT9iQDidb0csNaPC91j5+4D5kkGi9CMnsi5E23U/d4
E3TLf/INb/v8w7QkfS5aD5UKY9Ii81waJNkIdLUhmWLmyOl6nPfK+qEzKI4tRnlI4nocmwUQTB4U
VWgMLvn63lFQ8gj0hfTHNCq8OfDJm/IiIk2p7hZ82mHnhHSlaiHO7uHrFnIZ9IsplIz8H4x/SwAP
X0HebmfOslyoNbny7MCf2s3fy0x9dweuDB4SZEBN0UlGQO+TR1rGllNquarZG6Ysiql3eE2P3pYk
FneJAskYfqeu9V6hsEJIWz4Lo6pbrBKp0f1YprDfwZt7t3GrD84HkbqnK3DYvrKJhaLpBwKdPWBU
gH1C/Z7QRxPz3kejfwxnP05akRKjmbSCkKqBngnj2/yEhZZWF7bGHi/DIhfwlBOSkfLVr4fac7MQ
p4DWb6/Q2xi4jC0HaUdJCIJ0Xb+HTZGcqlzPKNzWWdEN8gEPz+jgItgH7RMEF1DJYvuce7UcOc07
mWuYEzknVlCuMwDsi+pkLre+qog4Pr/g0A+i636H+TDb3q8/bYZHaAoLm8Q3vU3H8QsVHHBkopkY
Hp3L0khpKGg1ywhJyHmrbnvIecXS9MjrxNXpDqR7Egs9kl+/hJksiWprEtAP0Jc1DGh2iwNp1K/+
TeTMQT5HU8HYA2vTcvzOfHj18zQ7QLMNMtZUK/gJT7Kmdy2BM/RZGecTe78UNV9Vi+z/teJPOju8
WxCk8VO42fbSO/3q/Mi+R+zp4Vnn//jRMyNj/m+OrUFIsVQ0SmGPgwld7iryifBPGfpiGpf4ZIAV
7/4NCHtKFbYWuE8RKvBPPeaZ5dH6jJtz9WwDvtjUXLBnO4sAI2Cc/I23qgkDJPCHUSl78FO6ctKh
TURLAC5nN7vKsTrfS8dkfexHiZ6ay74sl112h3c6gATP/+3kXbzoxRv6R93KAwT4n5qdlzRhbk1M
lbVuTqpe6sJymVrYp/SDzLuCV10LRXprBGF5Kdl24yjMNl1OAPKgs42sEVbEUmUrvBhalxorZMfu
7cmKCkzKx+WwdFFskA5y/oXSruzQoAgnabVhzB0qDS3/JvhagMPAMCscx4DxcreiSCvuHaICCUbs
siGZUJcAySSde97oNh0PlG2YiVPd33arS7xtcE0g4I2SbiXEdTQ/4VPbuslE2x2Y2jfSKCGLIlsh
8/WVrA99bNcMeeUL0NMKsY+o2kXVWeNLNO17MGvEmRd4j5+v2j2lTd0313k+TnvKbHX0WGnoUoRv
06JofY7pgQMEPOY/h/846ZoDFxiBeGMl8+SVveD3N2RF3vhaKXQYSn1fibXPW4HXyWm96opweVUA
FneXQzhk3tj3o22DshNTlo2uAHVV5Mh6Es6u+uQx5J5DSAVkIM0sT0UARyFLdzB6RyS+0XdK7fOY
ChrrI17kUUWIfh6nkYC/bAP3MpTZ4vHytKjEMW1q8W1Fo66ng3Fh5xLQxPQDvv4wPNjG0/5SKboB
vGJFSrVi29iqODGZszcLJmLFh9MTWZWRcyTNUf+20s2QZroQz2B2bFyS6L+hFEIzDMSTXLe2X+hO
xnCLED/zROIn/KFsmeszEX3+3fQ9notoQTsSPbxksnSf1WGKXvNE9BoOf4ES5V7ifZRDsUaBDkmL
xS4DENaQLYsUUSXFAD3qj1az5IWj2cIk7FR2hy8UoxW0zdrygl6VG5tIUq+haQEBNPsc6z4Vw3F6
ttFfnoyjC0GI483yJI3vEjEH3Hhi8OCDaIHWxcSnCZ5nLqKYWiguXUenlWSXoaN5wOsRAOA/pGkK
/UyeEZfwzoI7VQ8Yu5Sw0Z+p+lQSpLDD+Yh4YPTafoCfavhkswu8TBXoTVaMo4kAvO1zeyhy71pU
/c2m6wNmjx8Lj8qVFQbd+4C6KS7UZONTy2x6yO57nf5eIAPEowHVNTDPMSp9tl8js1+4+zE+PA5n
uVtaVWWCgxSqHlmpDjPL3hTBRF/PhT+JYuQenTs5XnnrsaF8oItew3xGcXPHbyQ16NRM2Z7xEUDc
dkXpqNNMGAhDrTW4PK5d3ZSkZ8pM+WksdJdyz5vPGAtqoDyR+RNVtSc0yp25vgDSRIWj8klYwgxO
l/T7mFMmaXTUSFKefN6dXXPSSaq+WCMo76e/8+Nk+VDprzHauPz/Y/v1bs4QcJboMKHm+FhJsGye
V4KApGN5YSJv6nJrD49v0GPW2BFykWNBhnSw13X3Qa7bleZydvT1qRsF5uSW3R0CaNO91IqDBIbQ
q8S7ie6EH9EnPuU6OQGfQzuPZduXs6LvEKCcNGe6rheVTOxss272W54qcd2dqOm9Qak61b0rg7bW
iYdom3K4tN5Q6BrKIqALy2w8ElcYOHKpHOBgykQepyXxWPOgkO62kFSVBQlIFNj1Hiio2NQIhuuA
y4fzLl2+m/tPYum7F+fDkTEdiyDQO6frUaEc7WuIwGTuI89A6ejzCwOwAIRamsZnfsG5fgo220hp
p2LL2nV7PO1JfFfjNfCQvD3iNp3Sb1QPsmuQLa8XvuIKIdXUGuiNY/00yplmAlv0VIJGhghzyzpM
lqIl0BiSlaBEPklL3IxtV1zkaZ936W7N/wFELuWFr++mQ1obhhzfNS2yEfbSTpRcD/7/vpqn9+Xb
UcQtZoc0Y5Rle2C2SsfNOf7TdPQt91nGjkhu695V2gvQEmqq7VSXoVQcG9KCjl1YS/YGnStJeQPj
YTk++EqI90BMSImxxcwZ4UMIs2BYquA5A8IHxq9aPUa4ekcPuNdIF2I9ScbznVZ/4MAY6Gal68/N
6IjL+qeuSytB/QDbJa26jrAbr/xx8ux/LXIcUE1kFUPzwI9tMnRRX7BV+M427IVhTgyb2EySXhVQ
3Dc3Vo8Mcd7YXDtFqomz53Wnk3z9VFe8zwXVr3aOyzKB43Faf8rzmKjFeezO5zNGJxe5xUz/yZmK
T5QjNhwOS/WvjmXPt7q5Ds2ZqqIs/N2RCrsjcwDXZc67Pu/L+xeOJczBNuY68FDNf6sJf066iDN7
nom2SPD21HyYDiJBP3snuSQbGLf2wr+9vEqD+RAOxh3cAi0yNIldFdn/qhERbj+sEC7h1ZvwAJg+
4XLSEk0XAcDta1NpNwE38wNKZK9s3kXipavEoARri8NwRC77TpknLoFkniJsDDj2wtZLwa/z68AU
FbYAW8GZnVF+AKaqGvbhQdiYdOmHcFyTqF9i0zI9wWEun1yZ3/HrbC7vr8+89Uqnk38CCVEAtMj9
QBrWbNAZ6Ku6pusIssAGA9kAfAlL6rNbYBydYdkkEyciyN2z0jXtKRdCoC1jN9Ij4zHxq2xYujXb
B6CcEmJ+Fcor75VXEQjYZjxNrDWvH3AIKEpHRhRZSVGt8kedefOjUQMtLX8GlBaTZ5p1ZsgqwbKj
yvOowsP2j5ZI5yOANxwxQyqKuMh4HZCkbB0lUEbB7cpiaUC5hvxcl8ka5asLRZaIkSKAzz2jpaKY
a0t/xTNxOwMdR30kS4Ub/JCVhQU7IkHMRmielZbgkX+7HoZkIyX+GzogBNh6j5h7re+k/LdvuG0h
43nP5x+75jFHHURWWoQE14D9wpXPK2RIvAVeBwUvcC/E46Moc9gmPF8bNm1LTAt/hT7kMLX0G3W8
Pjdsx8v8qFhUxbFjdRP/hRs6jNmzNq55IapzIYQk8Q9XcDuOHLLVsfiHgOkdZ4wObR9jRYv0XYTb
ZQ0w5uVScL+bSIUxVxI3INwfPKuouT6ydNPvbdAr8QwNgjQyjkp8pDXfzvZWpcns5pBq0rwl6sOV
pzUMyD3B3VWmJ2IvrAEYA4VOVXLfq0qpVQ6ZwUUngP2RpmWKUSWoPueMAqFld7TV61nSyC0N8yYK
4PrgLHysEBzx/l7cW3alRimQ/AnNisCbq5Xx15hyepESWth4YyP4Tmu7eccDUqTLAI6aJk6F/V3p
tlXEJSiiA32Yus+ZegB3uEA25J2TFgn0rh8px0xl9lEY8X1vBf6WUljKC5Zr/I3PqieQ+Q8UA1Zu
hbOqtz09M/jyN8Ns06ltny0sHHgNX/UkfSlw3XPGZNon3RZ8XRrg70bjfhNGijJdwwixQIfNVtNf
L78UCmihnGg22DF+NBa1e+vDkEuMhffPDaaZZAL/vAA+4CNieWNVOQ24dpYs54IS6stNxve2tOJg
stAn2tyWoDJtLZrzZlQPnxSmEHlwlvihtYFPAux+NOHPreeXViNwQy9yU88XvD2rSyTaKqTTUg35
wpPJkSooH/8ZAcNvOFLgxJdVd9I565g2T7WJHHrbpr/trN3QFcsszKvCOZGsOQmGRIBJY/tiN6Zs
NcjM5/Y4qw3RkIvR52trzQLhxRSMPrQgAypO3CE/9bI+TQVSEmjF3xON1+lIl6xcTMVNhDElJBbG
VZSfYNWtstlddzA10j7eK9xggUcCYZlThxF2sOe6NXSo1UwIiMwpXXDDiVkE71OjDzzZx/2gmjiU
aEMeLxYnJlpOdm2T2sPaJiiGWD0JnyYzr/8/MBFXTukIeZE/4k+f9j2f2Nim7Oc70hfAn1Ql+uRW
iU8XJ2JVqT69KHC3PC4gq6RnCcGPsWVoQjG/M2ln6/sKDhIe/iwDI7xQMx0zP01jxRAhvWmI+ZhZ
SjllphcQrnQs4jAOPMSaNJljgoL157IWc4UVZnMqQcoZir5oKf8SAtFnpqAbUr9x1ycVA9n4R9SE
rCqNPSb/oB9R8wbId0ZEhWykn6blxsNqVAIjPUs3Wa9e012RgBqn9ryBNJBy+rQ5zGZdLxYFsJPr
pR7HQyXTnbqwA5hOcJpv2iKp3D1uZqjJGpKp0MtqsLHelmV0YbsMuDu5QnOGwGBX4WjextSulgzH
RQqsw81/gprElpFYiorChWZeWlmeLTZ4UYp99fJN4bncxsi73OqXOmCkdiPUAwY7mBY0Fo1cGXmJ
Rzk03t1aLbYAvsB0xtxtt1ChJ8rGPA/1pXyXZRrkSMMr873GuXmEmRbBKMLvX39RZfYyzogaPBrD
NNfXWqdbfSP2GZFn9axZK+PspVQhaKjqq/EpmtVpAxVEOdc3JmiX06YQSXJf6irVMvFjs7hBWT+O
kwPM+BN9gFdN/JZl+H6iruaKPcVXHGbXJzjYuzavmywLZSK390uZz1i/RMOKIZNm8qeyr3HIg+8a
T0p4p6Ak7cvuyXrCNCqXUgslo8DOcUVHRgWcZyzEYGIpgF1wXmzhAEa+BPsUzd/UnLhMhA9zOb1g
MJkAkNt8aRGvyTxmf3liNzMuwoWaOHQxqXEL/9W5zDcETnhPPjwGofLXdk307piy6gv9M8JYgvU6
rr1sfzUhqVKQ6gCqDEsQPQ3sXD3FbNy353W2zIb/vLzJ/n0DLnWNV0NSdyHbyrJCwpMu8mxNRkfz
pAJCodepbd3rJIgLPWLkZqPI+7aBtLxsw6MwS/gyQcDhCK4B+JmCtdqQ2R6lgri1pDSDhQ4Yv1tK
iIk0f5usiMo8OURJ/00L/VfAUihEtmzmlaA0GYnBFGfHKByNlovLHCTFVSO8eRwNTw/1eblKW2n8
a3lGG9lfsONAXOSXmrqVcPZk6b6iKJLsF4WL9Ajs13fzhiC1+//deGf3uyT9OLb/S0X8+3msXtxw
WsnLwXgTmSL88UgSxFftB6Ib+a8QS1oJCF9Qo0Af68eqiMNZr1dT7eFTD+3PezeVuQK+lFU2V+4I
NC1ysd+Os3nAqAicnTG7MVyM1l6hDaVtGaIs3Y6LsG+EOgOofuF0ewXQlRx4XhAszyBgY44zUu3h
MuSpud7wdYhxglvYAiaz1Fa6DGjc64CMAX3gfoQ5UULphujtHFRFjcIjXoVZgdA088XjZcdBbNCZ
FWs6WT+kkNO4lSAsk7Fs7X/wHXG/rG45GPEV6Dsda9N+xskayA/ragbUdq+HMkhBtSvQfhpIbnGR
+jpP3cdX/Zfs2QN0Hhjdsj0nqs647YLHwy8TNofcieZbz4FDYJdzH8aXd/r+Qw4s4VmVm1nQExm2
+t7QxeG8oUdx4IfoHLeZ4dZCLcDH20tb2UMQhpx583NtKi5sOCdAupn3sGayHsuy4KlWDEZSguDQ
xc4N2Jc1QA4KxGxN91Twrx6kerDM6Q7vn455ACPKiBn6b+F1W6R/Z87S6vuVyJyeyQsg4C0OaFMv
OeZTClBCvlFBCDX3iQy+e2m7wcMKmhrfo2cmJOrvrA4Vc7/kiRGBP0oFpStGcPf+4qT7aGuyGutC
3gvfXQ9gL+kPPrnmTewddPPNcrWdd4n+7710p1oIOxvjor7AcOgzu+IUhxAxo275pdXtlpHEA4v1
63mGWiCvrY+UdiZ4pN2kbu0Gv7EVAfu2eOs6rtbFr9FN4XGyjVo1vY6F48J9ZkRgrhJA44uz75XL
04aLn74mWGjBykOTaMweZe28kTLAB3TV+23j2s0w2ssKmSiXqLgoPilmR0oMBWwaQ/ATe+zpOfmH
WU/VSURc1Fn/NpFL8DX4dNlSgR4YhuoFsk0/hyYa/i7WhQnzsFsNOjz7zd9ry4Iktc/kbBtYDSm9
uqASgJsUDC8q2jxHRmLU9J4yF4nq3xnxJqz0FCumJaJV+HPkXPXRMfY6dAI8MC/Rce/RRfw8/w3r
m8CZDHNxOYjVNMWTJ1nYdpdM90aK6EAJ2gPxU7yQ/oeuyhXfHyttUMnFLBobI4L59HqTZfRW2dUz
nfAgFjbBA47iZDnGdMT/ovQGITRioYgia/tDq1dikFthtpWK+o3RBxS36TXCBuP1bX+jSpmGZE98
wACrtUhzTqUqpiJOtlKoxYJTz2yhwsWYc2desGhAY+1jr4e977KzlQWmdPMmbExO8UwGnqH/zRU9
BU0eebnq8Yp9CiEHXLb10IXOB/C++BDRfb+7s3Bvff3VIsoZvpl+2XbD0ggYviNWr17m6EPZ7Fz/
PJ5pYidoAXthxzYfNDgkji2qblgV6IS1swnyb0HJ89G0JzUXd5y3Uj0J/OMHofF5q060uhbRY6Go
0s8MEBDqDenBdrLTnXHpy6zgOZQ47qkMpd/G23vN7HMfOVMZRz77Hw35F3DZ43uHbGXVollAo2Cg
vVoA53IPry8RjZOCo35zNfjzl+nQ9cNyHdQeUlrh6VXs2MgsaXAfaeWAJn/253ZhdtVi8upCyz1a
k8q6sG4MPJQKyquZ01SSG1uvdiIe+iXHZu6Du87VMe27iUT8JVVwys+umXxXOp13SwebIFFUKGC2
A8z2ykCBPQlo+ZoBPdXJujA8iwAsMRlTbNVaOfLI8AkqNXP8Z30aeVjjenPyj0xac3dSaqU+xzAZ
si5UFyWli3P6y3/6PNcSDYSKa+LM+0qk/xzljWplMW+An7zGiowPxQ+XZFnDNJ3keelblVBwKruW
LZOf6B0s60CK4aEf/0lN8zNZoUa5EK+gNrepfY2WB+lRCGRUn1J9Pwz4FJTNrJ6svN9OMSGIPf8j
w55x3q9ietniDfIhOiz9crS1J92nZ+pKfCqZCAabj/MKY7KALIikwFfUVre5XtmWy/H22lJgw6mp
N0bhhthGMUnigH3iEyo7c5SXQJrBA7usJxKfks5+EoW94Ire0wHhQMm2RSZ+e+xu21bv7b63DxnN
xXbY/Suvm8ixc763n4397zsEkzm9JuF9K6WpQpFQdVSpDHPzUZWfoLZ5BuHh4OCJ5QvHKF1pN7Yt
D7XQtbQMhG2GCDqAt/xhDtAu4fGvJIfWCgFURb43pRlu4CzGqhqdrbOeuJRx7n0px14iRMQaJEG9
GV6EitHY5Da8hynFkAY2mBSmHtvGMq8xSxP9H+VsLWrm7UREEy266EF0ZD+GRZibcrxW5ZjHJfIG
OHrI/QDaYXMxJKZxAGc+jdHIkwQA4ZJjTXs2KMiBAl/yigdAkRm8zg24g27A3KGJfkNkGwrd9bRj
5jeim9HXOxCfW0CExm5GsXE6t82SA++Qc4wXkZRwdiqHQO+By7l/JBE3TM7ES9IJbvX8zEYtNAV6
Low/0V6N2Mpz6aLYwgieceOWerEP/L5JiOR6rB2Z0yRqOJxcQ9MW6XR6dscJ9FncXq9eQ2csd/Ff
SyUwb4U+8MQqhUPyZjc2tM5p6G0aSHm73jRguFaQxio5SmLsBRwJWZPPa/peAXPxGDCIkCgxkA2c
A+KtuJZv787dvWPArB15GZpALq3L4BkxoJJtEy/sp1uhIHd1dgQKnPhxtZL+Idu4JXWS2dvgx9YK
f1lSPV4HwCKyCudeJ47gU0BVb2PVHa1vXeOCrPFBbX+aWWnU0Kw6bL06bEttdM+wg/ua9J3ja8PT
IVGbzBROC7fNpuc8HZ+u3kBRxB9zwINgD192iKhWw1+cPlrDbSr94NRbDQsTMHXkwtMtHGNG/89o
Grs6r9Yf1+rJzf1X5Bg46YJ9D0MXuceav4LUZQ0DVPRdZE+FiV8mbMX8YDRCtupZsHH+n8R6NEZG
YPzTENHztGSPOrLKptOvfKnoOrGj19C4YbbISSP0rk9bUpgxGH5eDKOqDcOLyeWlzoz8oG7z6S5s
AOejx+azE5OFn675n6qN8A8LtqwDy2OjBJcMcC26dDq8g095w/TovE+0Vuh4yYrA+xZNnOcF6YK9
6U5sipV6pwvjbJ45X/Ya59K3xcIKQUv4grXkDTHZzznAhCHd1ESuwrUP1JUzn0jjXo78sZLuaT69
297ZrBIKA2rZtMkQe4vVKS+ISQZM3rLce/tIQAnkoP3+S9whqQi6MFBpKE/O8JlveoU6sXlXuPbl
TVyhU+CskY+fnKnuMFIUi2WeF/GmJmogZXzC6Ye117yOtzC4nr7lN+dNHo8bO2el+wPWsjHquDpa
QleEb1aE68L+vaPQkHnW6fhmJ5cXBHsRlZ06aUZLzgOL49xvNd7eJblVYSHnwJI5LQ+Xa673hzpt
cvCa2xWWDvRBvUI323DSXQeFRDpkuLbJNFtARa1pWDo1yHoCVMUhM+neU95axmTREqrk03xQUFG1
l7WQxiGDNYIvTMo1xzljReuQWjn/o1mzhVb3mbr5xPODdU8Eb3ZnsOlNJuZGPfzB/6oqc1Ff+eFM
V6EFcEzoWer2CkeW9oQOCuX52OA4M+QALJ9qI8z4YNghtHIPiboIKo1Qc5JXf0F1ezkMlTm2P1jV
ige1Z2CL5trVvab/INrkXfvHh/Drbeo1tuMopM6PhZwWzxUgQ+3FBoOlfCB3Yk4Hm9oglTWbyZX/
tLnXl5NveywcX32YOaFuYJEpvmVHWAQyiNc784D+GKzXD8I5pD+eoHuTiLAqvjSrTQELYCZxTqFI
914/5tKlCjbJ9PaWTZ2K5nCOzO8U9RaP5RukkZLc4vf6mSr/Pk8IHucgYtdjOP3YAug3o0PD0DeS
Qi5lB6Y1+w3lnvGczZIcmaFAwN0pn9KP8H3pj4SL8PRsP4rC4hC/rw8EUB/KUygo/rFVZkqD/wr6
4Zp8NN/1YyZVkJD8F+VYK/q31cBh9daei0FotwzuK71DPhtjD/jpDIiYQvjuWyI9i6UdKyBQPhzF
Gb/E3yyaEH9gReqwr+njo9jg8MYcuMulR2vZjjnYMopKj1cmFtT83Dvt7c4YqOnMOZP3mInNMo0E
QC6nh4KmCwOX3lJ+SJ/9ocRUiljCLH4VHibkqKiuDQAf3dIEKiEY/c8GAFnuEOZ+eOdKIj/sERHD
/3h0PgozcUmopzqZ5Bud3WcZfqY94MnsirOJss0eBwhQxgZBpohfuWlqGq10Z34pmQyGJvdodpAf
cQ4jlkPcRC2yfRLsPZwvEMKWcPWiOrSPnE/UPwMCdaViXL+JNTB40pbm+p76whJ4VW/hTx1N1IY1
ywoc8AKFNOgzwP69zT2xVppBc/uCr5lJB7cYdXf7K70UgFhYie4vkyOsDPHXsPiwqq7JsJPCd2gJ
7a8910TW9Aca5SVCXCJSevg4p9XeZ7AyMfNZoK8bE13hglRxxd98201589KpRSACNpm7yXTTgYB8
RWkI/6SRDJDYiKi3hWTRdUZCHbHWOeSf25SvuO81TToyyBu9GlFMbG0wBBb+rpna0HfC1UR57LhO
MXgEVxWmM1iWi3MHjii4qnei635k7bSZ2+ZLwDY/OuiFUgU6NjAZ+aYnlqiE+H8zoc91HCkb5Jc7
iUJXHcwJwki/78BxW+RSCQnziZE0OKYfo0Z28G9SUvwnPI91b2gkDCJvML3FAx9mfc1zaeEgPSiv
obOVD6vM7vSYvZpU+G9QBI2v10JLdTdBv7OGz9aQKaqICt1VKcJlqdw4JPSO7pjA+arWkiqO9Nle
D2133uBH0OSSdxCBLd+N6jkc4jXI0nd3PmzNNedUh8pup0wTy7xFMG530yTa3CGPPMe8beEjYYCW
V+qPLa6W/2kexqkMHMb2PHTxYcNE29ezXxyBULQXTekq/yo2pv8kO5Jq+EmZr+jWNymhz1mzmvFa
+F+i5d8VarWC48T1H39mcFgJH5Jp7Y3KX+yRgd6gHXOZFJRmGi6+Jmd604qDC89NlXZgsPUfA+RO
5MJ8WGCPtxGjgnrvlHw7sSIuiIu3TFt/aChb76mPeejogLcQ3gV9Kxt2BE2uOYoZpXO4dCJG60j6
FhL3fcOJ9yjAsuP4efCgKrUGWOO78dQL3V8mTUzDBKuQcYPZwIOUTwdmVkPD5XCqgjz2CT0ihkue
PqcXdfuxnfpfNgr/iLpoTLIRTisJN7J+4BAxinnECi0ULe4wfVOLKReZIZ5pnGDEmVWLbZiEQG8S
8zhz/GCC7l8va4BjIzuvql3JXUsBe0e7vqplIHfWxJ4HFQWlkON+FrmB0OyBrNBryQbRh/OLcm5E
0itEfvawlOrO+KeTiHHb8HvMfVGp2uRfFFT7Xer2p4FkmSF2qA+JWc9np/jFjlWCXIG77/DcN2mV
kA78HbQz/fsAH9QKa9jz1YdNBbXIOyCJJcQXI4OmYSceoWUyn09giRTIhkKiP7p9TcIVLbPr0acu
HuUpoGLxmnS+vb0INVyJe7/JdOVoaveW0rys5ruYQ865+CAgqy7LtPTBe6FcSGTkpjXyCZOJJ/YM
sqd79Effh2g8ZlKryzeDBmErMdEV/Gqi6tu65/03Fc8jGqJ0bqHiTOREcyfCS4O2O9q2qvnc8j2v
Lyg8QRw1Ci13VzrpK54amIQx6HIWwnY8GWq+g7tNxDnQP5tGOcjv3IUsbN4CwiGodinTsDsOcVd3
w7md0i1pfgdbbIW/DSFQWCDPT9IP8CIBPms4gWe85YV7F0eYfSqoujw4evWcGJSk8KUO2gbQuOMK
XC140xwfgaIWBaJAPeAeVFxCGz31LXgP5/9ftKw0J7QNmE/BxqPAzvot2LRk2orGlcppeA7Gc/vU
58qCCc/kFAR+OYWE/Q+UKQE25Hy9ByAxAkdclmkcHnFdPYlXHVCyn0oD68U4fv/59AzhgdlD1Xun
xzKGCzVkv1uOYVqVl5clefWDMFebFUBC52uHH9stU0U/lLuzeM+K+UkkjMufVlTsaRH2lCMF8rYg
kjmC+2jp5Uo7RicxC1zWJQoUcCo8/VEA9S/FFHoTdAQHhGOQFZzY+zhKXAu64LVBXzNyKbbfjFzf
CaO10Z2UfJEzb3xkq2M6fvudhLXoTlB9JHovDVJE5BOpfTYRsCv1WIPcReeeWR7AGtpNDgRVSKlW
aPCVFIkPBDNdy5vHispn232hxtF9XXuy82kyjP91jp3tFj+zOCnVyOxR1eK629mUeriQ8V/H6QkD
qbT8dBijo7NeS1svSi/rAsG/RnsJ63w93wRWK6hGW2qUClYpKe2Ug4RAP6u2plG85kajEPcyjDso
kHHWoaHWSZAoo9Gu8XnL6+TbIMYm+X4oX1ekEKu3xP/xzX1PaDrW1X37yY+ninM4/13qvEOV37gi
MshzTuQkfuGXBNcKdW9+qYT9CspWcs5+w+NVlvBVa4F00e1R2i5wFy0lexgT/tB2UTfrw2rZhdWc
RKImJGwpwU3HUGFT4De7snmGk1FD8H69CVgR4bTC7w/F+/k25kwiqtM7a2ja1vZrq03uAtBDKI6k
I65dSPzJ6KwGVk9zPc1hXiyJMWun2W9+RZA7pGwZWaFN1jIk3ZFFB7ErDllGav7ybPIR+yOZPLPZ
OZRz8XQOf6AMIEIyjYMC6nQ/oSvRyDh937K/TmdJASnNsqpYeZKXDsTgF/4YTJ9DqeMd2Mv4UjQS
HetzUB96rf7W/CTPtyeOm61CL/0YYZ9U/DD9yBxpCPFpHr/EU8eimxfxYEflvanitgAdXk7eCk31
5w44q8CTgAhOfzwdNnK+AjKYJJF6rVpLl6OLokKpn7gtPKm0GQ7D/Cpbxzk+pJ/WcL711Pf1gsb7
sxi9A4wTTgQOvOYV1AAtE7YbjrdvwI3PYflnOsLrHBe2pgXtGzA8yC2qDqatXodcFeQCu9zfFLS7
fuf1nLjml7bXtec6EW9wWXtFqDuSYPWKf6VFG0YBHWmkWWref+Egj7+wU1Hu0HOudt7BgHEwSYsd
vJmZYuYBrTcuxjZ94iM1ziPMSRuS0hATdZDzkUyXT5X7BFGoF9To5LhBcf39FVsiuzsSZ++mwzqU
sp5F8QUmfNKJELxbAY7bbRCARpRTu+ydVv1szPdKuJORX4Tx5K7oiCINhnh31U2C6+67T+5OEE/R
p/y8fbDPosxXsn7Sis0xy7NI9K3x83jrJOkrAMv0reKfdqs3BXMowm2yEVB99JdT5EOCy2FlPQa1
uYUM+fFO16jdLT95ENwpcKKe2yYXktb3FxSjVTsq1PeWQKAtb3gar52fRdGQR62z34e07Gegqc+E
mjMbjNG8G+wIraPEg2BB44N95yDDovp2qhG3TCYAzqLaiKxfq1NDiSCjUW/eZXoeB7AyZ3C8fN2G
0VMvQXDnQqAujw7U/YC1NLWaNGAMnq7Iwiutu4XtxBrABHI+SXdjooi45ea01U3jHOsZCrOoj73Y
mq01u+kCENNlubvRz2KmNA2JULyc55LtQedBOVZNU+gIGpyCAeYwfF6QaipCYP+0JcRyGcp21lL9
bvn3Ihn3EIW4F0D/d96fJ96qhoRsQ2YsISb1UuIDIegTAA7CUgN4qUyDI/E4UJDTqGg2QxYcDDT9
Kzy9YP8vSd2ItRKHvQ8HiEuuGhiu3vNDhyL/rFAkpwGJ3nf1DUngsc3cEUhIpsCEgZqbwOGyOOH/
jIU3z/lbOchZM+WWvxETwuUGmhShyxesaJOW8Fvo3ZUqV+U3gJUUQWB0ZwmKUNmx0iQuugxlVG3a
p8IOW4ZrfspoCb1/azFI4T/qbt+KmKuo44agL1WRi4f4UiamMWvmohwjyTlpCBNwioXaoHqKz2mG
fTE3gioB5lIem8NPXYO/N2xF101JsxXGcO61+3+gAaCTJsygr78OfSC0L2ewUcOS2OYK+KxwxpdR
xgCSLrOYlKn4AJiKRAT66USGyox+yJYjUJ4ezmp5b5+zYg9x2UlJL7mvHp+sK1Bo3fKFWb9OfID7
tDXm5tw2GjviviEyKummJezevUoU7h/N4dGQPL36PPtMWLtfRYTQaqqyLxyaqB/ko9ATKi6T2LZR
KpJ9A6lhzMW8p6S7VSAr+bdQrAARV8h24QH7EhAg5i0vdoBywmfd/JdBr3TJfvQTm68O1gqimatR
0t/07rJWs9aTQ0HoCXaBGUj6znJhEK+G8G4v3WwRJy3hWCy6cEnfAyXBXZw2fgy9+W3EwNzHiA4I
jP3C5ivihrmtTT9rGSecWc4knx+C8mN1mNtS5xptwN/Z7w1RQ2hSmh9NZCPKDzS34S95gQ36fF5n
vDzqstBwqELLVTAd5s/7soy1QM/a7Ajih4vE8KAub9rXT5hgF/I5d7MMWo3btC7TvbKf29xdeMMk
MT+/0jaPrxl3u/r7Ng048kQlI6N2UxEYiCiQZWD0/8WyjibXgsPfHeU8EkHQAbg2nePk4IExFlUs
uCjC9wo1ysNNWtw8XgIdrMp7k0AMTyV6U3sZ2lC8u1ugUFR5jrv6Qgbog5S6xkKHAXg8sTrpAAyu
Mfg/Ot3/F1F0PS0wn7LsEjJ4E13K3OCuVcP+3uq3caf6ya2NjUesU8xQh/yI7qmcnOFSFtBPGEI7
8RYcT1MXQF6P6ti0uvRIFNKsWdms5INcb6dSytwZpzv7/UWgwm8vHQnu54lxrzkETp79cB+21P+P
NfzOj4MJ0ZguxkqVMMld9pD0On9jcfCzCiJ9N2FlAonwNGX6N3TlKh2mPR8NYU+bQy8XU1ZKALcd
Ruv2w68TjJ+0QMa6KctCPS/JKuzKJZDQ6Dx1wq2BxS97MB3kC8egSh7L2DpjCs/aysXIia3cNovo
uA4OM+GkzHVA0qymwzlJ1ou81TVHO1eJ0HsrzrZj4aVi9T3vgdyJ18udSKzSJbAg6rLTd3EnqpnS
PZ8Kh6KdlGQxLWN/mRxH33hs5LgTKub1X0f5urJcbN5x5Py6m31y/SXCmNCK2tjbRbr20Yrk6og2
FDfQhEYub04yPu6S63fn0S0OVLkw2ir5Apwjc8SueDI9zmVTczWdoXfA/azxa+yNLHtnSjqs7wrd
UWUPhi5hEzycjC74bQUwJA6ClvJKWGjTueVxz8c5Fc5MdZcTjtSSPiwsda0UGnFNQguPZLnge9wh
14g3Z3snGRSEGhILlcGGEQ7pbJ3iFzFMk0BX9dsKcPjWTzRxPWNTJE7wWOkh6D2vTyC+1ZVV4TZO
GmSmNWOvBnEHk24DSEm50OYo6meCYRy4fzImzdQMqV0sGZgnDXEVkWE2kXp0Gh7PYxVl77SVmLeH
ts70mFR9sYN/DLrkyiv5GymlystBT75GDSFESf+EA3Q8DHZhzC+VTmFtn5Ja9nOmTY9thk5psmFp
nL1Qg8tRgHkYHft0Ny9cUDFaBJoVqxOb/6LQLfmv1ECJru9gAcjKlO4wwV/+VNrAWLETaMHIA92r
qhyXbIieXQ713tLUHCnvrRA5ZrQ+tMYpJFi3Fw37MjpwtTi5YEEKMWnJRrM9J0mUEhy8WCIYdTiw
SOOQTlAtI4nHrAvSMjq4OqbIKd0KgwrgY3iSyZY2kXYlS0TJVyVdLN3ZhOA7z11eSYWiWDw5Deyo
pwIUZwvdC/efMJHjQigWNiZlMUv5zrNadoFYXi09lPtWlXvzhUVpgsrQa2W0dEMJR07mpUAEwRjQ
6J9CpiZlOY+KwPQ9yr1DydduMVJbpPSBrYTqDruYY+ARPpNwpMMdz4pnQ8qRYg0aT5/EgBu5sUQQ
VN8RAFUM6QHcwMm15eVNrdhGJwMGtGllaBebRB+hb41ws8I/XS03vi/s9AzEaiPxxx0oBZha4keB
ckkNtOzbil1LjFHMEYcKVAEHp9GJkaqMrHoi6m59h4otwMsghcuZXxxHi3u4PzL0NWHedxVPuJXc
zJJ4l0wcYrxNtaXCzgVDREB32DQUhmpEN/o2MoubG4sFr5RTVvarCeh0jD/8icTTFuuBuJTYioSv
ot3mhVCdBBeLSQ7G57/ssMfJQkeFjaIoCASRqvJJRR6T5vZ9nXbonFJJozLGT/IgHPhZD/3X3JOD
nBUQ2eJuewuOOGnc4W3nt67oSThDRQXVeK1D69l9YII24MZ1kgP0wO243swngb7gKQFY+JzDme3g
p9KCATT8MLInlLUfD9vI/exjgqxaFaqfV1epG6+ueLLBO9JgMJCk5k5u+thanZI+STE3lfNcZPvS
ip4f1wgka+DOoEYvKQ/jnbmAYs37qe+sApQbFJac4glbAzeC2nJvdV8y5NuKxlzG3ose4apzwRQq
Y9cXfYJsezVPxdlS2TI+JCzY03NYKJK5pAoSTp6yzrt+glolhA83ElazFFP/mCddj8j1p3bcRGZ7
ckSWelu/fA6AQebwaX5TAYnxDf2gEC3y+xbKylMIlP8S5kyvuUOHPGSAb0lc4NCIDmmsD/2iX5kF
63DvZw5ybGkvQXxk0WTuJ3xmg8R3+47UQOwNljfQyag4qjKXn0Cm+2TPo4FF+ozKRZhuzzlExFVM
3Wz2dxfo4RapEeOdmntIY0dTYUeymT4hpN0sO+gQYj4ajLovC0o1j1CD15m7jO65zUjUop5+lGo8
JgI5myGSN1pK8wQEXCScplkwmeDfLiWKJJ8ThtKm/sVYnAnsY5IXN5IyB6Uek2YyhLIFe5MRpRY6
sQKmXwE21y3bZ4wxD6xojZ7FumuLIkJXP1rQytJNcGvRulNqUfvMKtYw+E4tcIfUCBOdCIY/MFLi
dKsWJKO+QRJ3iO+rCUZqN48NDSJDCELMk7C98S13df+X3lxachNeHJQFB0g1+Y4VKl7L/qgVxaxd
Xg595aCmSzwmF41bwEK3a8jakWjOIwFGeOeWgOSW08lWjajJB0PWP64BbeXm58LgRjIMaCjBJwXd
0I0dp/3ZUjxzaUfuMHz0Z7kKQ+ftuvw5NAB3J2KUzAG55YYz4bvxPovT2iT7lUB0fbC2kFO0xMpt
8ejZjH30IyQ4XycaGsjfe5pyERZe1pSgLn8OfDU0U//kuo+xVB1OML/hXJsPWW0WI0UMI9uV5vmu
wG4xS/Gbt/ELIzJftUBLqGoiJiDg686vQG1Jg18if02NL0tLEVbNIh6Ru3sta2ywdiIpNsTUychw
CFlVpKFdX484sA/Emoi0T5yRrETJJ2vGaxGk6TEhT2hyh0oD/jVcTuSaGtajrw0q25Geaox0VKC0
VdnoLpEV5RpNcL+2WBiQ1V9CoKnqvdotR2kyHiDiKGp6u7v3qpkuGkxY9RhKar+P2oJhSwU/FzyK
x/yf1DT99HyogrhoKfDn8f3DfM1RFENduM1pIUt3hdpVkW8IgSrz63Ka+LhII5L/sIT0lKZkbMbQ
TNDeeMXptFwhUamg4oG6Ntv3mFIzxKiKBih+H8X7zQXx6vDxQFrfQGDww4sMcVAFRwNWVybK31fC
Vwe+xus9R/1RGBo4DHaKMcTXjKDCDT2HNgGP+CHwhzTcd54MQUnEJyKuCGIAR/taJiFYgLyyB+Mh
z+UtgfTrSJYDpTbjg90bpkXn4uHZHaUQcklSvWxyrKKp5UHDQRzY8RD7jm4yAGMMme1HDfSjJYt4
F1kBjwZ6jJapQ/1J9DGkaqPSjEX8EGQ0OjbResl4j9sDlGnz88P2Nv5zhaMnXXXI6ZsADaniwMqO
BfS/p10sstufDj+PCFWRjKAoFCQb5RB2AqIY8cLpA2DULpDPuzZB4mpsAD3fVpgKkwP0PgL/ae8B
z/2O3a0/F7iL+t77m4mK3tdDU8eMjDiYNyO8Hv4AQH1q9ggMEgcQl/6tDxJpeOfeQ+GB8cu9SFPs
H5h5TMaTTLFHUsad8kJa1gNGwFvKYzFi+DgwB8hdd0EqdcCyjoH/v9mZrTBvCK4kxT8i+ytNXCP2
IK+mDpqSfLW7IIOGRX6pVY9EYRWwc3MCGHDVFK1O29V986Ets2esPXiJ5bEHB2gSDTHFjL9HK4OD
JY2y/aL+zclx8Lz8kB7yVtdu5FLDL7Rh9lNeQ5bV2ijvechfFlbJlreg5oRvjKiVZQ6LrGzXFu65
MJ1X3xOloyTb+zzNV4MqzS61PXdKAPhD5agDiF//kkvUG0rIwRFPMeB9fNA0w6yOh+zDFvfRehFC
u/FHAO37wx7Euyg2XsxvuCfzE9vQ689gdTMFcxOU+Yh0vg7P9mubgf2Uc5aMWPcmcxqtSJ/hVSZc
iul1xHp4E6CJ++F+z3rDd4eOaHG7TCYhV+kSwfjJyqPGvTdCQO8RtvUzcpWdQDW3GJaADYxlPrUM
96WPOfWOnCo66HRlzZggE62jJkvcvkZW3zEUI6cTIZsjAg5Sz8vu12/KTaknV1a4IEzNEtM5wKgS
zSBHgRFIANJAW5sgMGTVNHjwsybVKhuwHXgQOVrH1GZl+wlDnCYOCMC7pj1nm6x254yI07ldTUn+
5gmbruNkKwxcyPD7YR1HEzFthB77hF2G90xsujgfvhkhGdOgLVXKY/+WWXieVPffzAKlJb2B9reS
VBGmCx8MwFHkycanbQgi3+6F81CqOLjSZfujbQVffzR3kmUzIZpW9yjIh69hZ4NJ2CrmBJegNzJs
uUALi93H7Y5wiQQxXhIWl5Za2phRewF7QemrnZngXysgPJBg+xzvPb4y6hN0GUwWtmX0/iKqs9a/
qq3p1BLoOHXmlSxO623g3yn7hk/C1LfNjigmT6mVuLjr/xoh/pyl+yNxUIhNiHhs6NTJXGsawyQl
W+7Hprbc5UCLIYMm1UmaCD6QTc2sIltnUOsABfU8p1O644tzNNErcvVZnrfMdRX1x78qmjY+BeUn
uyCiHuuM/q/GKtPC1WA3E66f7P/fP294xceeAybU6xpUyfRuufLrQ5RpgVgbFnPeKn4Mt2H5uOS/
cDAOrw5E4N1gsXy+ULDY9uC/gZ6S2lfhJQQD0qMFAfSJNq9640jGtkWM0VIfw/2q7WU8INJRyrmO
zT/NVVvSr1YoRUGdeHldiAcBl4tiTKePQBUjtqTQj9YjU2cKkeB1dJubBbhR5jacfYicHoIF6tha
lJrsZ+lMSsOH6Pz3yNb1WDRW3GdRMrp9S3e/51iZND6oaRrgQXj+CjuGoI8572cGpO9RerTuqF5n
vZqM+U4VyhTeB4MMixm1Sj/P8R0gp6pqWU0O1QSyYRohccwdxFiHUQzn03G27ZOD+CSOTeY0F9ex
bAzKrsZfgj/Jc/LIMdeLzNFuZoKyydKHYy+2uwaQ88aigxRtZ7G8L9u6tjKRHgqc2boPycYyBmEB
73vDk06a2/zTUcaAenQSrFtdw7i1rMut+2i+pILISGu7zS7I//2md6P8uRl2HIIWCsL6Qg7V2PKn
46P0q8j5ahE3DGx/VgpjBeCjxokds4jt895cI5IfNFB5GWhA7P0Zt80sZHVbjiLMqFELg+moX1d8
kVgIYxitnnGhYUBUlEK6nwilIhqghU9BXAZ4nI0iehqZKE4zVlYYooxlTxzMKaRSVcE1CZ27lsxD
D6oKzOZ3joXF4eQPrPILyAT7ggLTWJBTm3pcIi1p4G7uV854BRbs3RgYHdjFnLlTrJ29lx6BToGp
UDOISHY3LEggOpzd82OGmrBhicbn/0BAUx/vgDPp14+v3yGj8m7W0sE7j7u5ZgXdBhCM01K+ldwC
qyK3ePfj9gz50+AOf2f/wbv3tc7UBfIMNU28/zQieu/pdPdy6Dwog0TaCCnsStkDahVoH8u44xF5
qwxVHxjsFRnzryVmBrZxKCZnYxjYphHRUx5zHmsdVWyYSQMSNy31zFuZmn2sc3qF11bYON1R9Kzx
Vm+b/wM6kLtaC2BLyJSKCAz+rxLrVphyukU7Qdf7KuBVtHc2APXMfvhgAiZEX3AJUtVoA14cijlk
jJo8z186kVHSqGBP8CTj/EeMHpTD3qqSRuXz+S8khwrSpbP9lHpIzrALBrTLNhNHUWlJkKKz0fvh
MB57iFfWVdcXuQ4QC4QQyTwhI2GPZNcLYjoCd11KU/xUc7seWl2z/Gb23l940w95TOKwF7SB/EI6
n0zhqoqpzNZSZXTXxW0pXt22SwI0M1uGsARoN7xOlTeUQb4NEKa/NNnAH+F5WZ0zQz1MNKQj9RFo
9K43wCy24s+NLr0xCfyXsASw1qA/flSzbdebx04ApnBsHQOnOdx95S5aQhTUoS81m8B0aOUnWN7a
Yp6JniLZJ5Xyzm5m7MnHTBcEgSEi1Dc657ZjX9fKNcsl+uCSBcd9QxQYVXBLZYqclPuCnsQD33PO
pLzDoj0wHiSMecXPRlLwvroUwp8k8g1spg74tmn0S36TzvkZUop5JX69UO72VcDOTgAyTHQU/ulJ
jD9y11v6eRsQnfqU5uG56e81BDSQTR+qIn/Mt6Tg1IXBKHWZ7azTa7CaDnklK+6N8iHP2USRYXre
W229H7FPc0uyFXcu16q5+WtibYoLlJ3+rPWy+jF14H3FHMZe7QTbW3381hjVoFPkQLBqjnxt66Rm
LokrqMYCiHNFi9JYcAEIINRcRxkg/XSWxHlzbM4K11eUHjB7pfRAsMYByqTUENoCXPbidwv3jYTe
pZOOPRtRcX1T9uGYTViuamR+h1u6bvJXUoER4DvdLT8ESDCcrXq6m0q8zYLP+x4Yp4gmsbGJBI/p
w8MxCOYpK/f6jdIGGITfW6cBDiuDYDgN7W8g4fmM3bLq9Dixfys6FfTrFieVeBZSIdeD2IQoZltq
oFoSaol+3jiCIQ3nS4edSbauxKe3GrHsQwKk/3wGt1jXoBDn6sLqy/4f1hap4ritUvRML4TM2pop
UHq+Ozgakq0A+4cM2kvUDpR5Vh4k9CCXbnkxMYoKCn253t/3GIZOdogcW8X2WNI5BL1s8IZFDo5I
Ft9X1L8846ApHvlKwN+0Ixoh6HBIPLdK1HcxH02vsPAg3iSmLR9lDRkSXeGJWQG6X+9UU8kIP+nb
1vC2Dlla2Yc1J5rYeDJNyfr516i+gBMdcWUWU0kcntzOR4N1k/AfPk6W5qCBJDCAS/F0BpUUQc5V
gr50GYClJy+UlO5qOz0HKbUnQ+AY4Jd5wu/nuhKM5+RffLhpbLRZXFTuvXZjpfqx263yyOkQ+bzb
r+lagHqsYrEpELmcqiWZtoPu/cAiAGbPUR8LgbJcCydlJgBWYvz04PxxCN1sv1MRu44wle8oR8Sc
EXBKjEY/Jg8RI/MkT3+2aoiIYKLCojGElGVIX2w2VRFfnUhwpUupTL/dcgdxtT/caSYaBLNdMzBV
6df7qO/kpPyBI9XKOEeE8oQ+FnmtVxdHjT6LwCQnR0PWe/IKG9DG1ZtsoEY6inkzh1Dlm9iLnIEE
Z2sBmcF8RjF4Rx5uikaoye+7lf7N6kwscH/EiQG3GJQNC29XsueUgysClSWVqCMxwoOVaDc7VxQz
PYHRbRBiygLdSRpdt7/YViqsz9ftAdhqLgrNhAY0gPd2fQBmg4p7yBcUwt+XKoaWHFbJyoyNGFGs
78vi4KRrSfR04X9U4eSe60WqTjHAufAOcn5fEj9Q99FNjdaJD9djM8iw6+GwyJxY4WlNAFfZe8on
TktqE4vEsuVSXqFxN4gEl7/YtXDxucO4FSZdVTfW22bVXqnsKebgLTjSw4N5+k4ADHWwOKUJp3ya
uKamSrQmfDQNikgrEMJSRDSill4WFK/ig3QQ/jblP1c3ob5Pc7gaZqyBVdpTJ6mJyvtnQur1MIHO
Ou9OSADOXE5bRiiRQwPEEVOXP0Uab+oRI4xNQs6oZnjIFQOV0Bjf7QZzZFW/QRvhIUm88ugHOfcp
iBMjJdYVVFchYtqh8riuhvzIrYcK/J3AMQKKLO/Xa9dp8nPCa91OxsSOeT+lqgU0EodB3Nj0YbCZ
oEtk3biq4mMlPFgQLPuGeM3KFBfdHBXqW7H39RD74R4XSyauDUqF0tvBVrFIBS3gCdV0e5dxxRC3
tJs8tJyVLdnWtctawqr0JVwoBF0J8p7FNLk83e48xALRMBZkohmcZ0ZcVu53j3spFn9sfWTR25Qh
cyEXzjux+k+KiL/ZmGJ5tJN6YAHrCGLXy55xqw6xbCisfdDHlMEdLHLUdRAHV5pVSgZntdA7yr2P
dY8lS6vzv5wAhhtZZI71CQCtsEPDk57qa0BMg+YihXwHn+WXOsRe08WyEkuN1AgUU0S6HrDBwx+w
9QTEQe9Kz4s/6IKndb98AVTqm+LjNJ4YDhuKf/5ektlthrQHEFmYUeXvExbOX46uIQOAnrXB2NOn
xNp/6FNiiXSzYJAnLwSFnnHZT6lheKktWcRPdeF8hwhWvRD7v0QKCoM6dQHPvIo24iZ/sGEmRESZ
QUTfBXiFN51wu6cBTlICpCM+Tg/N6v8E9n50I45wA5x6gNmLpzT78B+iVRszgpCpYVknbQ6tI/PY
EBKHl4PVZYGVHdD3w5R5szpKxJ/zxAzSolHLgWH4KAnEmw9acbfOTEmdpiQGgNHD51mfhpKQU6XZ
uh3D8Yammr3hSkp4Y8N47SbspxXLzJ1r6MHZeVGJjsDIaSDtB8x0g0G0g1Ense1YSUDy+KNyZd28
kZnVddtHGj3hmlrR7b50GPnFAahLX+nj5M9hZo/9jC6wqKdVd51DOZbnT7XnaH7kMzoM53mg4XSI
d7/eLZkcixDG40gweR5Rb0Wtlla3k14m3TwSzk3TFL7VN4F49P31Oc1o/YIVhIy6mqi6u0tyJPTP
IHhUjtZkPdb+VYqgJaSZtBtLH61aWGvnGFc7FcvOkV+3VIW16vtI/0jyNJcVlfKQ9BfivbXfK6sy
UU09sSkD8HogqpHn91z3slP8i+Nx1xcOxbWE8MpAqUfe3FVoRJUT4NWtMhMDuLkUEG8L/CvkFIhY
rl/wj3glmpG3s+XaBaT6lI7AR8LxGiBBijWsUu6Cn+kpdXM5cQFw0m3ZtL0uKVSHhABDNg+e5U6O
HpLvVbiF+CtMrE2FKEBVIegzh/lcCua8lBQfJIabKpUItQykNaHKKOuBB26fRwGo7HUNznPXow6b
z7EROevmic9OlkfC5C54qSx4oi51Y+WJg6pln1EYbr37LuPABLXwQZt/zFR7zs9Q9s0lpkmCEhBy
11e8XTg1k5+OotozjVsrM001vaFP7uTjpcKcDwGQczk0ghd6ULRWOIyH62b2YkAFDb5IJdwQH/bj
eHSCUR2I9GjFMVAgm67Ap4IRUKYyo/Joqbz7GqKL3aCmcpj6FkEayiLrPW8J/lx7RjevVkv+vx9z
pEM1DWiBGyLMtN2/XiR6wJudvsAdXiCRP0Z4NqzYu0EXiY25hIj6UJq1X2r/tR0ndxXx5FkQJIEw
9tif8YhIcMzoS9T78exEH0nYmpr+Z9ta+hm2vc3Ac4AtpMImYAPfM5WGXB+8ubwL0ruqxEt/kJpU
haYCjiT2xlqV2Ox4vIgGkuwyu0mUGhfgRZfm9ZWDrVN4i/nHkF/jViu4SXDEbk/NaYAa74tqOz4N
h7dMKV/JfwvVIrVHbTPolukMsFO4eJrgUoEYhXqGLcyD9/JHSILeRL9Qoo8VMwsabJ+H7uSlM6S8
CVVyQ4qo9aV/WtNGLjnz8YZ+ZnTcg7ANvsSmmoOfub46NZ//1K3c+BnuHDnQ/oPzjBc/dMYvi7pG
ZaHgPVSyklkcTNWmW1Fi6AQDo1FploCARCgnp9YZCPqTfaKDg0kgrnvjF6oEaoQCnKjst544rZ/f
1ilUFyelNslbL67dqYpy9iTxdVUdcUqaVBuQ20ADgfqg6eoFVrsB2YqGYXGbXeY/duel407TFERS
a06ur2nMMvmPPH5fNAED3XY8KDjTGTSPa1rSq78+0M6gzV0WZNi055vn0rlBO2oPOtTjcAlOi9Fy
1VqfUF/ONAdpGy+bwqjlmbAr8VonnXWfMYxrk1tLpCGFKg5YB3cIhQXnBJ886nHBydUVQCDsuSb1
CNNa13Hr+A8QOhPskeuwrsJmHdhx9UyK5uy5w7SOp7ImKfY5Lfm6yD66vMyW9LVGDFFiDi/GL1sq
02S5o6Ltk+OhOFkSxvkOegG4AUVw4fNYiovY0SzrZwPAHYI9x7AFOSwrfP4nrCd7JdHBKsmScizJ
7LK0etQcZn7DcOcKbfPnxefmggl/etP1ECh8vvQ6irveNtFeytGYr2iAc0V0RjBbYixXBaOOLUOo
WfcwOXkccelLaXuN3cn97eutyt66EFMdn+G5C7e+UoM2/SodbvkhvkzF7RTqlkQkRlD6//Q7RNH2
L2ZdXf4+XZ4V64BRMugCNGdJ3u+RUOu3WLTXIbsjrlPx8RAi69pnldLySvLjlupxJCUuAhQiILCF
c2ZNcm8RXr9wj1WyZkNMFUKnJs3i5pMrdIEbzlwSem4J+rhgeaKi80p7dbgpCVm1p6qHybMbFMFv
5gQxsk0VlGevHJCdYakRPnaakwDrf96AnFBSluRCm1x55OfoFZbsBVUeJQ+/fxbxCIG2MB/z2U9c
GKX3Vg1rj4OQTfP26JiA2AG3YvmdMvzILX2e+o7Fr4oc2pznegVQ0BKssLsVgOFrujPwTfghZrBo
H8mah7aAbPAzSy1PaO/IMiq2/RExbQJHFcPeyBNJ+0DjfUcLjQ7csiL2E+o2dri5MjgNsLsjcG15
ptm03p6TBXNwkyPz6CVkAwP7eemiSSKS68+2jJ5K1MGqAFiWRwuMY1KtCG03tlnwJy+vUDa2FRvA
YoP67QXSdtidEoaCsGyWWMwlPflyyUIr077HXza7NRN3f7VFs7sLPJsu/5Mzor98rkWa6e087ev3
8a2bPg6rcT0WlQTMil3povywP0ihq0FHk6zwKlNnPJQeYg5a1H9mROIjy7Jzv/68kJdq/zn0Wf3J
OKN6rmwSvHAfUOPjubDK/y5JQ5A8Rf1VRBwyK0fiQPdVRN3/gTpWjBVkchjv3nAYlDlZ/qD8E5Pm
ziryU37Jea8Rk9BEAU5OV/mp/xFSPpR73n2s1F2dbD6MDs3v35OtnsrR4Sz7rBmkJzJMhMmQfqyY
vyZEUR13q8Ow1+afUKtYgoyH6FFVtSZE5QQTC4ftwDTFbkWdvpsiwYpNxnHKvGVymdZY2CFS/YEd
KQKTHzUXFVvLy46qLeUyu3/qBmR3cHi87wG08Vi3JZsTHIIy5UBeR4llLxaMO8JxmFtqSHrE3c+V
h0XTFAxbAFN2axsYR/lPHv23fGq2tT02MKTyG+1O3Nat9riYocf2pccn7X3WQ3M4/ZnKIi8BoWJS
h9OKCZgN2pt0Vf+uBj9m7PHtfZA14aMajKZ06gEE7bz9LRk4JaFDnyBQSf2YAIcFa/JE7kVoBZWJ
YlBik+Wil3NHLI9TxfJeOd7IULdDSUjBF2Qqt8JZQS14naCc6DKfPGVFg3WHyz/mE7TzCw88grqq
VUNSAQMSaajHp5FP1zIap7XXK0rhVAHz4cB1DjbuMXIJiat1BMqyIS2OEwaPLZyUR9ox0w6ArCnd
VzLw+iB2HiM4EDpo+DcMxXyE97UCHaGOMEQ1d3e7FdtmDPv6s3SYWwVicjxtfP6O3D64/DSWF2nf
zNHyJbirXS2oVZHjsDnYGHRBzOYyC/sXcqEtcoVhn7EHwrQXt2Vx1NUdIA++xiFG/zdIReLGOP9c
2Ft/MdeixY5sWDr2I5HtR2+QkuPY892V7THr4aOMhqj7XDeLxxsTlz24CTE+1PfwVUyes85wRf3v
+vxufsrdTEe+mj6vLMSk1vhR9ouOTn4u4+uTxj2txLxQTvyLpTUN0ozBh82YHr2m7tF8SphC0xa7
DD0A1Ank0RX+T5TYeDhvnV84JlsIsAVtplTjGz6tT9/GHy+fQMUNChbUTLlYJZXb/kYSVdZ+radh
Ep9leuPURlj+A98IxLM0JsZB15/lILCURwqj9Xv5vhCneM63F5ga8OtjKZTFOySet8te3ol0D+dk
JxqU0HtV6teBOpBjaPDyz2bPqQKotyGN7AZWBv8/O8BtJhGwIiVrN89Ejqpzkc8b7iRw+RZTrnbz
Y7oAN/trZj02+Y5A6Z+R0v7Wm5037iy53UvVgUnz/JElFbYW5pVk2LT4g0ln+MMBjZKdr53j4kE+
5/M4WU0TPtWFvs9J8ezt4dzwF3WEOvMxRa8SXy5ZkihwBjltpa62sOMuNJEzq+PLL9UyO6z+Cxvs
p1jmvkpJTAhETEl8jxQseRUJes9e1DQkSFfY5OQu1lthRfKk8CzZidPIAhiGGHuuwlQTlYUq06e9
yVNydxJMKPR634ZLAQLoBdshUfCYjLiZSlfIiBtjBauFTxIfuSkm6WyG+mYeMSldNyq+PnJaLRJ1
UpSBqgV2AxNBC9qi4C6+NqlBY0nS55URqzjFodVSPKrekCIWo01XeaqQpzsVPALOFfMDVKVrYuzW
fNnW64uTC4FJvQrlWO5/fMdFq9n+S5DFNoCmiwk0tJoyYiqDs6lVtEBqQYAUSgzb5axoDk9arAsQ
bTDhb9Z5zSQUEwrBpWjnIvr6yBpFDGR0UccBYINECHRGJrHf6/njl0cBJ9EY3NIwyJVermMyoBw0
POcdh3U6xMdNT5Tgv0lIoQMw29fQy69AAJ3/dEBokviViSFHjHluf1CAe06SaFIdkYZfgqBF0h5B
wZf7iVwiOgBiX6db/8oh+XLdPeuuxqDmcufEqTGpzWGKyVpCAW23snkYbP7VLBNWHX67lAXAD9sp
RF0oAO8KhllhhieC43kNUOU8iZ5W+hHMcMSCHxuDMe7cHVlrDCXpzJQmOWTHxbD0rxuGHwub521q
L3j/0sH72jEPSF63CmJKn2dbxnuOGkATGB7vi3XEYOaFsVKgb7b09OWBtPLkMInxA40VSrln3fq3
WB2smasCbnUUUR2PBTbgzlmG8BwR+tsQXDU1kN0f+l0uYoo89CODOJVtzOb5u5WIhub3PjKa9WPw
8ZFQi7jKNtUlRR8kLhzd/27BsADLmyt3z+6UTtdGTZsNNbWp/IM3MMDqsabafTWgrY1NO9Rh1MTY
ymwSsP52e0SAzDg7xQCJzmdSwpcqNRhNhEdv3ifziKyZk4FA3UeJ6S7e/z82izcTkZexeFqwBqVo
S88RvzDlCTzpd2taZHDGInson7VpXX7Bg7KzTsBzwVIkMg2VnA6jCOxVYHUk1G2UAv3r3b8sdjEb
38fzk229LtnEqnyyDKRbNCRJxVQF1s7VfyfE73+vBEH7695LeDBIRJuweMB957mzZUzAavrE6UJv
TDQsRc/vQUyY8+CvFnEBNeJKhUGwlvhNEcOGuZFTtj0V3CXG8teYG9owI0DNRVBM1oU0rPZ5rDg3
XGsep72o8y6KVhZmp1xftZgbUTbA9cocT1MJVRol2UsC94agJ43wkh0i5ApQ915EV92wu4IgmNHT
+jYgcjzds1D93mwX9NAcUHbO8cOoIzb82M0svqfsJuMeF0AHMtkOKcBSivV8gDrnkSEwUMuzH3db
Z8cTwrNeXVObSMPleYbfXrZjMVl7t+OyXo0BHaeKyaBQCaB2csKrpvIsxy80TYnLmRcmgopbdajp
cAL9OVBJCP/yapPiyYW5CPJQtUJMm5NWP/8EPYbGwvtxpAGN44YJvEVNhIsggT+YXp6PEZWurSoo
T0B37w3VWLmlOBS5MTE+c5pyqCW7hI4mNflsVxWnppQHYlAD+ATCm5OQR83BGU0ourj5lg226dtN
FSboEmM2SmDDEpQ1PSJj1Is+B4Qd2RLlmX40qhdDPHqqwseDKA2DkpKXvoOlnWKxYw8pf6IB2rMJ
JWspfNGKibXFQIIGYYeuyZ/2Sn0O5OSLtqNzPiCrj924ocNJczgAcKIHnbNs2IWnuCIyFB2e6R48
IxQVntF3FUmxWKZDC2NBSitaYSrFTX1/ZUIneElckAFirHlmhS3imkOk9usJ4ApAHM2Ic+zXXtQ9
+fznr/wYA3ZKskajRHSNITYMc9D0j3JFt83538iAtBcAs3BKkZexrz9hjqEOaRXokQJnfPcHqK96
CH3wKPC6ZajlBToPrT8v/1q0G7yPka+Bkqz1FHAo4oXdi8QvZcjljesmGJJdpHuygLWYk7BSPA/x
qq+625FxpR2eTLghRuDE/ckvbV6JAVBAaN6k5QP4ydnwZmVv+58XmKGG7dquRK9rFcAQOdB4GdZs
bAWGiN+YRA14he7Hhd7AcIf+lOvLqCN0FLJ8Y0/M/gbg4elqrBk9QmYNbKmhjnYAMSLnKdpZcDyR
IAHLzeFir/a0ruu00302Qfyp8XL7x/NO3EM7fEuMHzsjbMb8o4AtwHDLP1mWA3kL9L8W2ODcdBVw
zi7linFOR1lrkV0JMdwL7LXGc6BsJTTKsLvsK+Kp5WivmZdvRjTRY11InXhNIELD+f5GtRCU7aD1
RDfX0u54LZ0JPEGF90/hVNnbpmQBw5XV14zik2DxuFwXENTXIXlYmZ2JPt/15kmlorGwHGvtMF+k
uM06gVYB4mBEk+UJgq9eT+QD+9HIw7AvVvZeTm7EtWydeUggjeMKKhIZPVPrfVB4XCemyJHBI98b
DSH9Sk2HBfmQVrJVJ/CbmY8GdBiubSwuT9h7IuLxruSN/lns/kc7DofoIhfxhmZ/QLD/9k70Oubs
514z8hdRhvAmSGcs2KbFRiRe/1jh3BtHOXQNNFmpl+Vqzw/l2ZjY58VSMrO7s3dDBqvHDMo+orHF
mAJusHyN7/lTPuEAFRoqUIC+beX1jZeuGThRVByb+wpYawJ+0b2k+MRkItPb1CHHYXOhuaoJcIax
SFPaX1lpaOJgyddfp+REis+1HFMT+2ShO3PB7xy+6FuPqwZeGc5uDWcz1MhiQiw5lEYKrULh5jDs
9Xc5RG2FyrPPv4MinHq5QPYPVxDBtYngVp2i+KKYgoWAAuSIgGirOAyMJn3QPCiWkHpBAwxsV+bf
f9CPESzhbjUICWjNX3Iq2Mj0IQwz3zOx+o74NsgM1QsxiAEvQmf+aThu2iy73ob8nuXV95qq7Erz
3+ntXEpoP+qz/Wuj5gBFk3/Wjou9bddAibC3LctGdW9gb6z8j4lh3buBfCQYR/8Ov5jS4mmW1jO5
LiMw6jZScGol5QzL6u4TMQMAl0Xi4fMtSkQjR4qIveJd/TfBe/mZRthJliVk88ku/nEUEBslnxaP
kzzViRYoll/U3AjHyYJ+gOaPAMTi9B6JSG9zHyhj7cVndifvS3FCGMYfSEBzxTLxR0GpdHVqcYlQ
bakbwoFQCE76sHcaJ9yNxNDKcLcAO68tXG5GXoX/g+NTlsmteUbXwpOx/9W3jCdnarWkziTMY7X8
mZmXM/RsQmQn0wi7h9WQN2KRpTOBDBgMRjsgkipVFqZzR+T4qzEvBOIDojSfnRwiNAwSdR15B07F
F4QbTYDxpjI6UidWaCF3Mu1Tqe+MIcXGX7fQr/OMK4X4Wyj/M29Tpl/dJkn4mJEDMG+SCWvdAOLe
VEKbTNZ9ftVB4OIdeE9OQmkNeKeY5S6AqBnGvSSdzXlxXmWYM8kw2JSp4CEDmTjv2oU+vpxWt9ch
lKTI677qTAPaHytBOqn561kXOkqDQbN1vTgS5CBJ7QFj+OKwp+EGRzBe4AYq1WY0lWn84ogsv7NQ
JjfCAmUn1OD3b57zpMRFqbgoe9hnznspemIozVVHFibFkC5hxBHwe3x6R2TNOM8HTVbiplSZHLbP
/peM1N+o8TgGM+FvAHCCu2nHwOvPFZXqIQjSnpncWtA7E/wuyATuRK3Tf26hNr8a267ZmR4Zeg8l
c3aoJm/IRPTexGkdsFn2t97iIDKG0TLsVQE96tEBxsdVumiNvdasH6gW+XKZySGsWf2R9cggrFEg
gHmbOJNwo598HDal4yEVBZ+RNggV76MLf4d3tI6SHcZjvBfwEzRezQT0kIZlmJnQkm65I53DBE8n
JfV/G2t1QbYCkLX8gr41qBXcZn0BTBmHvb5I9gttviVSCGEL/pUIibQ5KAn1AuHHyO05z3EHYNy0
b2BT13ESRnygm+lmz4d31ZcLc8JctQy6woNAGR1pANUaRZEiWQbLGfnPxFq+HqEptfoq48TO+28u
Fe7LDWmwgj8fD8nKtCWoTLe4HRObA0z/DAGS0DeDrYKPhp2FYwwtHfFZPx/nYDToE3pm9SbqcYNZ
ipamFO3okkYq1+zXW1xZj67d/qekDgvdHgeN9hQ3Wnsw0CgTuUKkmU/bTFBhcQxIb/iTNPYqFowj
nJZIhTVrj2JLdJg7aMHiR2YDeiAKjiQ2OJoAUViWg1o2gBoLeWpijtyUT1FQr83vSeIpMUqnNhdj
JndLvygIttCMywa04Kj4V1QH1yd/3WesSBBt5R9dt9CWA+AI2O8dk+lN1HsZwt3NFeZVxmhhyOg2
yWnVyNcDS7rpWg2e1H0/5WL9kc4yI88R3KhlG8j9zDtv7hq4OsmQGf9rHD66A33Se2E0a9MobIUz
LAQrawYONDEzdOItB2V4ea/GnCCHDMSSo9d+7E7s5IE/lBM87yLmTLqjWlJwsOGTghIPL9m7kQkI
+2fmjTStRMyZmXv5DRSyqXFI68PRIDrLDy1svN1GxPOJ566Mvv0Lusz7UFdqqgL7ZQTViTc3st/l
cVyx2SbiqiaE2o1bqc231QQ509Inc49m1JYELRm6oBd0qKTOFipP1Ltblpo6cwoI5UYR5BGTsW1e
nKkX5iPbFymjeYqHP+Rh06CpXDqh7bZ2vFzsyQkv+rKzyOMzlIu1DRcv22vJhD9z1zviEYpDXcIP
G0GR5P1QKAwnAZlFlkvHw6hD9jCdCBe4dB6wUCTiwAvovETd8yMg+9rJVKGD+lXFZfcjEd1sbJeS
6+OCG8YiQX8ZeBhaHc7bD3bRxcPh3tcw9gUyZnuSEpsSM/RPjis13xXtca/sBWlZlQvuTgf703BT
0PBjvvSR7VOQOS0kSucqdcQGGGteNcA7d8A+hw/UjDQUkruyjguOzW3IC2QfWTEsUtUXsKcfO+bQ
7Q/j1HjpEVkJkZdQTb/52CdDw+Gjh0l/9wfEHw9Xs0Q1Of+7QewiOQ0ospeciXCRZ76EvQrHMuVW
rY+PacUz+ayCO/S3q77mhYqJeEXGyD83eM44ZGPBYGiKxu/gXTehGofbOLZXJqy8xEO4yTEQ1iED
0suEgD3UxmtblJ5OxpIkga8zEmZTjuuQnSzUZCkPg3uUB67t0/1xWNEuRgJRUxOER1TUbH6s/7y5
fbqWtSsOqUwe3oJY5AtO2xDyIZixRsOka1UZ7iGNXyn0Q1pZG6c1K4P0tPedMdPIUgZHFCZDSnFv
fWiY5ePBtU1BwG/EBrBJH/lk2ASXHRgrG1up6J8JmuaADOl7fKhfMncomNQyst4Y46kEYE5FySQM
/UYiWyESdBlPx5QZdIeIiDxLnCQZZtO+23NTHOMsBBHcjnPr+j08kSpYGK5pcvszkxsTSr8IvRa9
vRv2jVDBk3ObGpYNgswvQbcfqTUDAzs+WqROfT0K6E2o1QnZNI4No9sOYaGtWjKzA0raoRBOq2It
gmaEdgJ6YNxmsEM9CaZ9LZrJvZdako0AqriAfgkcVrGJoE57R+uUIw7hClGGlDGZW4RyfceMyD0Q
TqxNM0kJ18jqw5jSjD6kk3S7s6Tfnox9PE40nznW8OrbK+75bZXfK5Cwn+6K2PEy621aHtB8mIUW
FHYoiZBWizhhF3eFxM02S1Iatr6IstnH5MqLdC4Nghb/XCXHhtbunVYp4jMSZADCdtT6yKSwOs7U
xmnNfu2+WWVh+ovorXAu1qSW/qEJoSQRsZGM+z+9JOwx02JIxBClY6fgEUx8QanRfVE3vnSSeiL6
vnY+YifG4ppUfFDHAQsyxTtsvai3a1GLO8hbiULVle/9hFbmhkUBXqfXXdypr1f/lgOPzZQv3Gz1
VaprymFtOas1ThbOOWuA4qf0ac+5M34cJ4VSEG7GPS3kKmhnqZGT59LqJTK3hE3iL6bPR5ib3B4j
4XbF6fnajSDscbtFliVwVLe/+BWDbKH0vpa4H18nQG4cLGsIRGeuwwWknKNCODmXBCqA8fzT3AH0
2GN1MNXk48dyGKp5UOfxUh2fpnqCmNLY0ofc+ypx8GVuLNoKI+O7D2aSYai7P5Jo/1qEsgGCdBVL
UKCTMQTIKlRJZQbqMrkwHHMI6LOLvIILEoowuYFR4cUqbmyZfsvIgLUpXOxi8m0InFYk3j5bQ/4N
NeGAGeaGL1JU0qRyq6aK4Fgsz03qlunq97iy3iHWuQdlBH7Im4uwkCG8w4pW3NOETkqWaMvhF9HI
guPYRpm50n1w+Rs0syx0XHGGVdwCLD8NjI6BbgV0G5XPcL3ziODWkARw4Tt+iPAbjXIXsFUDRUjH
6oICyT9BBysvIMt9ulqz0do9wQDX/bk/VojXDCJtodh2B6a7uPlU7oxfYlwq4mL6oam1vwueF3BR
bffe1veAyF/9+U5nrDLyyk1rBNxLdf6XA0pFh+BvO55FIhefm6/vV/IuvXTG094H7uRN0Uubp98M
PcQ2l2kZYgtIBC9q86jPWAQr1K5tMCuAnJdDzdtNITUIeATETwAkU3PVOVpUrrwtMM9aU9ZyiOMX
AgIQo3Br6d2B6A6XEeFePCd7iAt3DxFhnNb99AVlpVjqHAKMBkZty29D+tHcJoXAma9w1wabPAq8
YnfmSQbHXiw8NLqCKTeO+0C9TYL7tlpfgldZPlxM1caVCp/Xba65l46y29+S9PWW6+h0PqkfMxvT
IBPGgfR4CWLw/J2Y5dzJ25neZQkTVWeGwoqN6mVd7+q+CM2MGlvzvx9Uh6wCacKlMjC8DLiP5w76
4Wd89WPAotZ9vGtUlHs8jH/YiQujOr9U5cwAksWKSHkvHdfqkdE7h/ZdqhmDRskhU8uSZJN0JarN
dF8yPiypA02O5t8ylnJqB+eIW4JqMdjeaewAQJMhfNFXL9mOj/fVx1VK42BcjVGhGGhA9c7V48ad
lQdA8fVmHTDo133w4JBhZpxzzC8RMlNHbF2JBlJaYaC+m8V5FOMsE6YlL8ePLAZUMZF9fGcnO5FQ
v0UMuKpKUNCzv4nz4UV5MiWeJilNca9pGOcdoGLlndXdp7pw16VBr9ATNE8zlWb6k76igUQTpPlq
qNwq1raP/ceU2B0oxhWevT7OD/l9IgYx92Zxy99PbDVASzWzcPw0OADTPVItCGj+1BR/oq7ahBSK
3jhWVeTZ5Z8De7HvrQJW64jbGnmWXMgKxRsrXG+HI4OyeDkLpsOoaDWbhe/e90DNTN5YUqBut47g
bgNlgHmDK4PjxnOkZUraBI44A3mmEdWLM1oUxytKzmbQ9v7kSKlIxf7QVeb0TiCtv8kS5wa8VkAV
tsmFHRYHxCNicK0l3+GwzbTMQ7ZCHPREtsAylgvmHCLC2Nn03QDmpxxjO6WRAdZwvXgu/vP+XY2L
N2JJ9hFYe+M6CvHoNlkra9jPsiTncxwd/ROifFBtK6vqIqxktXTT4jLVmYoVavRD7uuIkKC7PcWZ
XLXMOgeYG7ffPWEHFTMozroMpCdVRT35tytzSoKk7AhfIus+0EJjwJTc8zOu/+moNJD0Ody+uXhn
9E/G3eQRTjVolbHMDmPPrhRdBztnyvZhGjog8N3VbMCBqjPisypFH/RUH8ZGwrk5ikSwDA48zVHS
EO+5rbO/H1c6D2OvWJiaoHX0qOmUTfzSNB+WEWcWs877OpldJL6896uyxmzbW7A0F274D1JxWUZK
jCjVzOTaHJH7J4rZ+xxzzZYgVERT/7XllyZujXcQMbca4o19GpSPJS/ypYHZefdqo45XyTIzb5zA
+e8wVt3r1N73yM+kVrG7ymJi8g3xuhyCcEQo8mwrw48dS3itYvX5aT9TdPzQcawbOn3KcCtWLMbW
WKUWo91z3zDES2xH5L6NXS+NJ/pTKpeEl/n+6d4UeIRN0cvJlePt6g1mBBqTmijRjgjauswAMYor
z6drxjKv4bnL31EXx1vaAX8aKRyLt4/zNpWhwGwjEuaZernsr2F1+PuYCcja1LvSvUluhKsAtnea
wu/68WiaozdBYJs6kIen6EV8pTqBygRJB0PrcBt6XEEvB2/2RqaZ777u+nhuwCklN4k+EOqYVK45
1YytB6AJ10EVd27VtbsIxhm5CJh116KLJwRbJ/eABnXwF54cVfZd+a5kDjGD9+28bF1GDnLXzvGJ
XklFV1tz9/6xDY4qzx01fNzAABJ4hXxvYoQsbGhjc+tSlCqmqpgfbEwdzgYv64+hWRz8L7a9+LVd
BSiPwgjJO6co98AbTBmyjt415ajzl0c/xMkFFYftmLXNKjrBHxBsHI2k8qU+Y7+pJcJ3aRll43n/
zu22tnp+h+OZc/BEXtpEvDTF7FXOdkHRZg79Qn/2qVpHVjeuACeilwJ1rX8qbkeSI40zn9D8Rqb5
ik9+pHKiTod6HpGbaT0n2CzbNlNy145pThp47kV7mqaxVsk3bpiuUx7f7B/JzlX/bi1fepiatIG5
m6lIn2/Ok5MZOZnQVKLTlge99rDe0EVCr5Mt5YFRpufH6EqHGBoCGbO1u+IKOKg+bMwG1ju2hWFz
vQqNZBy4bt+KyS8e8WmqXL/fJWT03Iy1AJ7GXUNxeQN1z4vjceBfN85vL8cExxkdjFZh3PI1McjR
Kk+K9+Sg4o1NjAjRQwt++A3ZgmYEHUTh4JO2aZUbwL6bB5ceMXSDC1pnowV504znWyQcqMTgu2Wv
BD4OZob6xLjw7y8WY7QAUq0W/f6OzeGv9OMoDt45WUORkIGaKBeL0ZQcaN2B45HqVSVNOxfclCnn
HYK0Ehl0LFoKc1SObAO61XUE0/0tvXbYL/6wgE+6F+JBOPxkmhg0qYh7o9op7AcQLqDcCkP1Uko4
tssyLq2xg0aOL45qrJup3YqYPWWHOz180miXtl1V1m2vYrAkT5v3M+md+sa++Seb8LLPu8tf3UPK
wSv345GbGIctJJkPVdnyTMgPrUiR+WgFP+QY1Y/DXsaOg6WVoOifOYTaIcQTZRpP3Bn9CYtpBrPp
T04bta8B2Z6P2eRxhP3e2Bo1KlSEy5iztvxmY0JXJu3zdsB4v3RXqxeeO28gcj18SK0/+7h8g+L8
zUCvsWVswGGYRmF7A1ZJrf0R7IvfFG7YYdvzAHSMYfvAXBVY1po7bvIlz86Li7y3LozdUB1mlMYv
GMwFhUuYfakc0obuZXV09U1X7EUWFRl0i+68IBkg+xDxUAWSJLNIr6BCTfFt3DU/GTw647k03MVP
3CxqLRMPaG9s+uJtjDI/MyXLS2DwSZY/1D5k1TbphN2csvn4+ZqsdV3euoUEqkMUOYpONB/QTj5t
F5MSDnCAzN/gPGZDS7ny72GR4DEx6m1K+68rs9JFXo9M1+XBhBTzCFzk8tDgQYl2m33DuAbhAqxV
MAAKehzDcN7M/Zbumf5oOfxs7TltyBFrSMzN7HSN5bUivwytiWsze/PhHH5n8tDHKfn0NQ6273N3
jK3B5sySyzTIc+BADUNHN1wsIECDlXzZ0QFdS72gxD2y9mSgcppjYGTUm6c7NU90PXGT7iqYrySt
Ne94Z7Gn6rdg055oLcav8J7NeS/9ygJC03OEd6jhq9VlNYEfTDQdKiS0UXSCD63ZeKGwHwlmt3OC
L9SdSOB+f4/fh5A0FHggaT9674zvL/JxH6in/HytgkqKpWZrN023jTbjM/I8dk/2uj9PMC7ODKAW
qNRtvQiwfJ+KLQnT9mxhl3EC76mVilfAmwQMgkg34C3pOOJdwE95QAoKBvjDrX4tizyR/7PCMMHs
a/kVH0/CIlpFSSX0L0qn+x+0S81b9WygEANmUDra5662ufWGJW3fqPXxdVJtsGCzHUwRnNphB60n
4Zyxolm4ZOmEV2/beHBQN9KJ/7wWMcPs3WP5eznaw8JJxbJG7lXlawTdIbajyUQmQzlNO0LdUAqR
MIU9Kiak/Ls8Dzr0Uwb6yOZMRPd9Nrztly+Wh7cFhlLUcvW9WP7lZTCIWSdAqIlHfVe7yuBBIjX9
bPobUkaS+9mFbcvql5UOwDoCBX+eKp0pFlAwfl69eGsPJ70/ZcZPZ919fFethlvQZDq0aE3c8AFo
0hI0ZQhsZ/DY4VginS9GI6IKeKAujCIw+aq3af/iOETt2FATwBtgVZGA7PiipwVKFqDO6L53G2Aw
H+7o/URv74OXKONMPD/6DmjHKLJ+Ia+0jdoI1gcV3tZ17JqXwKjDo9XJFNLdzSyiMYMaSN988pwX
btbl3ahSjQdIHqOkrMXNy2i5lqz/1x9BW7yTUWUrUAMiHTDHlsoecG0zsyhhlMebwgvoPV35ZAAt
qUEz3zRhHRvFXiy15yY3cmqTO2Yb/TEnLkU63rkrKMaWqTqCtOcI/DBjjuOmqHHHnNswptqtU9E9
EhnrKf/5SBvoqV9RLpxRisAuKGyazyFVEgY31rEQe2wyerM6cmicFEJylsa8lt1AWHnqoFmOA24n
omusayucV4mCqXYCWCrEf0xjd47uMhH1uGFdAutlkqT2PokK8y03wP7cspclprkG6dzssuNewbLw
8Izw8deepgny8PzUp7j4Bob2GI+uVCrFQZsLLvugfDw5bVEQIqOX8/3FaOfAVM9vl5LJvQ1kSXtA
s+X5THYOudaTZbWL74LXxcTqgLXZtsmhgVhsGbzvftlA7SQKimIuds2PGHVhUaBjxdmT9PEgXraz
vFb1GU3w5wzAB9RXPriefY/oWMv7gc2YRH98s4cteDo0oa4WNuBDIg8PTH99rBiIKhRWXJBWGPv6
0mxOyo20jg+rvNaWnJS9yn57s4KiEQTBR96sS32nBxML+HoznVEBbuOourSl3YyjrDzP+aB8oE+a
8q7v/3Cz6WJpfaqGtmf4Fws+YZPOTgQhQ+QTqJMnFnrHWZDha9Vn/WgMi/7zfQ3gMh5wb1g48mLU
hK5jyBrgN1KwP8ak7ru8ca6/uk2yAoHk6KvyK9yqHR6L4drUIhk8cYG1uWREKiIk+OrUS/ftUaNc
3jQQGBOTxVwUMQ04i8AY5MhZuNdA5nWg9EEDZLATT2l5/yo0Ta4eXkdc6qEIiXmwL0airBVZAQSy
oYb3Zy0hQ84k4xJjcOuJ5noPFp6tOMVbMg1U8DbMXm9U8q7D3blgr7MlW20PsfCN+EyKlzvRjeY6
MzrOfl3H3PocEjzAZOuY3YCx9zjl1ygRNeLESD5cgEESf6bNrDuJ1e5EF/n/7gisxsT411kBP/dt
QUmht3w1bOrmGtYx5BlFu9JzZfh+tlS8nd1YHEAFhcKcqj5U7cXmcotBOHxVKB9wjxH8Hg9QjzQM
txM77MvqxxaNBgZM1Vk5Uwc3b2M74ZrgIDW6cvKTS3oKLMDTZfddw9XGYHsh6JcdANgIbJFKTb+D
2qS+MLdFgW+UFRDuOEUMwgeqH07M7hMSu9ksZxAHQNc+FbGTPU1scnHoGhFzhoMrYt+pYyI4JMSr
YYkOPBnTyXQdHMlT769/V8wG+/dXLap0+XjeA95w3tKjKwhQMmt1pEsOtt4w+fTe7/Gd6jlm1tEK
fxAwADjw677mPbsW07C+132qXViOgSmJdg+042R00CPBBIFSmNaMA7+hscCNOUlRPvUAyCgrOmTl
+/WI34EwVTsH956+TIKFyntdAHrDrsKaJpByGgGyOokJpJVfhNAFfazYsTbZdhDdVIjA0fWbp5CI
kW52uCQ/cxaZn7/7QyCDsznEd+HHFSe0g72JekKDlJOCnK5b+NO2KBDz8xcZtAK96X/PpEHWFOYx
uvQcmNGlenzKleaD/d7R5c3SvxR8FKxEcRYzm3pShuTlREZ4exfz3uL3GDgitPxOPcjJgdi/3RbL
2enR+EIfS80QvDGaa5O/xrVpSrx3HrX9wvLuzv354EVSqoXW5YRMJh40F085SS7+3FjWFXjLD2J0
CKvIqaH5wgUdQJR6siG4bn4RqlP3Ja+oXgOcrJFMcNIr5dwuSd1fGm7uzLW+ykWvK1gGT45Lq2Zt
O8CZUw44MxHDyO0fPAoXt3Z4UBvOVJFQZvXDiMUdhbB2whkqhtfMbhiS2+PUHq6+LV+QckSbFlrJ
se6Xj2cDT+bM9l57I16d0WHdXdK9pYGnF7zyHy6wDeQoc4NL5tl4usTihKabTYfnknuvZJ1cvqfj
gjCm3btkNtjMFRqfCRsXCbQkVB50PrsscjyAouOoFXhq731gpCYK0hizgNzp1rC7sgyZnLsv4RVI
9vbB//tBTO4F9gBCLHcAaZ+EU7drEAg8fqEyPStKXnXZKNk5jSYtuZdPYJMsEIBPFV68tEStyIwT
9nwa+KDv+j7hBVOQ0GZQfAWf8HmigMcz7+9YLplTwjBDlv1sDCLymhEpLgP3ef9w1ILJRHVawdPy
Ye8F7cszhnCi4CEYOEOJSVSZkGa0R70LM4QwzcoJuo9ftWXTYMAsALOycrGP9rs4zIwvE7IvrD+x
8xkIqBl8dJthUTyPnUUsODPxx/kFCNQlTyiyfyMFyyW3ZG+unnEkc239APapbdRCdeoj0uoxvNHY
9Ga6L7iWiaq4+waB12WG+ZKwroPS+U/SbdMCp/b6BpuHHsQLMk5s+CTZz9TI74NUGqJcVLIIcfRt
CEYZvrMOHtZlXsbyzCEKphUw/nDVS2zO+P0323XMlaFnYjZTU2yjfVLezfkdgx1eXzKiRxYm4PXE
hjeaCiVkozl0muMxXg8So1WzHBsLWpLZ/N/pwpBXGhI9GHN6Ech4spwVTcZULqfHFZUATjt5HObI
4KsY7yeky19kOkfFWn+e3iZv8PCnhDYsdSFywDUW2Nii8bfH0Iisr9PGFJG5dMXRbmuSbsn6R0FS
9iklYzQj5YMSw/0B6lBYltVfpWNZ88VWvR1OLIwsjKzn4wk2BszwZk5nsXSA1xWh72EuDgBfgwFo
AXOi6OP9rYQstRzkBUU4oAelGux3Ig+INxOs6u/ny+aFVA+b35yp2FTF+fLzE8BeywClmNa8RTQX
0voXG0NFo6mDHXX7GYIS4VXg5ytC6ZpLrLsrutH/IGvaZOqYZxItPddTpt13sL8gpB4YBa+ckAcx
qnkIHbVzuAzIAqERNp+8stbzdx48VKwpDBt0f4KXBwJaLwLwdBAZXrOOST1uzg+OWB133HOQYuj/
6b5Z0/EYzNsL5XEga/v/maHC089SNXjIBBeSNRQnMzbNTAoEYC4vuF0jY45TjrhZPB8gqBNr+Z/v
1wdpkWEQ11bYtDsWT2EOIjX9SsvVuiPMUcROASuzZqy9LwUhSBIeDVcgF69BUMFWm0GWXs4mFpln
1PVyQ04u8gHcwo1Dp4b77EAlHHcbtzdN8iVv5CJcOy5YKcWqxIqQVafZ7DMevcQ4Y+VdurOEcJN7
FwSHUdmTXZzm0UuIL3dcylVSag5K4VlVf4ndrrxbQrMfXrRohpg6fLeZifBX/o4eUSzbNvCml0nY
edlv1tO1gyJPKLe2RDz6Goma5cWey7wxZHK5T/ZFNaMVE+hGbv8Q4QWLBj2dXa3V+xR7DVd9uGPA
nezT2GHoRsZlVsGvh4DmoF4v2pn1LgAjcxbgg9Xe5x6eJ/fx4A34a4/gimS7ND097EPv3PqQwgHl
o0iq4yVKTrk/JEpM0+SvgNS/PFkB1LD03p2GA1hXzt7An6lZ8bMWkMMPv+HoYGE0bDcaic0dj06D
srm34AXcT94ld2cM1YCB2lmzNNxyGWAWDtyMd03d0zCV+xJOQc2BCNFsyQWRt0q52K2DJtxQkgrk
y14kSTLHKu6miC3CsY4p7zr5A570Nu4US98G8qzVYVtFv460b0EWcFeArObF29Hertcpx2z4ghvM
OTfR61uUcPyl5GVA4OvQGJZCvOfJUOnqEKeF1Zzp766UxKPiMi+KwOj/BEJfb2rxMic8caFEoKfJ
sbY9ANTejKkLsdUduulheyYOo34cjAQyKTCpBgw6jxC7MtWmdWYvLWUj51p5w6PYnJ14ecOrkV4F
Jg0hs/YLVxf+foRFMkBbbzZH3zVkawGLvxokKQLjnUzoL9Su/bHfVxVop2n8pgsQcYRZT98A2bW+
4JXQ0b4iGtdhj9uZMlbDHvpuiXJnp0kaE2Ln/JfNv3RadGsR838He4AH4ae5p0dvA3mTR5TKUYyl
Mnz7VCfnW6by5KSwkafoD9wNdJ1NnlY2phtMBhQPv8IElbnpzMwLIs8f8nf5S3/cpQP7rE+bGR2e
VGqwosAnTAcfRT4FjF6TPtjdYYjnlZdjCtrJHifFD7p/EMD3rjrqd50MXZ90y5Xfw1Rw5RxQRIKF
82Q1r8/GESMDTSxCk+rAA44+POka0IStEJeGLNUWMSwk2DQ9nyhViN7diKFqqKe1x/XqeUelwIeG
M2+LEuXB2w9rt0JtAW1uPvhgKQ7xMHpUErV9XgN640qAR79sD8N5fepLQp/kUVcJXptZwsfFVJq8
w2HWMFS3HxWECiWDCSVBG1+hJrzlf+W6T6xYh7uyXjKb2HT/omA2JwJkl1Pd5BfIUGpQC418Crxj
XiT88CY5RtvwS2uSpDMaGCLO2xYggWGhwsPwIpnFormpy6XJqvGw6RxvbE9NrQ6Dobg0vjja99Kq
XV3Mze48EjTQVK+pMyVkJnZnenNC3/LIlRToDeUwsferxrVn9EK8xmEOUYbrZts510XK/UBA8uot
3wCfEkJavWu0MKlCPUmUaX5+an0Z65AqRHhAkczZVDGly4GnCqkw2loUuLoGZeUtfpMnmBiet1dQ
HJZLO2pfW/ZLyibi83MD8SsAbcDaig66RfAFabqz4mZgXKBWojev5MquIu/Fd2Oej3Fc0jKaz7y1
1/eeNCtc5lL8uIVxMC/CI+08s9Uq4hZuzm3Pns1/uHQ06MrxJiudIJ6mI5BIMm6JGdc/rpE3LRxx
mwIqaYUdJ6uVcSxtolQl++cH8y/1yhko9EG5ttmNQum4C70bVNEb9nz6Zwvo0fcx6r/VagOEKbF+
6oeiwIoBj4Xoh5MMDGViu5e53tyqaUDKUDnfgSmDkuXEHwicHKu9kdlERapMUbvEHyOFrPXyUHs7
dX6Yrms7OV+vrAIjCZhMNdShuH1ylFzJxTiPSGLMlT/xOAyKJ9aVTkISNGP7l66E+yQeJwYEp0GO
eICflW3PPi4HUPYwiTLOKl3+vbk52hr0CXa1lrrPoHV2L9/PtUovVOmNH1YwVAv6nQhj+Aq0tcJu
fWZHskwe0SPw/MODTFzGvKRMXyHD22HJz81dhf8TigF+U1NRrshEsu7+nz4C8dCPXiMfrYEKigTs
9yXRiN21xnd1Q8jUm1nGogKpieZ4QgNAROXKym0mOVVY4GkKnQ8LKIbzf5BpniIgcSVFEOBG4w4h
+U1TRNrcsCEW//KMRzX4saZYFfo49hDzDWRWBdgaTGO4kvYsN2K0zj4XVXhJmd0mWl5tclWdogPy
MaC8XLAixA1e8mNf5aNxDEvmBgwGsPVLkOfx/tkZ+ehD/QTomRyvQ8LRrScDcqG11gQWWXmwjMD/
Xyq7NdbXKvcr+/vHfSFyRw7QJEqGX/M/ciJE0qLNbP3EzJztoidPCmOYCFo5pt5ZJxrt1dt/MMhi
XibiDZtPR79wySLL9DxdzMQGcKMpGhbIRkYDMcpk5ro1vGK1zZXR1ntf6z3varNA6KrSLiHO4MML
47rBFuqYKy6+IWQCFGO7oZ1cmkLsltH++u4zrXFZ58Akjd9VZzmXUY/S82gkrB7ZjDnyvPizHez2
K41UN2A19BdeTNr4IcqM99GCbSLngV3tsJODOnpos7gExyfLhkkhv5p45fIrNzlaIxa+fzmhBjuK
tX0cYMw270l3BXRowcKaSNOpCB5ajGsvrgWJOHRykAmifBKjEg4z4sDnGj55Xxwq4fZ6sMEVxDtE
NCI0ThCYzVrlIT+G/h8pa4Dxz7+ogWVmgMN4n2+cuRej3H31xhLVsPjtiQS4Neoqd3ta+hv4E5Qq
yjrs8TapwRTxjlFBiCXmWM+vMe/tSj/bfAYFGvSgQ83ew7f5IAReyr37Lx5uhsCKCbxKGErlCpEC
KrlRiQJLPFtUSNdoGvcCEiEEBPTVx5+23B59+A23kaXFNcPbqkvi97nLjhuZT7nVeQP+kEwEDvmK
sJlr9LHnNv9vEUj842NPTkAVNZFw2r4e7FGBjnTWbixm/KxgwX6I9cAUQ/zrn7xWd5apCMlNGtd1
DI7z3bsCy0PKP+dkXF9w43Utwbm+uYbxmMqPxja75RiWDcm7O5kLe2b8SO6OAUSk9nu7ZPenwXUo
sb1+V03Q/jXsD2IxFlldYshlS94ZtavUln83+STh4fCKo2aXXwHo4NyIQGvO/tA8dpIGh3WjGxS+
yKTc4LZ6KMmfdt47yHPlPlUO1zoFFS46mQXOgupcJEq7AV4aKdFyJ7sLSNYIm9KMmdaeR0P3LjAS
AYtMgPxxF/VaIdoGjlOiBu5bax2NrvhU4wkIQUFq1HcLcHvuYO6IRmwX/NwH66R9KK4wRsbYOwUc
9ousWsnhOeXvQFXn2Dr24uLrfRF+b9o3WBcB0Hq0SbJRZrWzjmUKsSmQR6/Bk91e9JMGlkaxjqz4
/GX3SbTBTAV0gqjflRXNRQHwewUOttHarbYcJ24zOx4lm+rsEfgPmn5Rw/+vmVRSx9tyeAn1LAmV
ho3MBlwy82GGE+x6fpJ36XAWskGAS/rCr9jsLFRfbaiZpvUDav8wlPSM+w7Bk4pISCE+d7RyHXc9
qLGtNqgjxdRjHKGl+TYrOtIB29iLVvOLmUY5bhyaQkTlYSa7tzvkhoN5lVCxRSL2TqzQ0HSOYNDQ
o9iR+Qh/9UxvxhFHRJuOU120nOhXvPPBhoF5k+PWYRtFimtyAGBIewrprFoZkFK57RJU+2kWaiIN
yvjt4fGkQkiYmehqE1AQzW4q4Q2qnTzSaCoB3HfB58UsmLxikFiBM7yz+oLwi2XDkh2Zee47l+pW
8p1QjJbAWg1ZxmSFAJgj5nvrZn/4qw2ljaA4nsAmLo9gpZc2gLt4P7aUG2/8HKHbrttqR5XZlvpV
5GOSYR0FRMU5fQ6kol9dCpi8kKu8xsOrLvM745tMrOLz9AaCvcT2W0T1yc4TK5DwsVgsDvAaPVHz
br9IAn0T5yCKtVeuC09p8W2LmPb+47yjoevP0WgAvO9oaBYJwMhEubl13Cv5w9cXnu2ofXxq8mvS
N8TtYiGUrDRXMCPYDpCYCayLsFL+72kj90lO1wQpYpuKVh2xReWI8LPe7T3JQCg1KgVOy3TVNKom
mgX0nPPjNQQUHAsymph5uuHqRxtKF5y82aEuC8NJfDWlA8WjczgLWRrnjfRNTva/vAuc7CdF7MVr
VlAzZkdw5fW+1GRs1Lu7c9u9jSMc8chA2y6CUgKw51PWEsGop4rvfJ+YijU7MVpoCS+pGOZMKY1j
TAErSCIj224RUndGYcnaKTVcVTcvngwoQ8yTMijYmhPcd7RjOLQxgVqrl0KnDdHeY5nJVuRlemXX
3MVcZ9yhYUlugLuE2DupfBGK0LLrwMOk8fpdxB8T9NPceMcxnaSaiLYvyIIRb6Z5vEHJS3Tg/ZpA
czy8nPZCiZXxJZeNQxcu0Z8aT70VWXfMU9lkVSB/fM2MjaguC39R6ywX8yTUwloTqv0T5weOmOrK
+rbfIbCSROL6Yj8fEYvmZ0j+3hbDwQ39e9+dmHV5n5LW6RxEiGUC1khnH8rdLsoD0KfUlzJRBCLK
IL9TOoirrSQtDYQAZOcI0vCMlSREorYt49wlJWlc1uIHzJ1+D5sU3akEfP/8mmwCFlGZl/UuY77D
IBSkh4iuBrLFkizY3FMXL3HpO1Fyu0vdqH3qnI5jlyTklQ8NqUB5vQEO3X7uknPT0qzo7T+UROpj
V5WyeXsYPpZM8HSxf+QPbXlcgOlhPcj+60dIBXZOvOglqO13UYcKSdK1rRyfgRpeyrxKnhjhEp2+
kf7RUqKqIdNG0Q3SWbGkYzM8INfa5FPv56JuY/pq0LavhjtASGVVpgczlb7kxZ+z4rf4twAjr7uD
HlyXXcgWhdTFc77b034DFXT4NROxJf21tBiTPN0qYp32V1A5A+Bf5wqS/onjDaumO9xgT2URkRn3
hbRGQdqGnYBvN6YwShjenBjNUIG8EULBqIxn21s3LbspMd0mWYb+Cdsn2ZIGvY4/CrpJVbyqVBDu
aZZoIwzsOLJA/T6zasewyv210yDZM/O9noY/YVCz8Y1WD2/4TF6B5ueb/hI+fsmbl9qXtRdNvVZ/
+J3G6jfy/7OSVcepveBKuCdXSs98c0bo1x7itToMV0b/O5vXtd18Vg8nIFCuZ03RiIe5aw0grv+9
X8dnw1vYgcYgJRTZdMA6LzF6tjWg+MyM9DTk37PolX6bwc5qbdkaozPv5PFfowal6ga9tQX3xu+Q
9kkhfXFhIS5h64wYdvmo9D6YzBqTryZ33nG2mLUZLzrnve6fE5hLRTbfkf2Fl+Mh9BZ0gCjWvZs6
QFfoAa+M6F8s26sZLtefb8H16DlxBzl5gLgPfD28voEuZU2cx/uunXrnyMb8N28lmS8pCWq8OXdc
8umtrtyVPTwBl4DbEe4G5K7VTNaczMQ+UFJtccF39MqWRC6w+FWpU1aBmn8WKE/dPvJOaQZNOU7b
A39Tu+PKFMP5I/z63myeqWJwTIBQYMT327blzVZgAXlBkyYS5/I4IVibFoheaBw8XyVfh95/5yFN
ZNH1pyR55thAexTO1Uv+BnzI/nFy6nG4BJ//wrvX1a35OZP8lFMiYdY1HuT3jfqr6o3O9pW15wiq
af+cB5k3JLCrlD1R58ScpRAnQ6UWVD8xWAg8G0SV7y1O1gBn/WCXk1c/4AJNT9DTgFPfCfIc4MiP
TDKv77qZ5BUy0z8KlzaS7VDowBniiV/bcEsiXqsZp7IwzdkqDg3VGclqnl4psi9xm+LIKh1+9KTt
6cbRmVW5YaUgH7kfsxB0iGpzUScc1YCqdVDaggObVOqPWZ6YNM3l8jiECMhmfiLsVWDg1+RY8GNc
vgFoDlbVUhM1CQrTEnjLonhM+TKvOhYR2Lh7qHYmi3y6fhjg9uYlGgu0m6FC0GvsXZeA5qGUOeHU
B7nWtO7n98jQ2Bshy+K5g+Kv9yYF8aUBT1FeIWzdj2hnOuby0ShF9WhRFkAtex6YZfhBQYArdNcP
XxqWivzYOouiMCo8R+cVKNrVhEcJcoCTOUox4ACUnTGOF7r0z5AlH8DpoomUJ2y+T/BvASxGmbYm
cwCd/0RMFetEopyIDA0+v4m7yXYIIROidqpaUrPSTSw02uemzkYHglbVERBs5eMXn/Nxw0a3PHIj
Z76oIX0vMS72GGuYK65YZDn4vjXGeziJMhTgDcCbw0lNRT+7nfFIMaIXdTbl+Pz67gxr3ZDi496D
1V9XljI8xTrvmE9bjexkYQMtIDW5HmCn++EIbQW0GPJ6x1HY79DYpxBGbSeETOUJh7tIKjYwQXOx
+nwX1H5lg8cNJCIcxwKAsxCCgh2F75mQnE1V4WQDi5db1TU1tu04sx+GoYQeAE1WB0oWACcw9cjF
PYH0ifHUun9T8HpOf/3QhHHOp3O9pTyjxVGsUiSD9HEZVyv0ZJWb13nLigWGv3HOCDebzC/xhxwK
F26YuAu/k52IoSqlALHfAfXIYZaArTVCbiG6kITe0QXTY7n/8xiJF3UkZ01XCkAUpA0z0nkY7mnM
UmcPJnrUbIlOtLiQyxbmqy9pqfGIq6vciCt8yTpoQNLnWdZdpWXIlYTcSVpbi6tFPYAoIz92+Klk
arhzbEZ9YfrXDIwizNCwz87B5UlOa91z7EvNiJ9DSRL5rHkX2mlZ9uCPQzclInHNnds+AIxtrMtL
290057L5kgEEpRIb01ty1qzfnH2z6k9Q8gppIBkU4ng+7WOQTOrmC4n9L9y1+5fRBUD54qPkeMXi
JkDXFCm4GncacS0ZkQ3xFkfH5WkcTHu7sdimQRmajEhGOW+6TNxhtBfHmQmd5HMwSoSCd8i2wAbX
ZKJ4McrC5NdOrNEvgXHFbkwQb5laO/JcfU3UqhWtqiAw/olK7o51y8OFW3hxQNDH1DYNsbFYZhjc
H36U2e2P2vLgMsfapfX0NSLLWAB2Er/xut1NB65/dHZWpu9DjNVqdZiDOjco5oUfDSv/3oUlk43f
lD/uz749jcezajMaEvaPQmgs85f2jduRE6BMSfjT6hyA6oT3CkaxUJ25krJduEUaMj036qbR2MgW
aUyZvN4PCXCZ75b6If+5kg0AWVEShHIGq4KaVUGBqeHz71f1ma+Hvz1oJzb5LbGpgk0Ax29hpxoY
YVWYxyxMDM941j1NZaCjROQ7etxa1kbrNGMWWkS89F8GDGgnPqwELTHGIDiGj/31DN6/UIYsKXSc
a3GoMfNrqszEc3BxXacMY1gYJPsNTW0K7bkwFg4vIWDWDB9uH+W0PNvqiWQyfZeu54jGBc0SlN8B
tKIRvxCxT2A7VotE5wVGwHk/FBrGP0guKBl3/GxM/OqCsb3l394HXtcDjCYg3iBYTQ18SbZalerm
3En6MTBUpX25xb6J2vM5PRDP3ctyF5M1isudy/SiKOr7b/F004HevJxsxi9kqwaowLcOd7xWHQz2
DRYugvS8ze3sseiz2R+IiWYKeSAXl0r25saY+7W3fGme4S4SWqGymEUF2osP45oW+SwHL9EbxYPX
WHndEwFs5Zik5hbeyozmgsahzcUjxvx4ZdIpUWHnXgZbTlL5HbSI5ZJE9RnurSnDvbvokQcgiTiJ
Oa4BNNa/AS2d5q01eLtEgBfDNHl0ddQdCZ4HNE7m0c1sIrJnnUZuW979K6GBNYhTAGkmwByAiCqe
6Qqt0ef7m9CI0Q5Ls9L5Q8RIBGws1f55Cv5Ghkvtr2FH7tTTzGOijD0c2lIk5MsbgGG2+KcYK5hO
xJRWF25qcSrh1dbI8d7p4yrFxJ1RWyn8CMdban3jE32liC+C4BvhMlkym7fN8WBgRvbA7+nYF2EA
3x29Yfd2wwpZac8sViVwvBuzOMghq/CzCtN3p1zs5Pp1pxy+a4vOgXctNADKwfjL0PkFM0fWL86n
3VDnbysnV2YQcBVbxjKVf3a4dRsHPdYmrkWckGOer3hlVNjQtFI8TEWX0XL6U7PsuISiPx69Xz9Z
4cGTWr2xM3INxh1Cvh8vSsOHEnA/H7Py/XO2GbDU4+qUzLApOOvSVbTEOlGZywBHf6PmSEu5q0bP
ESunDXPkp7+HOSn0XKCg+/E9vg4jSjl7o5mv4bLbG2CxuQB0u3taR9jHIY3mr2nLiqxfzTenN4ks
FN6jAl3HNZkDMYHb3i1oBJsf7c6lenY0j7F4a2DIhkwl7AmAE9i4hFUpT78B+lX3wJG8Lrj4P070
wSxke3MfZ1ptUdoD/429e+RZN4aMmF/hdFenNg60THT+6ZX1ULiBiW8CxspscoPF8YaX4XoQbLtJ
UCK2WeaAR0KbMSP79RSSIJYX5NwmogHMAph3JrsUdJPoTg5BmHOjwjZyimhwvKjbQxQtVVlUt0aT
KdnbW9Dc+89MJ3LzCtAA/A1uoAQUjEXWeKNtPCfldP57lGtWZ2dvwFSb/xEn7P3fla1XuRu4zpla
lrzqTILjUeRwSLM/ZkD1VQgfXfkgzqLqwY3HQk1/RjuLhIiyLx5BaPDi7DsmbZHJwe9CrM7ZDpYr
75GG8s0awVeIV8N7XXM/F3Az2bqWyjhmx66BprWT+qa0pqWep2/LQn2esnxKXDvP36brgswHQ5MB
st6X4OOjJDB76rO7QbmCFw1cElB6j+0bQjpQN5/XAIU7eggZKjWRtGdLfZNLK8TtUleDGYbJYgyx
u1+uFAsOSchLkdWr899X/ogn8ffVmj9RF6lQQkg3+IqxR1eh+xm783zxuE+XWBgetSW8wCpcsZOt
9sJyFCq9e+x0YYFWwi+tFqaFDBz89ZGz3FNn+QUOJHMXLXLqvjHuI6W0nY9ZV0AHgFqB8t1m0hlG
+vgR8PdHX4VIm1/bvq0rSyh0C0CAQcuQMU/bpzcZHgjgqhWE+NGSaiZeaNMv+dzGA4vhE367wWZX
timMyr/KT0U31RCtqWS/PK9RB0XmKuOMYFVtonKhSyUPdYzKsyHK2Jp/DMR9bBfEblU3+OkQlYSa
7bLel3EyjcUnvaNLlZe+uzHoCyUds+peuXdAPFBJ93s1kLOMYfegXMsuThr4F2lyCY8mJIzb09Sv
5TJpNlfZXgZrLSckUkHMTgmQjHySKB6HPfHCNMVsNokJoSD3vLVQcf8rmEbNfTaZ6z8eMKeXYmEN
KrR+Hl6/+EXXLrW3mUrQIq0pd0nNcFEGkV8uSBEq6vMvaB3b1wQdD7U4cjSTykeGuu0OCt5VeLrG
wClmflvUYNbRZFXfxHoYQMVcaAQTpKMgNNqS9T6fnHrLXeBsR8gWCGlVTbK5+nL+ykFtS/Fbhpb7
/fHa7DaTM2Td55tmhRie4auhLjZF7wIFuzBWJaOyi9EPuZMWoxkfOEtLS2Ec6n3Y8uCyPa9PWGep
5PZRLjOcq7LOQZbWUuDO9UJVbqQoV5JgWOE+fFaJD3j1PCVQkiMVIsdYrvG2seIG2CgPe0q6q/Km
Rtl6vNsxRf8xwWLz10sWhBXn2YkYrdoooqUS+lnv4+xljwm0uXS0KTCuUKzhNqHXtLo5x0VZqJIj
fHFBi6Yyi0JiP/VBPHeCqdV/E87v2pMwAhLOMYmTr7CGmEyGTFvoIgJ+uFozx8I5BNMwZmfDUL7l
ifA4xArlp15OVTuAXWIwxCfT18s0uR2rGmqQozgln8XWm7vtoLoGuFq2F/ryk+MR2vmHmTfX15Z+
lGZ7DrYLClMBxq07mzJPQ4fDVxCHb+NtZBvCpKCiWjovq9mAC9zrYm+IQ/0OT4OySLZy8n+unSHz
L3HwzbTswQt75z2GZfDXHc6tviWNUMTW0DFl981vI5EhM96L62jAnNYwnCQSsGoFJhffY70aM4if
4htfXjGS6TZgsx3Ls93MEBve6BcWriw/abMc1qr1rb0STIpuwKB9uiMe6zTHG0HLh+/T7lod+cgq
0Sce+k7Jiiin4QQel/NhYT9yiZ5ObRVurW7RXlCR39eU615xhHH7ljQUKJser0DOIvOtnI+Jp+/W
ITMWUg/9uu9YnfK3i95yQpnqoX6fDRCony2AIPavQRcQZmJHCCsUHCwXsxSLYSf+IRyw2dKcj2ck
LqewP+vOwnyFKg/5VKa18/vF1t9Hww5hipmuOT4XwCsfN+Yytoizcv8MIUNoe4Nx1HJbZ3Qoszaq
0m4mbU5ndohrSRlLgruxtIyBP9q0uPWBjyJdIxN6hlcNaiS7w47nRnuvNqqN4pzjxjvfXoDu9KXO
f22UUk0Ntqe7UAnwaxGShstkMBA16jQrOtWNod4MjpnMXScLQY0vG/Uq327B09J76RJCBp7UCNA0
Ox58j/yDbzJqGRd6zPABCpbuuYE2j3yCqjI1mvqEVgr1tvJwGjhwsiXn34DM4TdBrjf6BVWy7Kc+
j3lLtjjIFvG4/378rbnWeFTtTplABjoSOD/kRAE6VdblgN+RVM1lmqlbTWcog5UOhVR9zANaHfXr
cj2EYE2QfW1qRwZvqlJWj3NyBYvbgCnUXaHj2mQB5hQ3lImGZ59B36y0VW2yRjokHdTH9NT0Tk+c
hq5VQY+N7hbBOZTPBaKqHcK0a9Xfqge8tZr7XxKtItK9x5yYnSzKuiMfbKKXkPHlp3X8UYOqcjXe
poVX/BFuNiv65egAu0dmIusFuxSo0yp8ddU13J8YMRpZXh6WdYllIc3MXvGUFXyetyXKlWSVov55
78S/AxKAeOUtt8VbQ2U4ql6dkaDTSdv3Xuaa/6v1exLqcjOJ1nD0/URpShzm3BQtHkF27yAk9Dsc
GLJqrg10EKzoKsrQ5kWTgWoriUPubKxIMflVIEDgdvhd7BG27jUCS1Vu8fLYQyilZpkuSeMqTNQJ
X0w/ZjVYMIgNmJe8w/MwtjaEOAIpX7YJYPSQy+mbUHBu6j+DWChKBQZjVGwonhUcEBXvNOmTu2/r
0eDYrqMemfJhGQEMk5WWXwH84ibgs8UaY1lMVO+sweCaB6aMtzamhCiTm5YiS9sRQ+Paapzy6pah
KzcZPjXT6NqqvHNv+NejKtUrByO7PtdJfxqP2WhC71gkveJRgUlnfhMDLwv1a4SvQWIEAdoBKQUd
piQ+dJma4EFan/Y/LfX9Ms6iVbQoQ8XqgEOL0+LEVmiN0TsSZm2ar0b+IENBJyI/9qwnQU+NUMGK
+oRnGTcirOrqxXF817/KGRs0IIpdbIyx7s2fYJ61H3obFTEjQOUghgJBMiRxZKKLjQNqG+F3xW1c
M/LamWoFyZ2blF8/Xu2AMfdW3ZjDK4BVZDLcN0RC/Upcpp7ee0XXBS/8BBzD7iZ2fVJyCz31VdPT
nMF8zCTt6Yz1BhFv2YJ3t0kTa1SJBx4rtdT2aOUycpwCLA9AL0ZiQ2EjOk/MtsTKuUxAHZ8cHrRz
oPphNxQFXBbBIeiRskwyVSHxNnOsnJfxVraVbgEfAifoCIlKEw+ZUNnQQQOKDiZKsC38HeXMdt+Z
bsErscGrpK+jlVkOhqGwRsrqBEjdW9g1eKGcIlr0neo73o/nAzHhN9NdN9+BDgxf+l8YCwErgDys
yXnnBy7Kk1dnZvcr9/Xwn84e0jqapwt2ovOZ6dNMoudRr1Jm481BOzlbFJ8Dy+vkMp9WnbEMb62c
SBcVSRnoojnyrwNwvq+Z2Uz1LjwupM81EMIGzjEr3FLDdJlUXiNZoAVPK/35e6BT5ZpDZMp38qIY
0OvnFgxFfVOkUPKfGPmBtN/Xz1tDhcfMjH3oZ46stL2wsQ+/1KsrR0jQSR0W5171NSYgNu/4hPE9
j77m/aQtoDwNnResPAVVeKujaegaNrX+kKFRge6EpN/JmUTU31jwRbmKjXsEtLLoOmCqDrdeJuOV
dp/C83pN3nsCOsrtknXOYlJPbnk3s7paCDLYC6Gre+7C5m7wguBVTyX0Do4hUeALHQRuUM0BxjT/
RS5MRlYx1V8k6RINaPa6k+LKzFoWOiBYPV9iVORNy2kCyo7riFyozphHW0vmKIEPISLOuq8UO5Ce
/pORzsk6kWmG86o7jvuHqlMt7sfoQRzhKpkzAfbKb2UWjPZgJVjXaaVhyIF9Rt687zKtCm58+BDT
yGk1VovNRRGlTjGTAyOExdgZK8S+mI9nrd/K5+rDH9nAMoGF5IHiV3PVJkoJcNpGxYK7XG8ds7tg
UIdmXM3AN9rCHcO8eIVR8LKKbFlHVwDRLmnvMB9PkSpzHh8bft9EjXl11JFJgAbbGKGY3SE+0fGj
XNV3LUs0drZbRGdpsdmE2KIj/ibKmS4caLIcfsogv/GJzg/0mYvRj71YEu38FFf6vhTUluSHg1Gw
pq/R1Tv5a6ZF+t0aFRIPBq7tr/HOpKyNILih1k1Eye6/C5cNxb5nhRAFl8Or02i+BESJqCWPSTbG
85xQ1/sSCxHSzcM/Oh2CJMbcqDl7F5AKjcYzq3Qfgfr1gnPZOdhsWIcnOX2/yfaMv7dC3EJdMrTS
sZY/+sbEmpwQznpuGikn9ejxCcL/UTiE7VjDreRQYgfE1x08z+eQ8fg+LOEx1WhhpWdd5WhICGzr
004KlXgrbj9Kj5h0LdcwHqFORuinuhntrXCJ5Kt8EJxlzjpj3BzCNDF6p26ax7midbOMwkGMcqa2
QepR7u8V1/wKGqMSZW+6PSJe6w5pXOLw9XrklUBJeuR2PQdbIEh/KFOjdBX1SpixGCGw9Hr2Y1Fp
/hR3y2rOGI/sz9cFWk8ddjq4kn1Tbm7BoaGOOVc3+Iu9NRPzszmO/TJWiPCkbTNDmTm00SKZKj2S
mAdt9k5SumXDKIid9wSHdKPh9XfarFsCEj29KL0HbZbgvjZTC1uxCD5YApX6Vvi2NEMiZgZwozSD
eoTmPOK0AwDBXzJiEo+WHoywdbLsoPDhwm5BgDg1hoP0AsanV4NDbASk3tooN5ORLDlM8+nb9etl
410D5K4zy2EwMirr5HQPOOvPqByNNtg8L3zxr82N3+q68l1tx4P/qbx/BmLZD8DyR0IoPkLoqluo
xHDEk/g+nNLWRribZc1izOHPiIGPZM5WUje1jZKROJeUDHlUeK8RGpkGRR7iDH8T1axlLt8R8J+v
DBdVpmYJES7yQ2wIh8N6SFlqQaBo4fYvLfU43GM/S3PaF1fUBQLYGKcVgYOqITrR8aMu1Ys4/CDJ
62RVhwG1fXXvokf2V7jhHBdbmmXMwyYJvzZkl/8jXiaPZMTgRXpRnKAcvqEYpBomvv5tX/pzSYH0
6SAbLTNiiwmdHc9itrAJnD5wGrb0M8Q6SmyKDETvQmYnroX8g9Q6PHXVHUaFQh+RrAVpn1S396bW
7siYxn8seygmWyzTs5nCXTwxmuVRMjpjjBXGcYUdt/gGTIDOGxxrqNt03o6NJ5x0ZfBmYvnzsk10
XwmKzVMO1pjiMWadXeHsmOSO8lQjEklGVcwQ+30QOMgZe3LkwHjKgS2ysiwYYpTisxwThxXVifAb
qjxlZVhKluQo4MZ/JfZAlzL5Gu6Dqfq6yZBlww9vIZR6U+JSQJk7MXsvxAya6lDxrEVWXVY2N7lj
fe4o30CEfHJ4Q6xXUO/2oOWV37TpF3NPqCRkIBnsMAOu5/RQSzeC3riDMqip5zRk55C49IhON3Dy
ukf/q8+GiPFFqZLJ7wL95G+Ku9xEbYZz6+HFZmS5Ex9GZqdL+2zUVAueaXUoSrswYYbpVxYfGQgF
RT4zwNx5CGt0CgCHz5f5lHrGmqqzBrCoBHd7wvFP9A3Jiz0eRsRw/c0/YTZddtGoFTflkgGMUPNB
CgV8mHaGQm0fQI5iXbh1PZXzKvlHeN3kGGrpluNsrocvxKn/tH/rkibQG8KiKYZVnIT76FFhvnpp
79hiYhAjc+yJvfOkz2nUF3pZK2VkntNA5y2f/U7NybdDOMJpMRTFbpm5XGnqCaaRnOTGn5DlSm7a
OLSa9qONsWtQ+M4jDsjkg5paa4++8fX6uB+pG1nWv7rkN2M47JbrhI6V8pWzetaJ2RqpFO4rxzVq
WNbFraq05ga2YZY4Xuj5sm4/W/FTwSrWRiVKYv1N7szEBqipOXA/ycn+bCta7fxJwa4gbzfq4woU
Id6WAo3qp0GrXT2+5C96sNNlmAOS6qxKyE2LGY+fzO76zVGTtDbJ0WgT1c/XbP167FRxif7gLy5B
Agz/iZVbQSkFvmgNcOO/0w1p8xw7gDdwpA163CwWuVBML8jG4dbylQyd1it6IImckwlDPuHqQle8
PtS1AY+UA06Aa+HOCwxqrmdTCqL+pOUcYwkA/0AjWvuAQfk8JhWFB/7PACHWrvhNh5PepOYwvJdl
1rp0e4qy7dReE17HQ+uaCprQN82AIu0xL2ufm9KhQfXgvePfFXm5gK7Vhh/jdwJ9sWXwnCGZ2Nhq
kr7yR6JBGr4Us2XwOBBuYpMEmpgEsCPLTK/RnwJo9AbqooUZSCCRt4C23YbxLoJoC8L3i0g3V/P6
D+ptfACLXq2186RZ0YrfRlOGOZF1aLfVqSST1bjop1+V6Ed+sQXrnjPSUOos1PpnSajKs/L7VvGp
o9iCvvE3ry97zvTR+QAXMdd4P1CNiMhw3P9xHIYrZYneWzv4lubAqoE8fJCkKRqverijlDsYZrsx
8JfDx4qAKbW+tQazkXIrxQeYIfJprtbPTie6okVxQJgu6trB7eDus2aSueAmCqmJAfNuWSshLQsX
3ZRa6+nE5QpWqbnlajtpaEcglk4lmSIhVrwBmvWZJnvVY9ePKbhHHlUXRJHdVEJ1Ag631giqIG+5
i+HuX7aOZJCrcH0du3NcZceD7hZ+vTO0W8stVe38j9167RJlXeFqRTN9U8fMhiAo29S2Qha33GsV
IcbmLND6AE6lDKd9c44mEM84WXL93u4phDqnXQJrGXpbUSG8YY9weGz5l7tt8k0tYQO90l8LucWq
0pJrOqDMmornl5OmCv4BQ0yNjV753Ze1zp9EcqX2TZtjlXzi/xB/jyhZg1Gs4yqpHMty1J++/sQd
NfkFHxtxt/THF70A7fKO2fnygOkJFI/7HRfJDWrcLoTrvBI+QM1uiQPJgAQ3ock7axOMJ5i+uNlp
qFv5Sa4/taRSYhE6HJdTo/FkW/UFg0xqCtBOeID+PCZqNA6VzAm2OsQ22H1MusmmKmiL9erv2Hpg
un4F39tmje0ZyaA6NW+dLzhGAwWbqMYy8zCgSe68dwdF5k+QM4opfkLiinINwWhY3TQHCBr78qsG
VoTugRArSc2GlPTPG20xLCdmYnSB8GpM8y2fza/e3w2+nTnBEE/PFQ7alzMzhYVQ4qVLV8nMBqzM
YAWQuArniX7bef751Lqra2OP5OMrZOz5BJlm0hrxAVSTQBo9EkEVR656wsmuU8JSL9TaR+4TgswQ
MBW266Zr7cKpsg3Ts8QoU1VKEdM/WKsDPh1WcZPZlZkdcjcDrj6lLGfL2tuJXDoBNakVBgNRVFDI
YEse3j1RsdluHN5p0QjDad0JcUoVRLPhorV8Ef+FSkhWzLDfOMgu27VgPLibMGMFvP2K8LLoHuye
1xPNOZOvuD7Atn1YArLV/DJCk0bp85TdziKkNhiAISo6dk2w9PZ8hsWtRd1TwzTemx9KJQqOijx/
pXrkjwLTI5o3qL2XMPqhz+9q62veDDtKmKoJpbxhH16+0oM2DS3ZPIxO9lMYL9ouP6iDsTrJF9xx
kC//WkDgmGGzU5C86PmvArp0rH89pVjwcuNxhmVcELBcg6oRGdN7fTU+sE8c/++4wpALKjEyZnGp
+wR4YgCyDAuRkxufY2VffTnQdr7shoD4pCTIBvurCl05dkmfC50EAGAO/oOKVNqQeC01Q1LqOtFM
kLYN67PUYKd46Dzpw9Egqj+W0PUCC2T98Zur7D6q8dBRh4qKCy/ilcnma3JOOcmvlkaOW00PpJlQ
EIwOmXsdPUI6seR1oko/o9QNoAmjrwTwLltCPdhWULTTUqL7gXs0u9j9V2bT+aah/uCpwXks5xeN
kUVVf6uNVLPSK9+c/zCLlYPKjmscvutCCmV0/YswepnZFpwr7gS1JJv2hYqS10n1ioi1t7F3UmdQ
pHU/BxuGMV1kDD7VbVnK4HxlQutmfVXqLbzHA11V7uBoIj6xmlQDFXewxYOr2EmzOmsGyjfKXIFn
N0270pzuH11wbDdVQS6DooCyE/nIz4NyQq2TUSUHvPbOKo9K1fhPeWTHuEKJUizymEyM9Vz7F76b
RqxC13SKV12Q3ll4uPiv2vX3pVn3+BSlYcVDVvKo0gNeeHE3B5PwXMCkVl5VzIXur8T5CmDgkMtu
NbmR9J5WU6oxP+4W1MndW263BN/aHpBDhhhKqMsU29YsyC0RsoQcdlthpIqD2EsJ+tMHAAAtPYM8
+1OYV8sbeVIT/zWgSvF3jPkxNrLxCRd9j3jfp8KTGLMa318I0mOvLj5/NsMKV2K1hu2XhgdTFCq8
flaA/tcnH9jFbGRHjhfQfxu17hdJEj8vuOAQfwP6jzPqTG1uJEMGatCQbpvS6h9Nyud5n9zc/ARH
3+4Z/8+axM9MFjQwdy1681iXYQD4y58Ko+Nq/Nww6FUMiAafeeZShiGKjJcmi9vGXJsDVfA0t/qX
xLG2O3wgCWTAVdtMb0NgWwG3w1eVAx+j6mNu5bxRMZU9D0cRVHSs2SfYom9/Il3kIZF1xxY3ZYtW
i4NVue7cu7i693VD65NaQnLOgupgenxaOzkLlwEf9u0bKo+HGty1nOZLlatnnLLtX25IvRPHZRZi
URvup2KCxGBZxCmQwV75RTegYu9dDZ0ft4k0hHaqQ10sq45nW91YZz8TbTb/JI8lqHtJxxDI+DeT
9tN65c2/uhlcoqiiLTUqhJsRwrxYkJDmndy/AdvAo19LPK67Y3yCgclzsAaJrxiZlD6PNcf3KDZm
15pCPp24bgJjuwSsWtioDxdBoEnNpmqQ4n5SD/N1CtGfvT7dntgPov6zqfosIgTsOjhucjkunhly
te1BorAGL405fXe8hTDBb5WjNZOcKDHsam+CvF/sKW+Fi6UsHsRuLx/6gOnDA+SQ/OnRkxTRavpc
5YeanRMCZjWXU6ftWP7JkXxbexraYXZIxU/OdmFeHwfrSwtmSGaahl2CyViQiOrP2kArzuxwbuz2
V9bYfL/0Oyg6oGvUlPqOmpgc9tBvgbOYBNqxt3CUUOMeMzPk5kwTKe3xhGekFst0dui2wZrZkmP1
PXBimLSeWg6ROPxyczYwtLAV/k7ohyXS/nhvDyaO61gocweAdeuC0BvmUU1dvyeMN35w6R7QMaw8
EOicgWLqSWJDkzM9bn7SEBUJ1Za54twXX5yXtxi7HN61R8pMkrVcXCjwcLI6VLkTEzLdLgfTQU1l
iyzu1T5X+VKQOrvebJ7YXickB4xxFTjEKwz5T66D3PLftBdYe/CwdqZrfw/2UxFi1qkZGPCoWUYa
ursSuFsLf3fCSigqiumHMKpTMZJhniOvU6HUxMcQ5sHmlozZ4PnTZEhRPx3aIjuVh21UCfBpbHh4
UIc/u2qGPzegO+3lpVmYnhCbHNyu0wJ5TUBGX8JkiegmM9uX8i6MelQdzspJkeEjuTaDnodDZdQX
Ru1Cn1N7WjKrHRNyjWbJQIQd7BYbGUx+dBKHdCSQL3dwvGzp3UOaqynLh83JLVv8nGDn1d913sca
r+2focdNuQ9cBhvuNz1fSfa7tncOeCik+BZRqtAXnnifx9WEHvNm3wLIqa1+j5fdKbPFzcZBc6Sa
obVgD2uCXABKQAfkIU3pwdySPx/qqJIkUnW4VKjtWECryPA4707oY4U/o3AkhmrCH79HaJYSdsER
xALIsHBm31aJKWsM1JZlmKtnp6tOFz3JqPsHiCLslPNVEokKDkeHyfyrxyKiWHf3ZwQTeoP6+tmx
dKLceU5QY3u7hHD9uK99usC6iJ8eHAHTt/48WWKcd2LtKRgFe7t7danRIKc2VgtvBZGG6FR8M0B9
uISCIj+RyYZhBaJiAPov9lsbOWX35bAAcMClOvhl8sR+aQslNx9GjDkmcDfvMeMfiy6lIYb/+aDA
6ORzR/GwsCTkFxLEBXQsti9ji7fyRoUAfppGG7rL3jGavkcjZFs1QGdUYwkUoC5w7SxFhv1JTu2F
u3GIDOyNUNt827HMbams1U45/3zQRId235szf8J18x6zctLcGre5FE79vvanHZRmJ52rO8RYxmuJ
5UlvO9JlnuVOUUj5VFviOjG2vWb1l1/gxc/tEQ7K5XD3Qo05P2U4wMFnDzHcpdnbk1jp2oD1oLzJ
QuKeD54PssIIxmkEiA/qkZJ/terT80yL8JrwPENd5qPz5fBkokKSJ3EBS7MwR45axOxc3zyP0QuY
dk/Yzhvnpmz0tm7KrI7axnsQtSeLepAYK6HRf2SI+zLgWKRwYKxqHeCzGw0em+wEFkdaR28UvVSr
quETwUPY0PWdReSbwusTMJ2jlbx06fqB5CtUokNrrQLDZuII15RyEmLIikAOuTPpcNjTokQMPL6t
vGEoKi2i6fjHEG2t2HllnMoIGgLifsYMsoO6SQufIExHB0LWr9CAx9pt+g9o8q0E/Gf66Z/wzXwz
V6nlAiYLnjsBo2Dyq6tMzK6Ywh+55BrzQd5ta478MxYjK+Baa146eIjLlAgua23MPwp/thyQLDtz
JWYpcflgYTkK1LV0jd37yArCl3EQwcdJmQcz4+DB1kvf+0A5ucIBYMwQIf00Loktvp+Lf/PTf1X7
CtmF53n6iRgOM2RIVMK6O4EyPwITemjr6dpJgqYqkiCJ4+adEMoqcST9cHqQAgXKENasg5GYUqGQ
RRNl9wUUDlEsDFN5jDbqLtDwNWM8SS290tLYY1ZtKnu4cLs6Vn5Cv2EZShUTe6QsDdEveQF9iJa6
+5Gsfa7Q4f2Dft4PG1Wq7hcSccdEBizrCeVtyn3WJ+OcdeQRjOU3AUQKwiOwkIuJvZE4GjNz1qQl
0NKpYD7DXoa8Yz193ML2tSbtOFsUmmbtPuDertkFPkceMIk/9cRjWeCaFER7nivjV0synG0PTNHX
ud9HZdwdCBe7eWWYGKK1R+BX3YUSHblL1cF7FuBJux+QmmyaJJ+T3l/FTT28RREiNOXm+8IRcsOT
26f/Cyh5ZTgtqxfE7GQ4JFMefXupEk3SeDIp+yiSb0gYfZRnHdYIIeYx3ryN4cxAfNs2Tzj4wAy9
SpKnkrIBc+5PE6VTf+a/17cHZwSibvWFTDmCBGU9WxR2ySPahCMKaCRHe/bgtwBE2F3mwcrVnffG
Vxy2S6DlBttM1v2YM+BNXt/8E7tfpGkBc5ciwAIuAj/bM3yULaygT/kWUeFkkCYbAISiLMCqhjyb
fY6OK8ilhy6hsguM3kB6FHG4BoDw5IDkRpqco4D9v2FsqBLfjuLZsnPUfaCXTmmthKUPnHvUwgZA
EFAZGk+EplzXcHP+yojBznNe2JodgiLP373+05ggFyVQkYlxdWrb5ITEcic3waP99Vp83fl96n9v
mhOBWTz3tLslylbrgAiPvHltuRzeQ7JNQDADKnQhy8Ock2rXABZEff6HMhyto/wNGcCjil+j5g9N
A9ecgMLnToYNCjrniiWr5ALESLkJ2row9ZVE3FXLwJ5SUyTuwmy+Q+PkLfrOENwid0h8NgpaC7Xb
etALZHH5ud4ttYU2hCoAsCcF+b9VnM0LmY9gq12+KVk+bBx9Hl5IJtfT/ONTEl/ogd67/gNgN5J7
htaXiyHNsN8pC2TYw05xEBy130X3vf3cSXC03QZEv7EwjD9FMKqxkUlp/3T639eG0L+6Tbtn9Sk+
dQ4HkVIrxZ4LNYixF6R3kj6t9zvtUKCarTF1XnEEgpTWXvv5msK+KQNoX20ttnEl5MdvAkCBmHvs
UqUSZYZRgNhEjXEmLFi6ayHKa2m1wVmn8zDvPBXPR5NpFsm5Gjs9DYpTyKdDkMVIfrX5lGKN+GIz
0Bdb+vxNeUMz2lG32Ds8+sTwrrcZdoLVHlMBuR/i9s2q+ngVyJyt4dCWI2eAA2vLM+skqh9P04Sp
kcpn3IkseqgO9Xa/NtdIDy1UlyPnCaNTTrRV2QcKTnMdNQsPSuEWDTHNNeZzrKEZbXhjYAwGjmCq
KNpHPqjmEZQQghA91XiXGoWBnGj+kd1SBxzTVgkgCUKtWQR3j1KQgOU5XgL99F8+T6AaBOOdMb8I
4/7OoYnuB164RfE9M5gpXkwfAhIJAvYzwxpxUgNjRTAGva5z3m28/bEsFlg28g3fS3uqkwruIEj9
Qh8VSMLTnj6+Pw9guZ7/bk9vlpdDHaa0Zfz/HlnluP/K75g8vsHhVcsQl37GaY25tLElz4FcGwNc
vQmfr2vUKBbnYOfEnvSHAu0BzUbz1UYWq6BcIVV/KMNFacuSRL9rPIFjTSuuH0q6sBvDL1SULeJr
JJ1nCxgQ/sHsTUb6PTK1QyuMdP8dPrLxfD28o51zFcwn2RMItaDjm4MvvKGaRG8D8EHNkFRFjQRt
+a8ku9i1lLL3uVhD3FYpFnqgx4qnhFYuhQUX17FsGqHgtAMBcxhfe7j9FOsrzy4KjCsTrVHk/Uia
9bX702ywncG9VSteSHsNo6CGpcS/laraBjs+criiBvLr/hJOFE3QGGPIaJFY/wFx9HpHQE7mnYU3
mnooZIiDl9RcRLVQXX/AeoQD5upuldy56XmUOnhOK798uOmewfkwBn6k2SOFZmt5rprFKWY/6ge+
zb4rxCdk20+UkJkesRoyh6VWQl/g3SAe6Po2z+1ks/dWD6uTBrFv+KA81Yg6HCfxiI+HCB7xioGj
rNlDw895C+C9qL0XWC7I1mn3YllNfCUR1X14a6q0Ow4Out02bJXAJQHLX53egJRkk/8pYXMIVBZg
wC6O76oueRspveIH0dT4R5p8++CyD5lhLyR/UA+b6WRuMBGeHaG06ZXilVtjjigjp8THB6F1qHHy
kgpsdQdmX/TKrEEwROjSJjIfEvMA7YroTfYXH5Bjo43bEXIkJotWXhdaZeZq2yzo6/jckQ0IH4Yq
3SwA9ETDlfLmo3RWZIsd7iZuH7RzQz9XZ0B7juaUDRZtzzsQxuwpqjihv5DsVwBhtY1evH13XGkT
uBF+ReCbe3bdglT+83Yk2vl2a6dJsqOFDvdco9uvWntzr6lGx6n+5QsR472cqYXRNd9AqVWZ5rLl
GcL/ruvG7EE80DauPdX95mwAWdqTpVIOU83fgKhLWAqiibGCWq5UMb+eZ5AyOvcuoQFNRwaXVeye
9xVU2/WtO9Oh+E1j9qd5HFMWgyne2MqBdFVwGHxQfsZhVeRG1KS5VL9S6ZnYAQhgkvIYKXyvE+Aa
CjCejNQOqQAFEvRB4D4MYCp+019HMnBQizDAQSGpGClSv+QJMspnrfusbHLK8qlCudw0hiwkLMWd
idYCp9rvd9aTVU4iQSiS+OONSX/JGPKz22qS8gocRKD1CKubwNGrHVP77psTFoN2zsTshKe5ZgX/
PnDGhmvvubdfi3H09o4wggLSuG7QLhys+H/YvroQ3oApYoIRlfXdjiLEKNliVGeLorTJUr+KcGsM
3MWAa/tGCz+2GsdJdzT1mQG0Scw55BtnfSWMpkE4OkpxZifCfnFvzfeqrBYEqjikQbgDRq4w8WXG
pulL5VE+1P7roChnfqV4EX6G5uqfuZU5DM1pqC3ndh8IMSRWnxyyEU0EDDeE18PA2gEtcHybClsV
SiNiRYK5l+sf0/s2KKBzBohlLugAXiuYJ3oZKgtRnPXvfbbDXJ7bpY6pRVR9sE+0BHCoDFgQW3RF
wnLx68ap8ezhP8zE1AquBqfilp3R5hgt2OddoQahQJw60OyZjF3YP1Fmz7XZzoTf11ORxSq0nROM
X659k+MG1Xk5jUqAlUKjRHnPHL2496UBMlKTyaMrh3/g7CqbSQ5IdT9ZlwpQOQxfatcjDQxKbstR
ZuHg48xZF4kjevl1Q1zGBXun+aThB6VNJ4+e8h6e2dDMYZx4LJAIZujp1TsHVZeLcQKHtjjPXYkM
jjxJv49Gwe7wxcFeDh5XTHLuf2Tw6Bo9BI3TX/kAhOeuHwDV+xbqSq7qORE6p3vgI6NmC8qg7XlY
FcBWFfAImePBqE0ts8m2cZMbONWMBSkJnApJV9PshpBs4aO9Jf01Td7ZnyJUX5nGOvB1h2dd8dB0
M3pd4MeRAEBsgdwPKG+X0EkBzMZH4h0e+u+FjtOigUBETuIGugzW/AeuPoCEMzf7sFdF1KCVTd40
uo96wQaSQ1IwHbg5lbLLCz7ydt8NNAGKp7JpIlmNeQw1XNjLngAvJd2pK5Gqn6LFmxGoaqZS+38W
ccXiRL4SEwoVcH1APPDvV1S42x2OWKJ/FYWnK6qYu+WL7ki/mzxtWMYlrBV8+730l2wcwuh0o32C
0OCJamW/d3ob4MfuaeoMrk24sH4mA9NFOMNQG9xNlm3yt1YhFAE9K3BQ0mVKVJ9ME7FgLSwp4Bih
1x9PigWzcfpLiMpLZeJBkzR5Xw8F4Bl7f3PLCzpEzMl98a4T0Z+17QPrIVUtBZ8jnBzUc0gaaLuj
1TrDhrmn+VQu4Va07yLYdJcKcStkewK5wb8H2BUTsMo8o+kfO5I7qVm7RtmzeUjI5WXc1eCcfaDL
6fW07mOIL/NH2eiZOxkUUay0SBOlJfnLvDLtqot4slkJu9del+jovVwt0udk04XkkS1stE2/SnBw
in0G7wZs6QTGvS3wxLYB2NPSCE5f3Y3SZDMutBENzrUQCAh4XLq9yByDlJz1XkhsoDBZW9WgAg34
Q0CYhb4wQS5zco/K6vXSwYgrZJdBxK4dQFYCA1l+6VzvfX3U70IoxsQ071WbqxsSqqhZKlk/1PXW
QgDRh0spZM2YgwJCwxAlXJsi38Eh63nfC6OgVBAM9//liQy01PK4v3PQtAayTWoGmDkyO/jOtwMQ
ehBpaQGwMtZ0LDkJ5SWKcziO+R6c9dUofi4hDu70MMNoda8kPWQz3JQPqxn+2amA70nIFdfqwjzU
rBM2H9qvQ/Wud0U8IXpAZYQHAKoJNJjTZQMwaU24VjRvw9y2G9RMGm6B2oAPPfiJEWAeqQMJtJnk
j55L8F1fhZueWUC3Rw9WLvPi+mB42CfDuVy3qGkJ7RDNNCKaF+Q8KwBZ78ceyxuptCC6zm4pmJwR
r/73eyFMs7GAgelJNbz9fkpg7L/f7RJVMtSdlftJsVh16c24nBEzifrQbm5+/5ks6M/EfufmjBxt
dqfbdIc6c5Uak/7Xw1j9Q30wHy0cJe9uO18PszpkeTR35p+N6iRlZXlQJGEEWxNEaR0L8eMZmndU
bpDixrMtXEVeKrEgFDuFxnYeNPwKpvbjvMPmufALQK9Q6o+ikAhdMReojuX8BoR7AfcQm+XsQpn7
5EmbQyfvKspE30XGXSgQ6iezhBGw0/9xinbbqeSHuMPVDaZ4Lja7ayUqTFMGsXT++ULM0ET9vou1
XiPSnk6Mw7LSkh39TWB+VUcOwxMXBZU5aMwONm4cnQcq7Qjb5U6dJSQaVuyO///4srTbTCW3G/1A
DBZkt656C7qDZ25xre97rztjxf5EsgPIZjVFE4r4bLw9cjmy3LGC2u5YfQkmTRdORPQJ1wB5w4Vc
EXh4NZKLoEfi+mzbK1FgcIsNfoj6tPY2dXUQtApoaMXfneej09oQ29cYiACICm3/gqFRht6jeLZy
9Dt963wlN8kAJLvkelFKR/MXM9MxCElS1giJGo/ImNAL4yWq8k7cuqnuTGrqKipSHafSmcOthl+E
zfGPc3jkdKidB7wkIjEEFiBbgNWN0TcSOCtQihysyCxGnlqfkJTUjptu62rar0Sw4PlqA5ZRpNwN
f4kSTmQtmF0Ur9VYNlyKICoeQRlEbkDJNndZ7fobCH3ogAXidQJMnNgiPd7kCgmzBGYJ5I5j4Kyi
uGSDdPpPs4Z+DzpMjGDpS4V52WBSYLzN6+bMKC3IlX3Zkdh85UPCjEzMKa1yBaAMo2jFDhhZ77Rj
wYZ28IHwGK5OrwHM9QoxGdpQ4hjwNduQw0AydDzrgNxtIhHR/fsMVg+glwX+9egDU2boohXG8g/4
bxaz6Wijxt01RtsMKS1j/QCo60O349vnwqN2Yp5wI6ZnrLEzB1Dwj0i0I6VCbjuNDhMa1yYoPvE6
YMaXE9cggB5P7zOfzb6inoIeRuJ43N1mIQnheRQ2wBk4XNzJRSTTmM+bQvoGkJQxPhgVBr1xLW8A
dfzy/EutSoKPrlaGPZqFP9qVHsUE4vFoPSc0l5ubJ1l0Rq8WWNIY2h3aQq8u4Xd+VvKe/l5rDzit
+PU4UttL4rtq0CYKYNrLgi9PjeP6MSC6VmkrYvER5sy0rMTc9hgXaDJjQKgsNqgFFK6XSchRHaOQ
5/K+ic+BJprxcUnAzBidMzGMMsHUdHNtYrexyMz02rpcoThAMOxv/AZCDAnlqOaBCXR1PP8YWSbP
03iGHu1qwZrqVOJCZ/TXHWSD/65S++nIkhPnHDKLxEt+KYC40jhc43eStOWuNjvfkv+GNRJ/9/BA
RegKLISdIjfQS+8X8w/t6JrV+0EL4gp3zMUOhXuGT2/qE2QxJOaepVvsBM+rFKQIk17DeamafQLM
UTfoA43UuorKg8cZiyarMJfmKDAB5+1Ow0Ik88yvBeXr7ukgIZ+h6pry+sjRa8p+UenmCWHIIVKh
3jN7fLauB/ZUeimxR32PIgzP3i+R/cYD5jeYuTHA8INL/LifNl5nT+FuTR6VTyI+fT7vUuJw8Q5L
V1Fq9EJxrjHOKOTur5meR6TRMMd1DopoVH3bWrWH11K3vx+0fUWd2bGjJS341Ev2zBLcKGB173LY
pCdUeXXPXSG5HTP3Z/ZQicDkEKh7ED/M07PuyJtFLQO56Zyu55PIuLh/dVr3MbK/DYjcR2D6vcvx
JLqFzuKURy5lJ3MCBQYEFG+WDSdxXf0MtWWzRi309ec2bOmPe6AiqI2N07sqL0vaTeL3iq86XIde
InIXPY6s/TA5Q4NICvGYqHqqXyhj7RKanjl1nVWvVIgE167Xz1TSOArndyV2q0ipzKbHZqfnmNtn
oqloc6XYfsklTqVv532zFKpQcaUz3ZnoV3jX+9UQFkRgfWdB1IWWwaYCqWbYYjjQGFIzmZQuZFfU
3o+J6NLiVMBUuW/WKo+UMOCFCUg9DBiUQzRfI+mZsM+pjcV5IlBGcs03QDNRHHCjNdFakertW6vF
ktMg4Xr45PzCKWGUeUfQcTxDZcSwYjvLZB6Q+PTnYJ8hEuBJ3a1+VUchu/fJusOwTcqoexh9FA2v
LadBJMVLprn4PRXdvF7c6xhOjJo8nnMQ5PprM5wkLKkkl6uGt9Y1hpaQUn+BGYXHuOFaXcmPKvKL
JzU8jYljA51PBsz6Iih8cmhSF7OnQrP2pioKDM0R4Os8nmMDYN845qs5veNVMWPSD1VpbtOwkoPN
pzxdOyhuOIHWFuIJ2dnNFrOgVa9J1icqn0rzue5BIXF7SGSdsYcytipOnb7gZXsdqwP0ebiNSH5r
Y1DUm0o8ydB3zf4xmlgkC+ImBFs0pkN2RFeIZoZZXOuJZEbBEINAHCzlSZ8JWicFSuSIy1LtUL/Y
STZ1GEO0yyzsD2FeozhnjQg6WtEO3o1JI5mCURbuug4Z2WnCpz0F2VcrwfgQE8gunsm2pNWBjWfr
t3ROzz3xxQ3AlM1sYalxzPMoBzzjyawST5gk2R/XRDSWvT5e+Cd3weRScXM+82s4rr9h3cWdJnpr
SrySCHYgtidA1Oe0DeqNEBumkUmvMCWo8pNNg4pDxbbOz3BCSDW8nRttvsa9wX1MhE93ealCiNMF
hUn6nGcSHXJOSFp0zc2VboqZF8qM4qLnYLrZ+Mf+vtkgGRK+9sw4Ufh9BX79VwYtCd7lYxVYftTu
IFN01aKaxSZqQCxa4MNDqeUOf538fKSHIcj8khuMUfBzP1e3jX15UpHiZ/2Mi0gOyKctJ7TRj8R5
Ppthvcgp2vJcDwkui5wQGoGWu1tlslTX3lhEM6GIO/MQJeXYbcEpiaJ9mk1H+QAIJr2sTufU2geU
t9aJ1Wp1oW8DyQuKC468pf/oHc9EzZQ+kOZLXjlh0ywPjW6jTkfb1jzWuyPvc7hboH36HMNGelfn
DEzznNuIRrsnoWafTREvPuTV13HQLBtIl2uHHxy7KEZOmDQHmQKb5uumMbtK3cnKcogNfrsd2++a
kKlmCsloAXJajaBBjGmN+3CXaSVQY3vLlEjiZoaq3GetpOpLLK8lf3HWLMnXxyFcBqiOW3gpaW2+
GH18d+BLpGqazsoS0mWqDiW6E7jX+IlX/SpEOppTmNalINdBQOS9aZyvlegfSvgYXjNodJWW7yQQ
xVygJ6qh/Lo1PogP5MPlQbJkcex3bOXIQu9mFrrcsJXid9MCWZqxaVuJWlhtg3LDOSK97em2byxG
tJXboeGhRrn5hsfCni7K8jry4CACyPEBUGZsjxc4qGwqgrKFATTp2Qf7aZzzZrnbiHHEUXH77SRL
+HEEgDkJhv742mD+w8UcFGlujh9Tiw0l1pyVhe61mfOqXssTOvb8Hkc2ytyrrH2P7QnLIsDb7F1E
MTudCx5f0j/ni7Twq6G+RUDvz9YPm60PiEMoknwZ94oqa9OF2k39wTWepm0PIpTTkbcrtjzqslkq
YYkuLHGHIAgJNIphjkCUdyn+h7Sf6VUM0hFmUBMsuDTDVTH/eB1ANExFR2iUZyKQYq0wH4AThkkY
PClDHS4SW/yAF9kvZnPjqpY5J80+XuzzWaWmADoCizEIj0KUNtp/HVjlpiU9DDRBlK6uuE9fC0Hy
ywORjnkiF/ws6N54okQsrqNTZC4um28woUM888ZowhVcZHBXHVcbkrMxkvd3maK3GGsHD/JzOkeq
g13dSZvsiKeZ6P/0lvShll1LCyq/6k1bHZVdWuDYR6kmu0ShuycKDt7pr1rmZEzdFJyvd7whmNOy
MRmUKRh8mstI+BuQkhWm5Z2a4T4QRz9BoxeNsJe13RflQsKNVRlQEE066JvKQSLSa+eUtX3G/fL6
bMlmsUMDI5NCMPTWqY8zZn97j/glGpq3mEJrkhauDodY5Mzjhsfwr/pQsLS55+sfStipT0LDGCV9
TIfz/vRxtl2ZhTAb0Wl4ng1sOrc+kXKUIP5LYWm3xeav2x8dY9gqSwA1lUJatyQxvtfc7r2EkOl5
PFocd7mZgSFE/g733I1IAsUSds3gY60J/WCr/xAJv0ZSv5TZ4hwjsHmqQQfLEYGyX8pJ4NO3LbnO
nUNp35ZDAYOElyF3XOaFVcatx//KXwzH1ZbC1seArCFJBmj4NKrnzRvoFPhHJsIywDOMasmJ0Gs3
6S3HPWGjqrSWdT7xGPPU2bmceHagD5Zo1pyrTPkJxofQmyUo1OHMO9VthhBOJIMg0wlDKLTby1Se
BHPTUBkpYaz9vf0JliAH0GLk0eVCihzQT0Zn44xsRteMI5CCUV3ftcOlHDsjg7M/n528oDmXwZej
nrBqKDeRxP+YIOPmRG5NZgUTrGhSkcHTSsh8aRth1tafWs8KJu+WxariVFjpqDzE7cmYbNBHYBp+
Pi467s+ZHarAVzoogy3zDdp19wY60Y72dQNSNGpq154EzgkRfu4bTXYtt/xGQUikOZuMZXsLTvSd
zvlZLfPIAMT1XjExcKqpeIreZYZ7yMLM86M5z6Pn1kZpVSuiVjO7EXxLO9+k+QpbVxYYGIgwWV+9
jgagkMGsZPrQFb5PqKPhdt13OBMgnPjoEpTTG8DLMir1KALwi2A4l5et28EO/ZrA9TetIN9774xq
Nr1QugRo2vUe+3nugjlx+FlJtTT09xig+jiPzVU1nE1sv1EF2N0Xb5GZ0M2z5+1RLx+Bzn677Hqi
e8nTTh2MzMkAE3PNiIz11/5YOvRLEXFqzMm5aVdvmAl8Gm1ETPo6DE95IDLxQ9zH7upKoK2vnOUp
YESs4ht0lFJ6Mv/M2mEhtPpeFm4v1fQglifINH6biCF/wQGrHdw5gbeM8M6Jc0CGJZwU9Atwlz3c
xNKl5p00/7Ma2WO7622I7Ad2KIJ/dOr9RK8jnkECy4Xy/fzHkB0CgFQU8MTFTWZDsm0GnittCMQP
QoqIrOWeG4SkJEKe5m9CvDVkTfUxZjf7sM3YsDQf0A23bSiZL4JOpdk9Uk7sH5jybOcK9wXKKEsE
vz4ycDVuxNddyotDbeBvn+uhQq6MYx3cjAn2VyBRgwRKkkWwYI6Yr8NrbLhc8CVz5yLZdUeAK/yi
eyEXC6xdfyDwfye9N4xKM2OAndZyp1RY5gndbfjF9CUmcoDTZoc9ayqz8HOFLfbjWVPBoohPjY4b
giYe4j4JGPjakd+TtNonpaXG7RarsG/fUACaQlO2hOw3Nd1Gxx6Jd8eOwLEVcAXCkqsmc3BLF7Ql
bWDVGmZH20AKKOW7XszKMLRr4eWJITvgBvoNSi3zBeWFdNMoI317Axzm5GZOzScY1+eUoenJ3gw/
HCAai9ICO0F5a7uyKksd1QQiQyXMCR8yjsB61xU4IEXOzDo54SX4UaxMvK/Iy/B4zPaMRiXTt6MG
YdS93LxTdpCZFuFBMfWu4ez2zKZz+/NegbWKqL5sH5fjScrj3VwloGDsL2Tbyj4WyOp8sKEnN0IJ
TyZ91zdIG5KlvnXb0b9htEfBsuJck33ovM4xoeNcovsiWRmNMOS6z6NBdMFrG8eTU0hCie6w0y+F
JNeuj6HXHcdTiGbSVYWGoWweQGelwk7iBGuqJH5671dAmG5dEpcgACg1qUOGAbLGsNFkbwUlQBJX
bu6MzmIRUw2RjV7ufHSUyiz3V0RGWN466fYfsTeXE+QNkouYmAv6xF148KK+Dquj/DOVRZI9AFCk
fuO3oZObT1x2myo5tv5Dwav2b0jaGD8h2WSN3AdOUVsYMTzDqdOe6NsCmlbWJQ6EDCA6f4eqQ0Lr
+p+WbTjsHfgwnBw6k5ctd0mt6sdbe+P5CS3Od2YFZMaOtLQkU8j8s2wB5dMr9D/D1SyggASZJuAt
a96if4PbMuQhupgOhwjeTSE4No/DbVjuIlwgqrBT+FpEBp+lOVsfMcQyMRD7E6SvnH8Y2zuC4dWn
qU0khp903izLYBQJhd2AAS+6QLJehXW0LtYb/LVRgc/DLDe1Cj06GAWEq1ikKcweITCGu9DpAXVV
nhG2UPagDyxcTQiTa2YxtmWWoxowg3guPwL/Y5zOzh7aYlhARFjSGAuuVylYFw+/BQ4nm4LRbxpx
UkHza518GoTXN+X7Gj8fo8AM318pD/rHR/7JuhMzPN4vyRZt2AMfGI1dl6UV89hhTfKeIsOLx8AT
vdg+vyp2ma9DU31q4/7Higu+K48yUW9X+MMBMMq9qkG6qHVp8PE9vsSDU3I/7jrQE5eVYAc+Byh5
YDykn4TxI+DUgaYkZjCdXbwmPRF+cptkWCNoE9QoDZhoHECEPGE/pIIzgCLe/rcCLUdeNoXcj0T2
ePmvDn6GsCReEHyEr08DDxVOW/KPaVH4Av5cZ1TQo2lmIUN0DmLCiWuzHmDDKGm6oLwEBG+OFpQL
xFjUxD1T0C0pXexmDQ/UYIHamg9/iAZfFFH5syZkFlt1m7nPC2x9844EGpsFZA9hVdsU+OynqxB1
cQrcmquxiwQ0pAA64CZUccYwH5uW8aiYURxCr48FaG1Cv8CI0c2PD0Ithy02IrPZFtHTeLr9Bkiq
OIU6CKlzOAkkpch1rmCB5QuhtKMRgJs5P1vp/v4sAZNZ365hVjl4buRLdejcCNRorXOpf5jLIjR9
g7jsyephH5vhxdMalhn85AKwxaxiuXIF02VUG7zZhyLcmFh4XXB/I5MNxj+SxIvn84zWYu6zlcsH
oXf/FIw0TYjuknj28qS1YPw58CcMGavYw9FK/9cz44uSj2yAfjX/CNYTy/e45lCbLikJIzT22rGU
XXorglxbWkRuVbwctoxgrclytkMg2NT5pDRzHqYh/kndxd2a6eFWVyvJwISlzp/vX4p+S3+HSP73
SYk+Gul5Qrn+QcFSP/HVYt6Jdo/ENmA9X7k346lUj6Uie6j1VKUjfWuLcgO87GU7CknBczOoHG+x
RxNpB4qDhWI6VFo7RMXR58pgNkoewHwG24faz+f0bEAg8hhx7s8wxhRJxP7/9F1MGBf7sVuijp/4
Ff+lw8wA0pRZpeSMDJrg9yIyVkZI+vW3Obcl1nD6rAPlNjh7darliCF+nzye/9sBKAfSh4JeL+zp
iwt6qukJve0s2Pgri271pg0nIFoWY4N3Mz78SbuoQZroWqa+yBj9GwZ20d5GYjHg2eICpMCwzS+m
KaU3/io7yWPGF9hSDoFaNNSkS+s9o80BBneqIAuhVhiH8KUPurGsPMyqjj+QYE0H3SVNFW9PDQcd
vCqsEDnFua8jwfTMfjFoQol8XD1Zg9bJRymoffxVkXj8V+eXcUg/Q8BlrH6UTe2nz8rYPlJ/h9KX
+TccX/TM5SlergsZ4XAuWzyZcnyJ36Nuru7vehXiev5RG6s5ivweJehxhKAdOZtZhmW2eksahsDn
/nj7MMbCvomyWsO3BNLeO5HtdUAVzr/VPDJm01gvdj6EEpfDF9+poU/Dbxqf98jsRyC0pLlkTY65
P7ZDWAFJsp+lNjDCaCSGtwsJMI39naehXolnNh5fyqm4zwRErU+BlIAI5cex4FtC/uEDS4lb6NzP
oa4ITZGCyANrAAAHNrfCJbiTEL1NNmKgkmuoXojP17XwlXyh3NFHTqSHv8ddIlGjzEKuRV8PbKEl
GP2DMItGs78YkQfFzV1OZy8ty/JISZ6Lxw8wjftb76kG/vmt4dIicG0qKuWaoWdvAA7r4ct/uXK7
EznFUByU/J17EgQ0iOWHwUGQEtA6jdD6sX3QBXzNj41cQLRL/npCG/veg0JRw3+/zb5NlhITrTjk
Es01ccsgdUO0aF5EGLfh09+a43L3Nex9oz3RQGCAM7TfipGz9n94s1JUNPgy1g/XVLg/8q3d6t2U
mpECGO8SCkI0Iz3J4FQHTI0FoSRbDMP5WW/AqYCi3Rqq9HPwMPNH7nIDggxKkc1HST1xjrQlRgL9
LYOH/i0Zx0frVLrW5GWAdazjh2CxMbDqTpfbc12OxWogB1cU7RCP+VHLoGMxDJDtvRQzQFIAivMU
5wg0DJs4VuMf1rCuqapLpN4JQYbXX9csUWGt0XOJBx/FyVjXmBACv3t96MAFhhbjtuGitOZAj62s
GknovWbYT9tq9TGCbaebdEprGPw1DjrxLNfRbQ8rUqY9FgSAlcgy8egwsxfwKkYAxcD3953Tkcyc
x+vSRLQOJOKIuX+JrNvRCXnqLTABn7vy9PgpJ3bEBDAifnJ5u7ZUJjSPVSjAZcyUVw/+PtvRNu0Q
TVZg7zcYqKArBjn0H6+gM+zbYjEmDanBvddTt1QsIuI0dCMfWCdHx0PQ+cwo1Q2Vt/LQjh67wL/9
RoTD8q3evfnnY6ed4QdhlLeXgObTDUxOZpzNxoMzkiIYuRCpIi2nKZwZaLkDyVRPxJs3kKQWcFX0
vIjA2Mj6VfgtFtIAh15fe5AgBkeojzlOOdB+cmlGPcOswglucgyPbSg0LzBXtyu+9oZq5x8fvaat
GmwFgNq/1kkfYkIUS1fzvkMDNeEnaVRygPDTHmhQz4F180OE4kJtC3r4aTIMfKlD+lnbQqev4PV1
vNk99f2mF0QxDpQaWnXEuOkiESUExHxFQEYYGnYMFfqIUWH3dJMc7q5SrZJYj4HCKDS/4KIrtmcA
fiFWy3NzxdN6HqBhqn+QZrFHieo74F7xYMy7kN81CD2NKT1zbDlo9E4e6KpuATyZi/QzIqQLbFEU
gw1vmPolPBt57HaZMmjHuj5v0wQeMFG2aiA8LdoHLlLyL2pPXkPAEOCEM6iC24Hi81dhObWYuBEG
HtuBe/6cSUvLNVqZiUYcZdQ9Gfu207MMfeorSkhsWZV2lU+ysslAU9c6LddhBxinPpYkmicGdUQ3
pUK0dZKqvSSQJG7gV4XzE/ssWt7JYg1exgL9toQFgqKRGotD2YT0HabxCoYniepRn1geeBTzkAXP
zf5g+9Ar+mIsOe42muF1W6xiTA84qjXeat2JQw0wjNE8yWaWnOnlR41hZfloGSGA9NeXCZMPk3xs
+gKoC54MkhgqyHxH63RcO1S4XpZOAW0Pq1DkrfCCsVtSXeiOQvmjUcbwDfKHT5EexBSq25fNd3Re
dBQ08ixJGqOU+WlDsVG9WreMyFiYgiRD1tMoS7j2qMYGGbLA8qMxGjzh5pJYMxEJMMA3J2EsSHGB
Oh/XsCJIb38+VPFXOMGLmuTanOLsszE5+Wxv3sSh8tAhURyhuiDQxMr4RB2E2clifowiHlGzKCab
TN4132FMSMXiFE6EPAvei043Tk2L8Ai6QIHiwU9bzcQWO14skkHDDHA5ZN+e04nw2LHvv0nUseCP
xgRehj9njLZcQIPbt/hUQxe9FWJTghtg7iLNNXketI2SypBQARqCTlv6h119SPy236dekWc/6RMG
SO2ab2/TyxDLLYTkHFYi2a0ue601b49MxjYRDhgXx4vTQjPHw2uqaE98+T+hOu/wDv1nVhHmHZmS
UKAkDQbXevj0qXPIKu6Apc4TmhbQN058y/RJu5LscaNB+/RZcPlVw18QaSSCQnoftSS+jsdIV4Ab
D/K8l/bQqCu3m06/GviOcJHHkN8I4GCaJ10ut0y7YnZf+GkqzMtpoo+Evz9Rbd7si45Y23e/tGpp
14Uj5tTIp7ZkXwauAqyzJMhDHPagmm99aIQH5O6YQFeyqlynxqUptx//6LPXkYCvlaiHXxxkCSi2
kmix9TcJs25ey0jUXVUGNrmzxd1Cu2bmRWrOQIW2yKjfhHiDXvidNfuMzZO1Ug0AQs8XVMfA2uUC
LbYvqnm5Dtp1pls6Z0jTNw/TxQRaIETl2c4Gw8Gfh3oxcSvH1XonDZbBKtQKXy0VQrfhGYFxTQH3
CnhDiqFcf69xAYyEjnc3aXtV0RWF5y0RDMB86irq52Bi0f2qPh8GkQeftanky86yl6LWuRlrhARf
C09aw99/zRqj6q/3CeVmhFqyE8IrykYm1mwKpVwhbmjynzJR+Xk4BwXXhqlxdQ44dbali5kdtA/S
fLmoifj8hDBMNZO96ak/ZLjo8umFjVDlMi1RWBxmYF9GjQrXLw0w4Nq/dEZgfZ9o6u5EfWqh3jfX
CCYvMJv8RTqn4DrvegAHUAEe7WPSqtR69pnDt23hOwtYg3+E0e8+tZLXuDO6GJNWdYDG7QtWfIGS
qx/+aDgH7TpwjNbW8jZMPYVfqs+5JRO6qjIizKboJuAVN/niovJb1XNpISUk/tkIf8XOu8iuB647
bSGDokqpjxgJsxeKacte/MVY+uRoP0O/zE8EDVtHv+hlydkNHC1bTCqh5gt7lfIg9gD2+dZt/kiE
qyRnTWl41LW1IYmIg4YF2wePATPPDPHgLtRIIZKNsW2vHX6CP000ku8t2u+GjmNszxdG+SN91fLD
yfaDSPioY+2eojobWU78fSGnFVTfB1wA1WLo8tUhsr7bDVODPRKD5iagrgC9CSfkZZONIqRayCMX
58hXKQRC3+uuBLCTW1vj7xm6/QR1JdKu4DuZynDWD1iblDzs1iUp8Ty4+8mPJCbmeuTg5faXOgP1
/qB9iALLeUAt3C2SozC3lOaeyBOtRCXQu8AlxB34nUgYtonG8ofPCZbFP4WbwLBYRBotlCNzbxKz
uZjOTWFvkBkWQbMBb5MvWb+29tq3yYdV8y5EYPGi2RMnz3+6aC4+aZeARB2oIltYnTxH8NmmY6/R
nLCTFHDpiS1nB5daYlQtq4UyUieXtMmR9cP4T14hkmriuGLl8T29JDWwTvX6YjvZP4uhF74+RuGH
k/0H7KGow/EoPecuHYML/2A1GNaQZQuXTKBoCytvriS+XJbFI20HldK9Y8kyzLdX/mYHpQ1NfBxy
sxm0nQwck66BFMh8Qc20PpM0dtQg1D+arQv9KaPBArE1T4BSiEgC0SQgOpOjG9KAsvImZGwHUbVe
XKMEGveLV71d+XmNPgIR4K2X7zHUm/xKPxUhGAuT+IJVxCbsQHqWpVL+2c0HDfhTmFJhlPdGd4t9
qBmS9+v4UOdyhXPIz3UGy8EddirdShAVuaRbys5KngWsYFPIXMwLY3+Zx5G1wPUXeuNkXm8+Kz9s
ANfZL+KscIQjqmbIG2i6375mJagfglsLu9LIyw7x2y0Ztek6lCzlwD+A59YEdaJRPTORmklSM2P9
6YFEIBLJ8Q+Y/rjgtyIR3/6o3nseMjtWD/cryyYfc9lQYcvTXYrJ9xr7//x4rYqUB4SxmSYkFVIp
H5hK7QqRKVJyPnfAgihs7THUrJbzOnf60SVJFSH1ECzGVjfqPTlOWreryozuVtTqjYizzJy2hdYy
lKHqu6nnDXix9rimtmaFsSaScKbf9LMJn88xtxiyfxLLCmXo9E8jFo09TlfUy9fWI9nkTYpIhgne
YThIzyTlgQ+5KpPOyViiGTRXU4BnziLBXJh6rVUq7kOCghnB5oqJrb7hSpyUD7POIY26SOolz2R0
qXYjyntmU0WYOXnb5jzts2/THBNyk4lT92pw6/+8p2/lkjVUyqTRbWw9lNTRtSSo7z64YNABurK9
cy/qxt+IiDD335RbgbtRid+WIMUI+PhDPcb1BWAsmWizv9gm/vQr9n1+/vpSgyx/9rYTHovGYe3q
nT+KsMFkdCW6qs4jjGtQZlXSIkpyWi+42/ni8RFXwWQFz3eLlXZJZof/eluxpI03ZUdFkA9Qa0j2
qHkJOc78LhaEZBDoOShhaIjy15pEt6HxqSgBCrYevK5YP6G99vtpQsf9yOnBL5PNb8D0ldfq+aTI
f6Nb/rZiMgkknf7rwYXdb/ziyRk3Q+oIPIg+hrGUbCnBmFsn+DY5avG9V5bXsoWRPctMvEfGXvVv
CKK6eFA/wW5GmXDnvXOCxtr3AUlNacmnF7omMnBd7CW9rNaUXUIc/orXe1dgVCD7p5mVri+9YiCr
+J0V1C7F1jqxsHkVxZeQwCDdR1Ba52F3PIFH2eQM3ZbUbWX94al4fWGqn+EYrb7OqEwkuYCB79v6
gk74ZdCKuhe35KMIulbfm6+mpdbj4tIZglVi10j0a6/flXUOEnC8wYnA+3kI5noKCesW753Zm0kF
NDLP57ro4TZ2ZU8RdXQFo6Ne3gtdU/WhEsNCm3p6N+OUZgHtMKRTiv09aiLdq7oKmBnCcpW3pJU8
yh4h/Om37TOr9jp8EJwNUNSYScxCDmbqmH6OBHamdjHoFfGhnBuo9hEvBniZ0zjNjhG+yobmG50u
S4Q70QeDz1pz0hv8gnz9KXs9vOsxsTVYekay8AHOnFBtdg3sJfEfkAQNNlyibX84A91FA80k1l0H
Krt7S1OukYBY2cqj+0uErsbxvSn0XfWJ0GZeZBULd14KbVAdVDuwY6yVLLd1YGCmXzokHXzvCuKn
UVhMi0H7XRn65q+OdemLJSbcVcHpVqHr4noM3D9DegyeSjuB+XuAuzuS/Q+WUrEh5kQv4QMu8Tdu
RFf0K9CvuD5JirCcl6v2DO1VZ8S/IsOs0W08ju+LJmp6pRmdh5ft3JokClIf41uSmuIGX+uEnyE6
tWYPkfCA5mZhFc4sPpbif2TyhUlO2x+/B+7Ca84Ijw8PXuDAqDo4hKNDWt4YKZ6kWCo0uFNMmeU8
8Bk5O8CKIib2iJdV4N4cqFBFc6o2WmkPa2OaPvyol+DlCcjKQHQOJzqnKBrtacV0oWVMTXxSexwb
22BcA+Ugmc5PBovdkiCREY8C7SsTi5LaRCKi9BbH2or+uQSn4N/vgkaOKlfBvxhdb8coavBll7uZ
NODd8dzCwJbAVYTXPhtpgeQuRDTnlGnSMiKQtV4GL/Nm8RjGaUH0dJMmatHYuwRYvwFQhm2D/SXh
d0nvehK1VlazkpUnNZaXXPmMhHpBvchaujEbLslOEAqMbzEQURLDso0ijohlAdE8jps2cZx75ROi
SWcavQ1pp8dUS6WQQPhp8vhIlGfFT0PPAQopjuGRGHtdmKsNswi7Z4yBj9uETIYvEh+bLm2EN6p1
UvUb19hqb3ji0q2jsnxSYPttcpWIElVCpcpsnboeY9IrWPG7YAd6pXRCbLaRc+aM68k4xt00qM0q
Bad33U27IJZXtK79YkMROo1iPnU3FD5lLVDX2yvGFEXKHkNgNVU5BB+uhe+Evleyf+CaIMG8NwKW
2ilVnOMJCFZCNJIlVWUjg1MXa3JUtHC7UaA/8A2NyxrZZYEWvgi+WTAnFd6jTUwnWmjOZsHWZ67V
aTuhZ+OhGwnda+NY83XOgdrDyWnKnv+y/Pgj5N8KWJUjJdACGyExEgbCt4ygBswyyuluwJTBWBZd
0QeJKtJrIMEgMq9vbWepC3dP0IQYVVhQr+dEmKQdURLzlK1xzWA1QisJxWtXNVIKTP8FvP1cOFQ4
kpz/VXZTSFAFUN74QD71hUBtPHbygFLHXMh2P1OOOrU+8pmFd2U1LQEyK8kSUZy8rMmpr1NpIgUd
zpSxC3gMYoWogHq3v517iI8tCJSII2aTxcAPjen3gJRiJiuZ04BaXf4vrZqDjHFrl3o8WFQJ4mUN
qTUt2UrkcvqA30DZxj8e+mn4uum5T9ANighxIhHqHRAmeEViBlPJrSXSX7mM3jACjDOyNsja5kil
mwy8Lo9LV19ytv4Bp5iLb4VxxQZO6n+Cuh0BD/yKpFM8r3HbQcxkHm4PQmdGvHYR3lW200RNmexI
Nx0224rYrQ16BoQrmFiJqeg4SIkvLRumFGwYcEBmX0NeiA2KvuVOTB6rSHk6K4QfY39Idfrqd5L1
AnLqzxz4WQL/Cno7vl6OUhkw5RQk8zgZzTOs60o40Dkc/bX2Z24d4yYpq/HqTMB9sRtKezPazyy7
4roFTiH/erjfGj5KmqHXR6EOPSRIztVaUoE1OyoFlXxKlqxTCNIPfJV8AypEWNqb5G4b+3PZEQR5
K/bYJ0dAc8FsW18mIzxXCOtXmjT4e1hoc41qJ0vnOI8c+q1dmZyq/2JwZXZhCgEjSZeWnby2evLB
pceshCBlDkxSd5pt5RVKTiUvo6l9chbM0Qua33XObC5gejVhNTRPzRlT6BMA/ED08nrnGLYX9PG2
yzKsyLs4EepBRKUCjRM6CqQSoVxYrGMSf7rU8iNUmKXhht8THGU4nSF22cWWMF2aQgg/xV3/VHrQ
I6B9UVzRK1XzKD9uWqBdIPJJVp3AhLgyVcFbD1CUMqyKosCcsixnn2qWVLoOvslw/w9rFLIr0RXR
TQs6eNjY/CnjJKKyLM3cz5MyPDWFesf4RYmV/5Z2QYSTrKSFihzFtnkYcRSZ5rECI3cnTlFxR+fp
9+3rfQ3zb4DPQqFfyVaJLI5PLz8NiCAyJ3Wk6OoxcMWjkWTOmngWh6k2Hc7Ien5ZEPJMQlJitgGY
fddFxEq02HyxRk9Pk5Ai00eXUqjyPP1iA2mWSu+7A3W2R/e21LWmThDAhvfSn6jd0FpUWpVAL82b
mx42zv/4Fwwbcv6djlg1ZxQkaaH+jDzpNNajW8QMCwbFseuWbTV5/v0v39qb2D0tljKzaEGypHCw
gWw4Ty31WWF9PYVuAfPOHR/oAG13hyLyPAvoek0AOEpG7wP7DRLGhNonXYolblKOiFCIL06dJ69t
VCPYVPdZGTwR/KML2rorxv9ha1rHCVwKrtOoH4odO5AasPuOrbhDi8mH2A9wLftKB5BeYYNpZdAL
Zl3YextV8lbwgBxQiPFkTGFDECBCyRwPN1BoqFIElhMhl4JT0K8ETSobPRcUW7kspRcitAjl0ZDi
ybdVFnpczm9SS0jrhUzWSSRd9vCa0TeYZmnEIcdsIxa8pkQS6hkimzYl/prsA/CA8iUOExb3vB7D
sauQMpI6cxryoXEzn8CNvbFOpEQIdWTvVbpZuBoMGItg0SO3FUiNcUsSNyOHDWPBuYYCmfxLhdcq
hblfJ+ACxhnvf2gvHdzsTGzNZVTgWja78ybQCS9uTPpEpYkCp9PuXZEP/qgy0Ws1tE+OrwoGIEay
KqK1DLBBUuLQ3rDEv/6FGMl2p32VaQTJS+6V4dVBwQ3RfC6fY6697N+gZho0ARb41DXwHKAB/HXD
1D0zxnYgSBs3TUZG/oh6FGndtAwOQClu5AGefHItguqDm75boyblk1qML3VUEKm8Oq610cvzMqdQ
R8q/dwTAsHlkMa02zwdTAXVWHyx82iIYsZBfPPemdGOoOwH3IEo24oQ3iWS1/tAwXWh6LAn8Uwfi
8v4/+taOSL4L7P1GG9TyMlTcvggfXjCb+htzBZltY1kMP79OaXGlts0FwdPWbiJope1eHzManyxP
/9Ri3C22zZZPemhK4Feibv+vKqYfwHIfotZi6RiAe9jISK7p1otP8b5+a9eUeBao5L2Mog0+n8pj
VSVS8EmjLXfEM7uNE4lZwZirr4iZhMxsAhG+aId7CrjyXHVlG2Qi6TdVhb/vq6NLtj0jqxae3I2M
gI1+zGS2xFzEoR/zyd1fvHgU14j0TsmW0w1Qx4DY/QsyDG3Ou9KImVzXiW1e52bIobHBN0uNNSxl
h9Slgi2vEluV3+AW8U6ic8dtJ9O0r4euPh6Pz1pZ+aS06aHimsTbQ3QKVW5DKWfOa2cWNhtZMm1G
JxaghgmcDQW6oukvZEKo0CfCwXdUsfpTcgtopkW7Mr7vAig8Xa2MP5pmdtxrIApwYfdtuQ1t+csc
5J2bseC2pVSxAO00em43688MZw8vwCO8uDCcoNUa3NjfTcOjjNr8XfObmFKDC0ZhUPLghD8FiMSf
ZwZh7V1tFB5qKfxRzt2C6YOnpw0hlK8fmzFagjDy+FmVOLZW1CbizP+3HgLwQlsnShE9NrUumCK6
HKeVlYlvS8vBYcOrhpkXnjkrRJXSgev0fViSH6XdfsZDQ9eMQEi/CNZt4qPFrT984yhQdkU5Xkl1
4Diiw8yMHjG4n2NjbzGRaOCZxo8avFntm4yZFXE3xuFaRnccABIKIsmTD8jtz9WaW7yuutjtQodN
Cq4s8YMTSKXIi0xlQhfCo9RLaVe7qe9+7CEaQ0Qk6eSXVId3xxhsur8dh4F/z8jrbQ6Eq9V5IyEH
e5O8/nAZOQARU3w3+Bsg8rqvFFgQqLOIUU8A9aELb1ZLYrtnGq8kGqN0OxGZoLD/yOgDu0wYzKtN
9ZMfBrSZEDkv1jTY4vVk6b9s8x+LgGfeK2n8q0SdpWi6Yx34tbVEmn3EQEhnZehVobhB1Ws3DBGS
qbhh38y2UpKhHFhJ4gFN+gWGJZNa+siB6XrsEnc0qOT3lJJ7/D280qRFgY9mmZYjGMZGqWhd6qUg
kjWW/2X3Re61tKkLsvWrpieRGKneEEm/S7yYVU+GoqhEcPEglSWmPoXfWeav9bBAMgx2CXjbkyZh
LwNBnK6ouqzt1J3sN82wXWPspIiGyfFbmazIwYohsvHRXqRRHGQ/eYLEgZY+SpkXzZWk4lPGLDqD
T6HZYXd2rlABu329MUvI3yj5yDbWSFBSSb4pDCPvBw2Wqhl/45shM+EM+gE42zq9WyCFQo2pwscD
Q9I6/pCpeF9Zvzn97BvXLs9nrFugWQUMrLVKDdtJXBwhfF0CXZPkisL05Mm9LgbEPyqVCRnDOscl
IAZdz50AQCWEG6/5GtC/o0FSiuBUEmXNyQWdR/LMUjPlGpDjp08vePargCD42H4o01H0f14RKJ4+
q81lHOvDZZiLqwm5FuMRpE8gwJ/OMFXdUyIMcKvdgWTrdoB6/ScBohb74ZeTuzTNah7+L+FaHgOu
IqEaKCLwvGLMroxKQ4mpX2mNOMHWjBXDv2v1mCqZzq5PQx4tCcS/0L9xJpQniD7egBiVzCHX2jXq
KDuj/z4iuw01PHO2nKIf8FKvgfsNh8BApksPhx3xgZNten1o2xWZ8bniCdsV5RQZtRdU4O+fa2Aq
KIaCbJ6aoHGASVTMlk6VS3dCGy88aFA83aUUAz/0FcD4KwklZWdExyVCBbNhh+bGvMHnWShOoPuf
+QNi5xynavOp1iQZ6bmNbrIFhUoBD+uWMiWktBtN3KDDCnw0HOkvqoRmI+ld920fr5pzlJwoxwrE
/9JI9+rVofN6olSyuNvoXtG1IlKC5reTBp0s6wVO+xj4WI2iwBWx6lqB7MWqsw/ksbAS23GBN3+K
Gk8Z8QjbWZfuuHxX/KdtdjtMfjVwVE5tTzfDyf55HuDChkflElpwoxoDz4CKJA432WSNkTk6XNsm
nZXzJdJZGmesL3Mb/6rR5wU5xZ/GOHJjF2n/BiqQclrUZmawKZqlbEiKH6gdM10okcEuI3ZgG2G3
Se5zDevpdsULehpGTzCYxZU8lgWreJaWYEzgblzT6UJc9M33unAa/AxlkGojbGIMd1W0yeB41KSS
HngX5xaVjq1+00k0hCyvSn/yp3GTQPvmkBX865kZtVoUXVBnzoLi9PuTLDYmaaNCGYdLweBihlfv
QO0+exWITDjyXRf2e0GN0BKH7zLmLS33FQNrgpfRLHZQWxUmAwXFf7LXS1rzzCWzmSpBHZkQNahZ
ta+mkJhfTgUggV7EtqA6e2RmpYV5M5AtcUnXoCiXsotieBSW9cEj2CMi5hUV6ennEEt7oBtyy12X
xEdE/vvHqATIXK7HAz4uL6KGwAI6XE860MddcZdaNWiw2eceNxrhpx+kFr3RxKB4Jg7yikH961bB
KU/My/tKP7mg2zTyP5mQWkVbKM+BGAdjD1zKNg5uSe1QatwuE7gU0QyUrTkmwHMNlRe8HQhYQJ1r
S5G3tTEpKS5nhpgFYF5cT3umuAAy2QtMiiBBJDLA4vyJjZR6d8C3aLAM5z6/qtTEfUIFfYu0U/5A
svTSuJ9iSRsVk1yQgX53HEHw2J4muum7avcwMpNvxheh2dzV5tD8egH5YLhcq1tr8gs7hvpjlZgu
vT0XQOJIcVOPW5SmUWvKNww0st/Tc5tCQ0Birr8kQ2d+TnIk8wCDpTR06o6UAqPJytkOxRpNEHMP
RbdbYAEtQCJCHeZl5noIkfr32I3uqfnzBYHrdAe2Nw+zIqg85PRZd77i1JpmNZPz4CZbXWwmjmvH
pIpU8RRKRHQrfOdye3/yWLAtu59e4u5zpI9r7dO9jhmQKCsVNx3NWErLWO2AIrTi9vl7WVcIwXsn
h4qZr/zU43CveIJCK9dW0fTSvbYrx576jBHGDzP5VFvkHTYpK/yzCLsW31knqkrDJa7fp5gfuuZN
wy/VMy1db+M2k+eJZmgSvZTRNVVH0SSTwp5Gaw9b1qs9qaVvVTWgdMkvyW7u073Wicu5fDbExf+/
Cep0rqbxwEfy/SN1xFKAInyRa6CMuKx6LUFssssQR8HcooD1k6IdsoHK6iBhO8wDVYwIaJc816Ws
PcBVPiFA2zoOXMaNXBxSekTi3COUoA2Ti0TlqsglreNRUNLRvrGzKnIwp8UcMT7pbvdRnJ3SyqmV
swc0F0LzZ4ngV2f4Np3Bn6QOzwtxLdh6uCUvCrGdDRMqbIICg4N10HuRUIb+/2yPeRos5y11Cbqg
7e32CHC6dOTlC5liqzTxC7O1MvRsA/YUoji4tzBv7dvRT5vNskoi65RetaMXY6wm5XqIpAURdOL6
Y7Zz4sposu3YOlgeroifW58/wNp1YhKydFwOoDa0EOU/DhdwYXFYC6TgkndHUtLYFvGkZ++DY9Kp
Ta3J6sHC88OxO5EM3qDx8T+zJlz3Evl0/P2hi14WTyU4wpnaluxd4aMZU8b3VNUGw4jrY7w2NnYq
21TZJQmVPFVoh005EzhwhDS1fbyaWUZ2RhZ4hjyMvNxdF+pbPvmPuo+GJMtQwgOLogZCwCx3oM+U
WNI8zO73mUdk/JtN0kin3yS3bMAFJQ6Ghef6jEZkaYmMYzT0Wpo14FMvYwJW6DrvU9ZRa9FtTYDu
KvfojaZQYO/7sUX664PX/nNFa725bj8nl0T6NgId+TXPzFxoSngceRlQ0kq2obP85xXMJcppxlez
HH8CsW5Hm24F1TQ6YprHKyY0djmBLE43b/i9+RH0wRmOpJLjUmRA1I5KMRHK0yr5fDd+2JScop5g
ILKOHowDriOc5K2Nr5LBNK/j7nz0poIox2dJJMBHK5mfnbQ++0RSJRPNYj4gOx4bB0iP8KPAr8ul
vKFeuKT9G/YHTKQsq29s8OIaTN2RaSk7BxWucuoUgwtvmeWs5RUfVhwk5dWfx5UOkVtQ8nNiLg1S
l5Ps8pqeToEhFh2AK20BTqExCcrEbP1SFGwrXcqkPveinVdOqk60tIGFO/SN8Z5oBDRgS0PP7IpB
WV0lbJhJZT1PFgK1l5dWR/WiOMJAAGIdbXWlTboCEKShXrhpJKA+Td+x2cNfBXyyBHr8nSGPHHh6
7anEnkPkzZHUH+KICOEH6IdM1gENjjiCUljvC2KZsQeHpUSBF+w8USCzOSTYd9XjzlqWAfqg8AaM
+hr4lj8LQVHYC59qGmz/rzVEt5YjtE3wR0qHfWFQb1m7KQ9Afkz2lhbBslYz8wQMvAr71x/ID9f5
+nPjEtqlhLtWFEAMmYzcJM0WhgqUFRhTTBb9nwouHeBkKM9F4HLTUcnLoeixP//ghbNLYApePWwT
pYMfbFDf9UkYj9zoGJ1P2FlHvHLvvvHb3++bDB5kXnv9NdHA1t3JH8IzFmWeliUtMhEQ5/MU4JZM
C7N9AkdCepOclXHkpDCIKEvFQ9oATM2JeD5qhxUOuvY9EMICH5yvec6fGAS+XShTx9SNylsu9ars
sz3PtrJIE7ESec9LVXwHa8l20lHdIn5gkWCS6O/fzXgM1R5Syv/BzkFAE8F+wEmEYm7uc92ZYzM7
XjWM+EuIYq/fOXGGWDyaQHt2kOWqCzjshdn/dstOYYkTZhDvr9K6dsNPwMw1TupMWOCag4FtWtr5
b+lWGDHXGVGr7q7k1QiXBiHxYHku9rgAPdTBDOgzXpiKdMkt5ZhLEpZrL/naCLpJxf54wtr8YjdK
iU2+hrmSmNDSXr6VAB+Lpo+QOAV7g1dRcHiB5wwar7np7VKQETwsI6nN0qTEeaz0dnqDG7jUTZMn
2S3/izNUcpdjeo+qavzuEPM0hF2KYfwWbXPgUSVqA6at4a9j9893YEmpZdUZPnTHwl30wztGSZ02
qvyPb/XzKr0D3ztsdxXVpqkjzPJRldAFN+ebIb2p/M/AZTr3AhEGSsIN1l1KNamn+uZ5ATVox3Y0
NEfyGBgC1ruc6Y1S7mgUnfufXLo2iX2PUTfveQrpcKV8sX86OZmDCUzMY0XRsC+p38FbYuhy40yL
biPb5ukTmUHQ37aVmm+jmPmy7eLPzHLzdgrGvT3xMNaG/xzHd/XxtWTqVyI8or72qHD7S6bkDire
HS8kpdRYdsnej53oFo0Pk9BrHFnnDCuWsjJl+cAviQCDQ3Ec+kf+z42drWBbaeSEZaQfFfbiH+sD
6ESPa+0+nH/olpdvFce+zg5HFrkj61tn6rlYBjS0qzAZ0SHSsd0SuM+ajjb0DidgBEfVWV9Goqfx
5YYMLCyCtpWdDxaHV2eOEk5v3jaGkBC0AzlXO5rK7z+pspTjfFosJGgGO8JlO4Hc4oKoVJS0HZdn
ToznonU6NTL3NP3jG4+nYFb4nhgtCvCSn9cS6D5D3+SjvvsLiPvl3Eo7KhgME2LSJtpOMYboISYL
9mDbXmRBj8npzjOrCcezsBmVkkRUO1Ni/JO5fuWwQEPC5w6i/qHDG/QTT7Ly8lK86jkq/k69DGEL
jX3hkXMBUdgcNWa+sGcyjRSumcyJ4BAs6ItqV4QI8sSm3pYnafDum9VO/2IFTTgjHlemxray7Csl
CwAFPFMG6kFhTyccvsBmPEDlF7cWUzxYHFOT7TZkD5jzsVAqoaIATmq25Uco/rIGn1vjKozrITV8
8kRjN+GEzUQlf0vFBtkdUp2sLnWhlVzFIU2cqdCehKv+/z7ZwS8/f5Gs6+NJvOxKkqjvlpE+6HwG
q1Z6srpllx7ziPKqLT9nlxc/jei6wMBPhK8/ESjIU+vhFIemb7cuPpbmlJ+E2ZTrlyzOWK72uw/n
T4sPQfk/BIf2I4TA48tyraAKygqZ+fQsDnw7gO6sW2a5wyJnbJgtgdsgAtZShYCMQtiFRcSgEvFi
Q5KabNZO29BH7flS7kl+kJzA9yeSS0MU9UEcNKWdaPyRTgWqvqcsu5wvmxE56/sPJz3S2M70+uW9
D5K3JXekiTxIan5h8JSYXZLds8OHDAuGHJrnY0f/bjzIRmCVn8T0KIL4t/DEGAkOVgT+24l3boq2
lZ58o+RX+2zhUOUwTfeQfLpDSi90I7uuJH3QSYv0DKIHD+H7RX5Hnfv2uDfBONh8eg25GdDXnM1G
JU84DI/BcfwXdYRMYHEPxrQX+VewR4H/RLIpp6YT3K8vZj76/y1VxZG240tRrN26qzkLGc9Efvi0
M6ZzFTxFwLHs5kXc6O7Wgl9qDzOoPVCsyiGI11d3g2kv4ms+3MqOOPgbHzSvncx9Brv6qUW3G405
X4McfLhJaB93qkWnVHTIA8FoTGT4Ps5skeiSHqQ7KxUS+T6kEkbyf3Fk91f2cjR2cEFt2Hr5FlYr
jqMKsgOi7X/RJcQTSzGn7a6cyevK/k7eDipPYVrjxx/jC9en+UGW+8vV1+sf96G7+NXk97/mLsWx
FsRcbELf1Q21wEeB5q2d2t9X0EoBtQ6T2M8p3C1hy0zzUwVgLCauHQndbBhhL8HXtAYhKfqsR8Ef
85Fk+AfX37F6YS52AP0/khpNRQhjSk6y2d3ETsa/5UxgcLVFxN/GHOSxc6vFCSvvOOXg+dzDMh8q
vf1boGqm7BObEoehiouU3KxH/YgLBFk+YcjakwVDFcJpEGivv5eYju6MYC175jiHtnnvDHv1hUZs
fI1ijlzh99G3NUFw99ECeJP4cvSlLyIy4SSe9MdV9Dx1VuJ3UZQiEcGgolOp2BXCtOmFB5G/w8Up
SLNO9Vsr6vrOggA/iaRrVFIdyRF+XaWvQTZXqzp98NBfkppCA5oYYrb5D7lHGrJyQisrgI3K57I/
XODkJsDCSbdKVQTDeScld4euE0LxmkoO1aKoD2/rnfxy060zRy3ZdtoTM17etBHtyzL6d+jio2yz
6WsOf8l9YITIM1mZuOQXagEpJ75s1WQ45WeA3FkUzaSFrJoqcTw5OzMMfJdCUG7GOURbLuPG6gi0
z2wOBIu/jnjv7VBLxDxY/5K9si/FpbBBsmQJMrtNdEtS7AIsIyLzYeG0bElFsS0Pw2LXxm3bzscN
cWxDjpT9L48io8hIZDzY+NSRdPbefyyOuaK8PR8VluyCpGUdvCuEzvHMqui40FDlLuKhb5gjGH16
MH1dogYuKH/oaasCrCEnKtEOCwGN+C2GFyuFlOzgV8vJRaqMIkQjACXJWELC7hB7CSeekgTbuZcU
k2wf/c7segayaziffBsEiOfh3zaIK1lyv3XjoqdslIWTfBYAjjaPQ22Ojt03dw33WAX3rqBJW4tA
FrdUWUZIF/GbO7VGZWz5JOjv+mPrZ07nJmBQ2KMdJMGAYKss0XMvi6esgbu9qorfUX3rVcu+yf7b
N5vIUxwwf2bVfqITvzc162sKcDSOrViJgKpTsa2mBRIlpbWnTLz5sxSZlwJFUfhZpzAkEQpqlHjV
PiV+5G8wKIFJpQdYllu+8b/lVp74FYclYFFpYqQLo6Z3YODHZs1F71MUNJ2+oDvUyJuZtppCHMdb
gQM08T25mU/YW21KG/gZQq1TVKK0qzj2fnV6S7kcQk6+LnqwJRrTG8S2ll6anJhVtOigUcW/dxv7
fPhFL21654fRznXtOYmnrUckLQluka35LVp633Rqe2I4PTCjHcWgRb26qJfFeNz7lswnZ37fvN0w
d7tv9jzVbt+KWSdOPi2M/OaU2S8CDH5s27SjRWwcBO+s2XOsJe3JED319t6kF98vU9HI+5ZK0I/h
9xcwJkbi0XXmMgQ2NllKSRwcHJ92LbM1MCe/pgFU30OAtsWqfd8pATpnXC0IOaoC31lxQ9iYx0uC
viGO0dWRsjrZBAtfj+sm8IrSEfp6KB3E6Tcuck/QcT+xgIdYT/P913n51S+nWVozZL1TMvPfnBli
Y3PdQW9YCAzCH0/nga3rcisFZNPVuLJCuZelR7K7X5hENL12SU1oIONRIHn6jXDFakNL/nRrUyjX
uQxiA/iNf///zopnt5Cq9t84TCh1bjxzDboRLguvJiObN76YGJ5y38urkNkQ3/qHBloS94MfUAr/
GvfIijYxiLcDkoyf68RGWHfpWPyZIXykiLFL9mQu0J5GYXSy6lDrHmNLeLn1ltkuZ7XQSqQMn3k6
4ct6Sq6iWoOHGJVk4XQgbtcJnCEy2znVX9rrlzLkwhBq+reqgABDdDS1QGVAC1Yc+48SaeGqEb2W
7NdqZ/Hg4jjQmons9/CQ1hg/zcB1UvYW4BOwMXW5cGo4lv5oN2VGrFzNI9LYsKbZ7X0274yf9d8L
i0z+cS3JIaGy3U8+SF/qjHla0edUD2puczyrMf8YEfpAW4kH1QSBiHHgXtiy4dmjf93G6DTfA9J6
/4ol8VnH8rdnO9iE6UrhPOPWS7YFpSToyGiO9cqMjt1Q+QwBMe4Bz+bLYZR0e2MjwD0/IKClLCNX
rYGX3F/fK73pca0Ont5R0oW8O4Rsl2OK9QUs5elze4ag00PBU0GVoJwINu9CVWmr6TvxSEHHxh5+
Ai31IgzhNUtkXsInkhFKsZGQYm4zQBbaWkXIUOeOqHPJINaQ3AYDnaLRsofUK7b2mI0ZKSGlza++
FUjjoO7jHcJDs07gYOjfvfFhpxO93qWe0wid4umgXRoRh3KY3TTN0P/ZGGn8fujyaXrD1jSjs+el
HvEBCZn2m1+7G/w6NALPBLwOjTi7GfExt9x1f3df4z01vsSZgnxYCwrvt0luD2rbtFvF6ecm4/uG
Zj1uoWK79NmH9HCV2L/kljaduS6PqBG/Al1cBdqHQp5ODHi047h7ld0ymE1qWlPzyfRxFDIlU8Gw
1Nqal987EcvZIajQWy0b8geAwKcl0mpi/bx788DYK66fFZGDhRwkXSNtP6IduGvt2jvLSiXCh9xO
EdRSXaVboeAwFFHvTsxAlQ+JoVDoJVWSg7NbKNAkB1+eRb3VzVRJBaJtdHGexgUWUwGiUMQ6rFyj
giJeU3MwbFbuiRMYnLbbwt0fF8xxWEPHIhB77ZhPC9q/CFa2LrypAhgnFhRU64LBwtCmECEWrmPR
5Ewalsz2CaFoAGjfxUsULs82o7QcUDb3OsQKMp9CtzK3iAStup36PgKQrBKczZis0XT+y5BvBKnM
aK3BADV8fXNjErrSfQpr0KIM8Yip0ShzVBrvJXFKNWHgfhrGsNxh9/UVoDp/aDVqgLHaMUcEDE8G
snA3mQBgijr8spo9sUZxzgDW3ziMdac3+d8AjDrsKwg8cl4h8zjKWuEwcLudgKEaoBk2DPRizDRz
juKnkqvi+Rz8szGPIXnr99FD3bqvyh9n13jS8ggdIsurQFgSybfO77S0rNLsn1eCR5SzW2tKZt4e
KMCoZ0G1UB0vVN7kedUMmOM4rknWwJxCSLlPI1EEDkRTcXlJO6wSB4w98de6+hENQ0CW/z7h2tN9
lZw1ZwVFGTikjcKovbi9asd9mB7OZPeCG+ZrgSBQu6fbFR4dh4YaEGGM2nShyOpQQI55QM+Pp23+
8zfCMLAZfty5QDpncUbB8k5FlptebtOtviNhwQ/NefD+qFLql+D/68TDfk7opoKlzMaOClJnlMes
cgn9S0tMyNGlcptzCwe+lykhAeUle2GbApD4mVlP2hnnR5XV88/5hs67PuYW2RISTnKH/szAplJR
41QyvhzqXTcBA6/QulBD91uMZ4ywrG91uu/oQuE+beBdv8YKnuycEC9DCXbfE+AlnIcYlh+H6Rll
juMKwHSKGH+5e9/w9d/dmUwqpL6t6iWG0veVBxxk+thnPHoDnJGKhT/NZBtmaNUbUA6MFb6ymcre
OnzPiJ4B2oJ0+6QO1o5ygvQjUB1+rPr6/KJP2CsJJQZ6ogwP4D/ky+hI2dWJYsjLaQquDYvlu/Cf
JTTL6AvmKm2HBD7Hw7rsiyDHRm/C7MoxwIq9Edq35GPzcOyFxCgF3gTOp2w3KiYY/YJEJfBfnxrx
hZZR/iLHZ/6i0UuExV6buF2yaNw1ckS257/92Xo0Pd1Fb+Idi3fSMLBBtrmKC4jXURgdayqcQP9W
cujHSYLuELpzQp4lxnsVgUnwl1MP32YZorwq2y0KWchDtgPdeMsOV+Vz6cvAX/8sLx3peWx78RqU
oFFGgmHzG05oWsXynknkLOSZIUsTGIZJzUx0sRN2hI9oyTy+8CvO40gc4RDU1HsO5ncrJTF/d6tp
Gw0zIVR6qpaLxyd5YgDa6zJ6eXcjT7wpnJm7jtqGPyOQmCQ8reS7Un7tGP1CWLgrR49ZyaZH3iQp
EOipqGhPx/bFf428Xb1nxCPAC16Nu6BRZq0GmAitzH/WIFif/qFWaN5Hd0eEJcgiM94nLw7srej0
uRD+thP6DSfhqsaL8sjSclGvU/j6Z+N6VlsHuh67n9IC8klGlzB3G2V0K3mygSOixhyzZ5GZYRKo
ffkzM4F8Eka27Ik5BHTlcDeD+r7WQmt/is0TI4RcngqWxLXhNniE9OFIpAsd3gWbOY7S8YbjRxXk
lyCwFG7lyBZLzNb1hV2ZXIBLsrDxHeJNDM9rkHnwlpiw8F78Q2BkqOu89yxE/FM/FRdh3hDDkwI4
bmJzEw7X0H+3areetfese6TS/H/3SsI0DoNyKVb0P1e6pIZvyNbjbOIUWfKRi/gHI8r20n2/XdeW
CFVojqLFTeWGeppHcxtBYQUsm+s9NBJcSPoZR2pXOpBwAEH+dqhis1fFNBOC4VSFjjAMtRVYifL4
Y8mZT/MgnZSjA306kzkQiWUdhoI5eJ2f4F8NL++fZ7MWbJe5823QS6NFNTDDTE2TCwNYXNl6jUGc
dyvB7DTYmsGDy/vyM9Gz22zACcDNtZOj5C74vt2aqTnxEJRzErZGIlDfzgqqBRQnf/zlCKe/C24r
QVaTJSuk13xJwW15vUgIP4fekKlwELNcUZh9a2XqxiHB7fU+a+uelH/ieKDU/ThW09X2gNaDMUxJ
9fXJUPHX11qHCkTcEgNAfL+v2eJJAqJMYZKNoj1lBM3vTZ3sKjetsS2os/XlcKNnBkfomfgcwfWD
n1mIFV73sJTNwp053ftE6l6GrPDrFSNR0i1PX5auJLd8ykwlH9SYnpYWJOy0HbEjaZrtFcPspHfH
BOiUDvM+hcyjfycpVjgdngNnUnnoZuNBLiTPIaKl0WCPfEKyTZx23XSD0169KiUmh1oCI5YZu+tX
882essyLNW/sOXQu1tnuKJqA11wUIyrSOMjtO0qkh/GfKJmdkldL2erGErWZ0rmAYrA3LRCjQFY0
L3TLYh9wDGypTsebYR4h/AJq56TWdSKvOMkosp6H5Yj1f4Km+DJ4iFK7C7cMrjfUD++BivToBG8K
qeXr2Ty7zWpJEM4rnOm5V0ViqQE2bo5k9vdMut15fCjsywkvd2AKWxdc5lu0VffftZJbRdf+jwZu
gfg+zq3B87ZTYvxlL4RICDb3/ljBoiei8WlDcBse+i0yEYM+lX/Ms/VfTQSQac2RCibhkWCAI9iT
UNagQBq8nh5tAses52XSPU4dMRtq1irDGmFudZl0YEBIELN7+DYJ6fgN6dN7GYbu5YZzfk3mSSrR
Unc+6tpezwYv38tRGMR88FHJrWuJecVJ1j4tAzr8j9WDYHDX+8Lhgx+JxJjJ3F/+XysGdxRUV3IM
ZtEiveJGLrNHdz+XvTVM0WSxFMhHE920QOpv6EWMkn8kKFfj8D0eIWmW2rmnqkDhkVeLBXtiCVS7
Wwo4dcTOiAsa8zaKCtpR+1nRerstQKxVrNAtbIcc0k33PanaIsLDvq7GTn46woEMM1U9bl2SuepJ
lyKkOYh4ClBs1ICWN9HvBBCojYWK+hrp53+nBUy7Sd1Otn0p1GoORkr1VCS18ThREJqbWV7ljOWt
XHZXU7FZd56nEyy6NBv7ROdAK55QGrpgxqhPpmVI1WTwl4ZBxyA9Hx0h+qoY62Rt7tY0GUzZhBeB
g5Z8T6rwa5fV2Y3NWF24f33IiRH7S0wEpUZP9V2oi2F1jjAwB46i3qCYVby/zEgUQ08CJeE6rhUV
5seM4pxkhfUqAWqormHiLrG3T1we68uxM8KRHEKYGOoC4bn2BL/nIvKqVg2/6pV+YwEOsJGxwRXZ
/Ct+2ZJRn69bxoXgV9lkK8zVfOIX/PY01jUNyZp8jMt2Kf6FtL2gkUBKavWsF7D30hPvbBXgK3LR
oaQj1QObNA64GZkQ7y4lkdvM0IkFTa+nrLfhLpylPfJzYuqr7T0jZz4u0g1VyiGIMz9IL8YeXSiD
1hyT+7OxTOiAMO0O+FJmP21uGP4H80bPjiasmE2xIz+F+1CZGB9VVcg07CRbXU487oO5Sxqt9rYA
f6WapWSi8NS4yW9hW0dEVmnq6sFfaiIDGGILWvBpmGr40mgN1TJKYnD9D2o0Su1CCJ+Pewd8lexC
/88+YJA2eL9b/MZl1mkGllIvrjQFT42uU2N6tBhE470xPq7PD8Nlbj7KDPCLUSY9yjU/zw7emtDq
EwuhoSsvHfdv97SpPDNOyjgNcRQraF/HRZaN5bbb5sixAiHlSlHaTnknKt0q9MUmfKQqj1uVaFXt
S90W69T2LnA3E3GxLh+nAURpBI/UXc5pPxkcum1mPnGpiJpGMU94tOQKB/HYnCN3rSJec0NXlGlY
cRyJbk4RiH8Ju2KEpREFWfzfHhaq15ej5zmcK2I24CWqiA2a9YYxFvXu06tYnoucKabo3T8TEULw
c4Ce3WFRQf8hag6IHl/9X7MVYNtx2gxoIB0P46hb04UuzjI4ly3kBS39A7FIjsFoPz1IgYVx+Kqd
WQ1kSOiBCgrk043NlYaqZBzQinvOIhDDY903KW339Uyh27wqHbbNHpNjBuYPp7hhNvIGHf6Fo/eS
ULKW14s7rm+pcgkSJM9toev1XNKr1YX1OmPhaz/JrENF6hRXOui92jn0RZZM0kmtyg8szkCJKkyG
Du9XDI8NmeQ/AbaMwrHyPW0qlJViE61GmpIQ2YGUy+5ldhkYGSsu4lkuw5gnt0IjZpca72C4jcPJ
6xurimorLEhQuvWrW+y//Vbgs0y+XnEG0FFubAgCNpbLtI0LGtQsoH2cJ+R9JXQOH+ubPp//oFz1
QAnx0QcpfqUr3zxK/Ld8cYox3JyA6TRVxOS2uakVCbuxGnPza5/HFgQ3v4uMIRj8mp3szesUwCJN
MAb2TjKwnzoa3CnOYgF5beNpas0c+IHY8OYmkDht4fAc4+QL+t/X3UqjB8OFAnvfp+BZw3pAws7a
qAytr2GC2+TCwrDBavjWuSQD5zB0xmO/4Vj56gNoWoZqD0wKAzQiTtHjK+/qe2gJxWy/o5o2sUNp
nB4jjhZQLJdzNthZJcUM9MsgXRmsJ2I7RxyVOEwR97ZoUzUUe5pRPBin17l5H9e9jyMKpPEmbpFs
gFfJ5VTL6wSPI+u/DHDUzg4GtwwgqBV5X/YHc9AVm5+nSpD/gJoO5sipGXCy/O+Y47EDR+E/prJo
FAvL7jTU3TO6Jcu9qe7pirBJZ5HekHT36SWloIt4Uc+kcYpzFvdTsQ4WqwCHTuK2/Z9aFawgEEeS
RLnkOjx/qSwd7Y2dM7Mafnor4gNvHmtHUhcRUsL29HQCZTJHSCR+wWtPQOmuLGvPyAGPcoMTPUBA
kus43QremRotFEt/ZEu8nkcD07ElkKwsFlE3N/TDFqI44clt+wKIOlxccFdNPBb3txzY9ZpEqIL0
mHwtl5JZycc+bbpWvbvShBlkg5WUIhv+plhvkssfD9d4I9gb6dyDXoQoHB+576LItHsCVFfPb2lB
jmsFeJnL88qsU+1t4iOlvhKePmp+8tzwl7/AZ2ORN+opUmW8DxqssKDKupuJo2ceuX1xjVfQBFUP
XD6RSjalSDp94xWklKGD3kEUjhpelmTzM8O35CEJkYAsubERWy+PBIrp5qoStAXnqJHVl/o/TYZW
nTQbyevNgE9uTlbMIpJVTd6VdFq+7NrMVn7hW0TlN5ogOzsdEXoEN04TGqspJnU/1/txLnnNRtpe
Ay7zZjAZFtrMXlnulQQVASPT3AlxaiK95Qqiw36SeyiuppwzWBvNRibWYcluT7F8DQVpUm/WgHLo
zLCEI/mqYCnhUYSHoKUADJ57EKq32YZX89bm28SeFhH26Pom4YywkQHNPLqmQuir0j9Wyp6dkfsL
nXX10l7+LxPexhpZjH67C5pyd2FT8uKUuVe+iiWPfgwT93+zw1LWffdahAdBo1q/Hg3OZd3rudPK
kzsVlp8iXLrMesjq18RgIwDciCYqPh+8b6chBOSe+OT47AYh+QiqLVuBLeA4Mm0Yx7RIyyYzGUR1
zCysqrwZb+NUsT24H3GWuexa6eyXfk0nKMCdk+Ks9C+aC/2aICt+1QC2wLaaDPnSTRt8Gd+GMIe3
WlOAYGAjylIoqgj9HGXdbx3pIVnSTtKgHEKBm+NvzsYpZS36kM7QlJgsbazdNHlcJyvVnD2u0O+1
24Y7dR4Y8HAow3sjAN/mnZLsWi7DhtvkqAl7gGkecj4PzwA4hxf86m82FtfFgREXXpb+rvB2OTGx
VIfs0tgRZJkuoiWLpNIYz6IicvQe8jTidd8CeAN4WmK4KMA/RUOXnxkSSzkgahQBdAK549tEA/UR
A1Yvwbzeq+xdC3l72i0o/mWtU+YPg2kjfR+P5pVjJ6gvqx41VygtYEVyLeAu5RuqYki6lsnnPicP
uewJFOdm+kkN3fImdIeBINY785Xn8FsklE8MIPeeMKIEcTtABI2R3m5yONLnGOSDnChqYL93oW6X
mE+UvqET3w1geTQSOMtwe9GcpDGuJM8H8hjVZqd2VifxoiEsZSWryIxfFQB1dVoVozhy8OnrKB1G
eC08L8bApDuejk27SQFa5pbH0D73AYEynnC1Wok3wwVj3gI1b/m40VFC/rZVuYWN3k5W87+guwaD
e1/+sKiVqslhSAoLv0DTm367h6kBQFitAX6Y0KS/MWk1mI4CB6xwBBUwMuHXde5PGc8lIZUWzZX4
bW2s7ZfdO+3peTX0+ebMu4YWejlcQ4gB6I6DvIyB5+QUjGdqIBTfXQVDh1PE7XH2YFv9KnO0+TTn
EdW48WSDJeapZNiixRcylTHjKdwfMpU4Sr65Dx6yXgClDTPpeNpMmNvUNWV3qcjUbSQZWyDIGKMs
AJrPr8X1Rtd0aUxQ4bJEoXd6AKuxa4GE+SZJR/NaQwzl49Sc8xD+sY+6T/RYnHYYmR4yaWyyMJmU
x8scGODfiRvBwwAi67dAU852jiOSbvvjsF9RpOy1aPcW01EiO+avlFmFuEAs8lxaQNTKvLVWn/2J
cWuLavh3UX9MyNu2ru7i9ibVW/S3SVNE5+aL37Vf1u5pVzBY+6UkphKjpkRtQFKM++ZytaWrqsu8
PpsNKodEsnaGD67arj9pPFjXPX/K1DB1aGS9QlKAFEQs3cYvRH1OOhMGyw3/jgq+/Lq7UxsSGlik
VQhswoATs6sZn/Kp1pWe4Hm4IL4fNsWc87JeH9+zpbQjkhAOF6YSisK4cKYssWWjVsMjiDaWfP8S
WvmUCP/uJNkDzbhfczADPZxEeTfL/39bbyjjijfzDr5zq1HZKHe3UoKP/bY1ztbMAdqpRhumIdh9
yfblTnTV5t9llrN0vdD1wGmHMNXnmZHd9NcweuiHigH/vgKJwO0khVjqex3Uu55LD/POkRajbIwb
Hz1Ahta3yySbt0UpXJ8tqxnq+iFuKmbReawXTuOPWi4gZunhYatFHABIdJTStGliV/VVS9B16dBb
cyOjAgmJZETci29IeXOdI5lWsq8RmEqRjlo317oxtRrN6xlh1uZbsIc2W0apOXZh5d2e4nD6VrEO
hqhtXnzPWH0XL9UKcCyR9MMVUmtnIahZcW0T6cpphbLmAx/3kzi96IWRs4JkkscwLntLr4ywP9d/
/YyrpihrWX40TlkuSbhFNgsFoKoR9mnF9/guSdlSbsH/wUuyadLbOrH19i1jAGRWBtDnCxw955Ze
tfvT0gd/8lxDxWQN72qrXNG/9GjfJPsFOxr1ZGwyVR4mkF5odOQpOArUQ2k8vFUMvOtRaa1XGbTk
/i3s492lcHQQ9VnTrHh/PsEfvALi+e8c9kqZUu8h9DcMUBCzYJhnf36VbEz9NwdR94g1mRE/9Tpm
4ri7Mhuh2oVs/f9kImliTeHMTQMzQj5Fh9n1E/dXpvMpwpj1gfGzJBZ1NbhxyDv8yWrUdWX3c/ip
Q050Bp1KxIaXIQw5oeNOuQu3zkPElxJqV05CkOU7QVxeKF2dI9UvzXeirUCR/lV99te/9hoB+dwI
88bCQbDkWPUaHQeCXjB0Nep/WcUcbFO4nq5kT0IvlgN4o3m4YPXuCEXXvZIva18ykgjGsMpvrART
WlN2A8PID31OieQ+yj2xXCl8jtWY9t9M4jY716nHJuUz9nuychJP6LPq6pyJfXg69FeECgwMESoi
OImfVy+Day6tYnBu4slCrGc26zALFyNA99SUHAkPG6mICAqT9rXnXtYPP69YBM6qfVEHQUAta8B2
G4VAsBbK+n3OfWMhGIK/c9AIJ1peMafAlS34UMVOAJSSnDJxYTgRTule8+TGc+sIJ/Dn/eItErxW
H1cWgGns2pSHxddzdlFIX290HbzzNyA65maNTujwXEr/MpMmDKSUvDSazole/mM32868omGKQ5lo
J/QIslVNFJ+Ll5NzOujosVglalwCPZzMlfWCZ9afosL7AYnGsDxE0jDRa24AAGp4/r0gnZ8yT235
e5Ye509KaapuhOOtFErCSzq6M911fKIiLlLubrw01rUx+clnvj4qLTzqzP5XMW9lo1C6j02M3RcP
QnBcIIW0gssvevjGKfXP5onKFvWl4TechlPROTFcpEQnBQbMsO2Djh/OKJ5icmSp7LVCjo0jSkDt
NnwBjjDQnFotbroGkXv2sJl8LkcPxarvOjJwj9XbtJobzv+dHpzqpBq9igk29LSkk6bh9hQmstm6
IrLjqfPwBlNHuhiOPeuTLLRWbkaKAvKjfZeIm9pDS436Czd+ofooT6jN5/Y/bF7WYtKd3Wni+oT4
XT/ombvknWDKA4vDQpLMqDKA/V8etv7Y1Alzv5IUYFfkOAP1AfcEM+N7zWj4dS8pLM9H5GyE+9Mh
URQlx2ck3MRYgyiw5+mx3ZzNJ1ep7OE1ctkLqLqm8XbNZ8z5eMHYhR6qcqZ1GFzdIQc9xEC7seZp
e3kZYtsCJlsJclOxg12s0cz2nimp/hOAmtE5IVs+a22/em3iBMLo/j/ppIh0ZKxYluhcOfV/7UdZ
NZY7fXsqfDvmas49fy3DxuIQ5wu5XJ3QFQnukAMiSlaqSdfhh/s39Ucjt/xlhP7ok4/gPSCTn9HB
HwCivT5S1T3vZZ0rn0dnEC4nhpc2uqnrgOQQhbJnm+4fx2T5qKnNDA3rsWegEgU2YlUPjyZLCC7w
ottVaOieK8jJ+90J2LqbIPX1k8NEAKN2MIu1g7NmS+p95Wv2biSANKl5xCx0CqZ05SVMnSnb3XPF
Pi2Y686vrpL5RQpCucT6tJHgu/irURvUza9kgNLjLXW32XjU/D9JUHFVIEooxcyI1N48XaHe5cvM
hGTIYQUrp+nhBYTL1ohC+YwyWZH/4am9uc6tZMLNKKBR2aCj+tmTlKVwOlb0MZ5xEYoZ16RAYfzg
yMM8NuHg8OFMRrvfaa8tG0dkac6punlvZxfBrGtKSGsddm7H/VN7rsalewIPrbG1Rm96nJg97xfo
4hhUUaxuY8JYBqqjcMRuZAZTv1K56VIt07KDBijL2X/0DEee7m2Ulfq1WOcuSuD4Y1wcLMsF9iFU
Ixk+r//lqs0YwHtGKMrKSebfELb2ytJMTi6P2RtGEbtqWFC+lK90V3xIqYf/OS6/MABiEbr6yH/z
9dlY1Kp5T7fjlsuXh4aEtPTFSdWw3C7CYx06dav+NcwnMPoVcHrxhUpdYZXDhfN0YQzXpanhkwJ6
e61ILQeTUbQmVw9sni8KpimRd/DlgkQ1/pGn9Ra1bI4Cid/m5aGIL62/jBaECqrM6RJ1uXlaD5SM
JCyWPSVgUpjuskPlzMd125L90JzYjTwBT2pboaChQojtzUITNWYNVvs+1saQuhnd8o1UNOq/CfdF
TbA8gyUgli9Bg+O7UZbnELSGJ6cxlWrMCPi2nYiZ0QO3tG+PQtwi2rIzxSGZyM5/jQkzT4NjJVa4
i60GA12tHgeslsg7OuNsoBlTYjVbgwoU3XNjRPdPaGmBrWoahbGzPWjWuq3JYIHjC5xNknI5oZkE
HDKtASEd+tTDZRZtIR0oqSzbJFaXV7dVdiaixXq5uDLZ/Spj0puPWYYw5swhfGOouFhbnVl+4CLa
xl1UUpq9AmQ5riC+uR6JQSHylcfCw45wHNDZ5HCgNos3FA0mojoFOAIzzlptx0MZDdz1y6NxwXJv
4hpJYZ6GQHYbbgwLHL0uGNIlvMLHFEc/kDOwgG0rNFzkIRfw3uZ3jcKAvZ/8Q8to0KvyXAJF2MOP
g0EwW8GBZ1DEPQlDtNI9TPWctNu2dr36EehhAjDyn5V7CG5J4o4WtqcWiPRoz4vkn1qPrpLsjajV
goZukFUqfEazy/IamaxCLZQih72fjENkGtGfY1LsmXoqTZrI664rM/jOWfGDnnYN1C8TXwx+mk0R
IeqmFCvdR2H1fzM1fTn7VG7NlIZlYRYY1Zb08MMwbuydtC+4iQJLwQ/vH2Ic3z5BYUOrhop85K9R
aZwkodHtPjeifS+x1C7aR+zxtsuRE+tvFI29o4/R+uGjtyIeylWheaAq+uvd/YSvbLO7rNAC9ikz
i6sU2ebu34dsBK6HBNQXKZ3xMSvMNxMw7Y3OisET3t3zeNMIWFV10ubURimRVpOYRXbnMKrgCrdG
GHZEToPF1A8Kk/al9R0/T1/ubswJwWjYBVhjh9ppkd++7+Jec/HITga1TLVhIWdbABiVht1MV9O7
uLsxHEp6dtDdnkMsgkFA8Y8WxhG8lL4guwzlS0YX9ZHHYTJrhG1rRbYQ4bg8fNYQlkUhIzhIRO0H
agSqAy3dkvwwS79l6NFfxOxdrwSb4AllXmAGvTUbA6AKP0XOLD1zw8/SS+9BzxTclnabhO8dlJKK
tZo2CXX7jhOJPmPHhizlMaE0GL/1PG5bd4wIITVODQ8TX953A7L25003Y80UWj7oJYw+xc8+u5cz
k/8h2E7NU3qgsguC+PigVjCVp1PmhguS3QR78wPJrFTeX9Zq0MqDQ/oq2fC1M/U/e+l95vty5lSg
cOgLKsdPpko84zSGydhpFxYvvG2NZ9mQ6F9VJguB2rD9qyJYfQtHAvAHmC1snxPha+DAau/qPXcE
qJjmjTfhznyF78xBrEoXhKNg+r3eIeDXpfpOaLq5cSd+N5WySQnemHg318Q4WyLv/t584O7x07Ni
+RKcEF+rnO+pEpCHYV13/D+YrpaaFRSbsdt4R0DI2oq5oayTrMljml108p00dSIfwsYfBq6ltTGB
aLO8Ox48uQKklxuAOR45ZsP84fUAkxFQtO3k4YUzd3iPUeav/thGSQpSqh/cN+a4KslQEDK3ZU6r
iz76oEQA4+qSemGduCNNB64oArxSCl4lNPPpTJkwOkyruekOWqi5U/cp7DaYL4lKlGi9SEGBQywV
K4DHnmYy+P6FuelxCNKNd/cipgI56S54YFWFo+pjazDhEBDo7rnrsT6FZ0nMpuLM3dVyhFECanix
8/OSg9tmH4Kn5Tp3oA1YwMfFUr4xI6rVbPxSTh0qJtIiq2Hxbvu1PtuLkOgGy8RlZtKxgqhFGooF
sIq15aJA3fT0i0dZG11NoUher2ufF4KBvz+BTkwXOaZ+0hqIgVZDiYRhGLnk9A+ziaICO2tgAYPv
VANAPPuD3fP5yPk4QCyFaWGQTqK/dvLsBYDiohxfzEqVV2qx+HKP3cZTQ8gQGkAESVnbeKbL/s8A
qQWtSRotUl+gUcsXLhmfR12rAZ3y/B1n5Dv+jS3GE244pqQn7kDh12DtAgRvK216knwh8nj1XnkF
v84tg3JidCGv26dyp2qPUiCD44TYc7U8LpryYfyG8fdOUrhXWVeYzBzVjIJEJlVpSKixS7np8WVM
O2t1YfZ03xb91IBsSsWssh2KKBvcMsP6qLQj0yFDEEr9x2yB65vSJNQITu7khsU0eBYR7vleX14S
IN1Dw/tO2y9EZDAX96z90gZ4UQNzpqgGveMlSbFZ0fUb0ep8ofMvxCJG9R2auw43xh845r8U+LD1
a+nTeJzSzrcfh+voug3WWrLBy6iweZUkR+nbY1cEI7SO/9WK9RRNlxNJtKASJEiEfoefClB4UaF4
ByvAYjuI0Ow3ak8izj2wCqrs7Z+BaKr95e9OpHuRIvqOE+rmy3IuTkq7KamGvaNIsswNbPiVs698
/2c/O8Eg0WcwlaVCEYkqjDisB1KxxOCBkt1EZ1x09BMMIPIOq/fA6WXH+J/3Akm1HP9Rtms1T0wV
o2W3XH17mGCloxgs+1KIZ/+V3oFT4LPsgZc9tKbhYBHdYZ1aNEvx8vsFur4WAL2kgFA+0ZHOSKHL
IEjUxUEfpVhndmOE/o1rWGUQ+2Ydq2U3hxOL/uoN5iduuMl0ioYY+18uBuhN5n2ze+7lB+K8UzrW
cpv3GjeypZC20J6c3H6+JTqLSGN75RkQSf3EuMzkTv173FjONVe5g9smSyUGA09mrFdIRKCdZr77
xKJ64c4wZWFe0WaUWRJJ/NtHO+LxOGft9dl7Ct+eGA+1poFlnp/cNEazqHS/zEaN8H7nErDBoroC
FjGq/9k3n5ChPODCT/CNleSZU22IvxsXfY6QAmmmtorOsAwNRIXr5VYvhgkNMyzV9BfInlJKAa6Z
3jaLusMjFZlrW4ViNbBjvmR32Ac/lcVifXSa/tE+WQqbh8mg4PewtVpE8QDyuySAK1RpeaSNtDp3
C7OGG4T/1z40WZg/yy/Gik+BJ8etxa8tGVyyT1Y24ybg0lV2Mn8PAZcvd2UJouO/1fGW3Wf/Ypn0
h8pSCSclQQafjOx9qbA8ind8FME01VDH4HbE3H66eOiZLvFpYrlv3xug+yajge4c/tY1xPO7ynqs
lr5rf8Ny7V+D9pUg+C67kBZh9sSaCbuJ9adNV+axMaENg52SEafLFKu7QtNgK8vcQ4HcikzskqJb
SAKHiBZQwzLdBDYnVASaf4Z0f6Sx6sRY/7acqoXqnu/uYyQt+7oK4e+GaMtWuXMNJ6yAK8PpEpie
aDWtAnj79VuyrGBSB3eYGVM25KE16VtcgOKNNq70w/VBw611vyqHq2SLAvcNV+IDOMwm5uQZJw9u
TaJqt1ESmWhgCQ/UjtmqW/0m7xqLTKtD/mgGhPdIQLx3JtFLgxmVLaWf3s/EfimH+mpJqhllthBV
9r4C4VwHDvdti0HXF4ZlVApNHtugwlwq97hYUWJliHlnb7DEupbNmH1s5rg4OPc7C0rikHQI7oQk
bpUR3t1Cf/izOa/WKTKSSGaKjJyvDEQmtIWXvTM1wbuvz3oNmIrTxMU4BlRDN8926lngA4ckZaZW
zmQnHbTmXTUseIEk48V+rvq4qe0IQSLPDwuxzfQz0gUiAa4MXktspT4g7aygZ0hwm0fkk/GrsyZL
xyTBEdbDEtxyegLS47BcSo+dmQOg5TmfJCmZ30wcsm3IT1EifR1rfJ8kpEU9ybbarz/OVo50OwvL
6ufuIpi0iUUBxjtRzXX+vYxZ7gVQBLggb4ZB/F2ptZPAp0PyScMdbSNXpzFWPj6uysVQswp9qHCq
aUsd+E4hTzuWmaUAQwziQSn8IeNy2RzNyOsFYn8gnAmemxJVPLnV4gTHieBBUsxEJziOhBRk79yq
pBSZr0VZIsYNHdz3k/ZF57PvLFfDiDN1uBIrOJATwyQuDijHY9+xHtYvLdPZhiGIdx4RI+cQIy6V
Q8kvTH7KrTe7PAHlyz82E2OTz7ZOPR6RLobabCWnkNrYrwZ1CHO0j/BXoItl8pReq1eMD20TMR/4
E4+kCjWNtJgbmG9DCOSkpiZvj9ODHztO7AKx4O0ZavrD7KqNwwWUAT3+/5TetNNhfh2Q8R78m+ZQ
QeaPUxxDj4KtLkNDR+03SYIbrPzpeOe6eCFPMbHqtIATRPSeEMt1lbEiOBFUAMh087S6ThFO49ZP
WKlxLfHEgUN4afBbds2qT1uxLKN8SXTXh9jau/lzmiG/UaP8RKncG3woigwHrrhma2ikCZUsvSdo
0HdoiHTYvumd1+TuFvj4kmP2xwY1IQf7CQtZA+Yesopd6SjbHHE16plRmbwsibwPHXKKmCIQFBNR
J3eyzTdSOSs8pqXKGXxOy5/Z6/qbtWzqKxXqHYcSdc3f6Jg2YuMfjROuqVOxh2nKjtFwKGjQ5IO7
QEs61wk9BsxANPKJw7OqLjr00RXFTngyraytTwXAM532nJIl6IKCpru4wWVgNFdv5NQCDw1siq8y
SjfD70pREB/Z0r2PFIhfTF11CinIsVL1LS2kOsBZEh58hb5GwtFfy7bStMyV3EKek2EsZDlc71td
3Jj04PQ+OCVA57AVgr9wvQABL1yGajAobi/yupQN/Q1stOxq3cPKuPwofeUc0bQhwwZiURLcMdVI
SaEmA2E650bNZjOso4oIvAjeyEaKZy/bX7CxhkMvqdXYnfrhge/EBz+cXxs1LbVi28p7GbdcppV5
4pHCQAX/5b78LfTgdXDNojbBScRLC0hWPaQZvEOOGQBrlt89ngSu/xH53u+6cxdVuW+9l36AFHr1
azWQtxeh4UKzjPQOm0hUph2x5/LX5VxlaAzV8HG8yeWq85aThQtqqKCose1BIN451yMg8tKsnWXZ
T9tBZgI9cziKH1dzIe35t3XwizRJLOwQTGKhMrXbSMzoxn5LMeflAX+cmsk08w7n+jkGP6Mg054w
/zyJdAMLHAeUJEn5N5ctQeLONYgABd1+dLoyierbb/05OBVS8PPg4Zj2hH3WAONCzVghuEfR/2S8
Ix4N1vzqbTReAkHFLidt0SLnDi8gKJjzTOPo/y37sLcP5JbSajOHffecOhX62EhWG51uWYEglQSo
rQVhEFFYvhpI/O7DSax8sLGjsAK7A4iUjlREo8WHi0P82s35xM1oMQZ9FrVKIiuDz9epJFdsMC5a
bJwq6p7knGyr171915mM9SfXvCdTgSzTQR6vDtWfUU5Y7R4cdOh2s5lW6FHDJxIj0KvR7hW4I3sm
SOOBvaGOjPAfSqqmB/ONMfGQzSYIU1YTLHiQwuDMMPahVU4ekJYkFHKnHW91xZxao8MDNVyAPxyL
54MiePEm1naaS0rmT/HMSXFPhDWLWLqVYbd4D9fvx4AZPvo/Z0ddZeFCoze6pF64KUMObH//3FmS
e4xokQuTivlTARSdPPyDqesM6FffRoc3D6O6Ck/v247J+9n2ha2B1J/REZ1H+KEQDTqDqxO2c5Ds
cwKfuz8rgLUHKj1LF6m8k55txL5E0TnhrGt1sK64vzEOLQ/MbtiFnp5TL0huP3C46cYVlHJ+szxI
eWmkYPTqmzIOxdwZretMOvNH6PVAi5XN03DCutdYYyD2Ge0yr1xC/bXkXZp61wsjB3ClMRjAVsWe
3DJF7UMuW+b560jQ6C1ZYpyRdA2RgZLh5O0Vzt6r5vsH/3fLfudb81iwoSxZRLj+0Efv9sZkpav7
zodZPPsqd12w0qn8AiCYm8XRXjhsulYgvapb2sDpph9LnfCZpgtjBTHDXdlyUpnrRJEIz0LZMuow
psKSm3R91zIwajrJcb7GCX2kLphMn8CWBYfjXa3oUzx9uoU1bH54wkcn5E2BaomBnWWGbxeFlByz
VPhcppNQx+mJPZHNOoSWsfcI8P3jPtIWW/qrsGIlAUmFYLoRXW48NWk+IN0xCT/gHW8V11ZFeUFE
jD8yY5JZW7sf3vnQ8GXQuGICzN775CnvKhFuGuBe4rtSjUCvTeowi/XhAqANsHjLEdc8Ey5X30Hm
ghawu/qh7YH8Y2F6ZWMm8hjEyZJv5h9aS1e9kaJc9H8uqQPDgIXLm7O+XyvBoXTFsfn2C5p6b8hw
okT+YYO8YDrRWmSaDgVpjbZXUPhWt/xI5S2jlDaUFtEPbbJb+4UJyB4NpDCrrBjPgZUJ/9WfGakq
Q3pZXSlBhygyVpGDHZiztFuAaqJSaRiY2Wxyf6ISDsA3zNJgi9yxiZ19gy+v0EGRtZIGi/cpVARD
ovZY1i7oeOIGQ4ENDEBIlC3rspQ6lQFIQErFoEQcMXKxWVTHdJR/MM1XdkdLarA/GTflOsdpdY/B
JI6pNZAxUkjmjQnzaRwedCxgm3QPh14T7kC1Cs0YKcmooSb3BW1cgTOOfuCvzepYKSDzDjr2027G
G1ldCVr3FUqnn7clfv9Fj9zRuNx/g0qW+FJOAronXLdDsyYwG2tERUvsBqwy+p7980KBrBN8Aoey
4PbffyBZp+19WXM0pbJW7lhjvGfwU0rUsThYeerMFVf0TeA+bGMwY1qfWT6Xj5wuDJk3g5/RVFvJ
yhQQ0MYpTZCwJoAJWkes2oUiv6YNp3F7jjEMyvdtRR0gzjQFFwCeYBaIVe5E6ZR2VrUOLGXbHU9D
EQyA6JaR1F1bk+G/C7n2/bOUZayzt4lwJCNnTxleso9jOtm6kb4Ye0C3u3mONN6onUpSS5cpcW3c
neHOiG4F3ttMhFP5tiGLxZDygsX8oTcigkTNxGbCE8rNMJwaPf66TCnzW4Skhv0A5GqutCpANkbG
kN/2Y46jBbDPLnStPUZPg7icqwMQ6QKFYVZdQddSkRYIxHqBe+yWvZDIz5jUAGmcD2wW7Wn4OZtu
6v7e15EybUHERo2DE+Q3qe1GbkquB3VtEnpILOUSeaaATQ7te+8buuv5PCduvH/2gqmsOG3aJ0re
UwwdRaeUE+ZHsMKxVnKlOPnyvlgSwwa+onGCCWCox/JVuNQyALyAckMtXmL/ZC+nB1wdJMYprIOE
nVBoXSJd/KHHClCg/5w95jTV08WJX85OS/ZEpbei9lzvMK8FDruOJBSjl1k321wkAZ3Dmvfpw+xS
83KKMkavlFI338MdcznqQ7n/fVAAjHLYdsgwoVJD9BPAQbLdBn8RyNmqFz5JiGlQ29r+fBWYk1Pa
AQxisEAVlHchOnoiPCu8JZd2AdJzrCAhlK6cifs5WMcv9/XvK32/0WPqmB6/8t+jLU9Zw6k85Eeo
hBikNxTpSAgTRT/7V7Dwd9lPA5pVq7xf2DF9Plg1BJ5jBt6thBOmc6x4w2zHXk2OLMGCm3rRu73M
wbkx0BjlIc4P7CwviIS9/45WfVQs0/bidFjfsIi9bDbJvWWzdsDl4dXfpQcylGcHVP53I2U3Ra7u
Z4jyR34xDjFzO4szPFWrr6HEhUVcnvTHh/fxRNDo+4VOiVRhuAhkOh1nJt3SQlYyzV+2iLAcAYwF
DvmBQOpR4fQzBfPmERO6+Z3OQyYN85OYrKqZa7p1TqDp0Iv66rFjAxMkwowPNYw+2wNXFCavmuk6
Frzax6RuUltNrby43TQHqGLAnqL26S95JNWmhbAxuMuFL9mrpnvqxlciBqP5Dv9LjOpGwodx+Tmd
AiC7gskUUV94tC2C6zXMbpqbJvN5B6omzyFaFNAq2xCktEnskstph+luGjUUWOpvglcOEni5JpDg
T4zDQpDYhLRJqbVMaLcbQc/DIO1Lpjq+vjXN6MJ19Hqx+NbY/d4nqeXlXkwUBrDdTqg7qLc6ZrF6
K2SVg+0QsLh+FycTVicDenN8Ivr1a2EHvrbHKUvhm2LOpbgl4nljA3JSpXcoweMBSMWAnURP6Ves
WhanlAMHLbkxTmIByp87n5wAmm5r1FjWCu5sObSa/AgQPT5TW/Ij8j+Qbc0dhuu3ev2EW3XOvgy1
89OB5spxYCEh8f/8JiPkQgbKuALdFVe3w7trlOM5m9dRRU8WN7u83wfEC5ueydXvTnAqVwqZDkod
W86qmSfLUlQVUJHWUbxj0XdNjemwIT+xCge9r3RnP7rsUOMiPkQnb8Z2i2ZVr7PHfNYXaU+eCRib
kOphTelUdNfs1vy3znDJvr7u9Jqvx5CVPB3jAt6WC9Nu+JXrdW0hEuHL2dqJAP/ujqkd2AQoHZh9
UAZC8CSndxhbGIWikhlaBuUxYdCttnj9PSHf52fQ44UGKQYs2nUcG4rYHwrgQ8AttNQxByUWh4Kh
VcptPkPeQWMltWjgmcQSBNm6qc654kTApK7g/JYfexXlPQBtnOkxdi36oWrmVqYri5ucezOmAGtA
w8OQyfcP+hRYObH7qn7D/1FZvfCU2VTeabeG1Aqt4ECxfF8LscQZMOmihe69zg559y3EDXhOqIKJ
Zt2rJhgwUtV/aqYtLUHYaukZF/nMyn058JOHKS6t083oKeE2ZkYM0V9zLThUE8KJnvzLQo+TMbwt
V6SgFBMmBSFrfyeoI6o2sfTzDdXBQkktAEV+B5vyKWFK0bLoFWGAjOMJAzNnmU9KEUSlhJP/mIKI
IfqA3jhgW64Jek/EITLTE9ZWh+yPXl2/knddJi19CLgKfdbl87uWd8sN0gyZ0F/VkcO7Dieps5QS
N0/B3tWuRfhRbpLJDKCTbfb9GZUE4IXjQbngB4VgjIq1FhIE6LPsm2lZcoww0NeSzHPHgz7klskQ
1yS+65akeGbqmJD7m8TIVO0YESCgJ4a//cs11ZpOPyHIPmNRS69QrPEwGlGrzUNi7cjIvNZDdgkP
uXL2iCjnYlSKEBMb8GyamKGl6gvkwP3HeHdCe7L/yupJcFmlNyKOgjguT8ZJUgQHoH1fRJHietAa
UBgkXRx0AYV4Iua6NZP/iVZPFLSM1Lrh1xbia5qWh0Hdjys67zHQrcD7sayRxeS6Nu4IwMZG6L4B
SJBljfOxDvVIV3eP/ybnIsVa4qo0qrMiN57xhkfhrnkaLO/VobGkz4L9yudvdPoJyAgnS5o2VvUq
iVDUJeDsLatSRDPGIF9+/tjslc9YDZ+ELXO3xdd8OQINmbMqchYhK4YzvS3zYZg+JP5LERRvG0sp
HaN94PSdjqlDsQOwaB0nQe8IELt6tuTE+LUZM407RRi9XdD8EChZa0YcaZ2FMV2rIJHoBTjbn0B4
zNUfSmLQLhyl5UREPn/S2r0Gd23KffIGWfDCC9a/jmpCwuhqnzJFLFi14zu4jPc9CqNZCjkDTYeq
qff6bqnJ3BmpSZFu0Y2o4WvI+1ItqLVmj2SeKJbstjyRHu8HYaRBn1TT3RzxM46WlxBFIFjc2KRI
xQDCpwa5tx3+RgYmh1zHIKSOOZm0VpxNl4mUDnllY3wK3GpBFQkzNBBvfzrBqeXhf6QBoxso41p9
624OnUvGGuamTaLoL1M3m2N0dRUqS2zEE7jvTnk+RLqtw/MCPA0qVUKor3PXw+lqAAI2ZLpykDQp
/8H+cmQUTW0x0zlL/5vYhMIf/uCIUQg5kVOE+EmVm7FYi8uE0r4crcT3bFRDSwdsX5V7knY+fzsS
rVAagyWzg7tc6c6PPOuTf0bWhShx5WYP7UburgMUBELfupInhZD3TBGnSHzFcr0glry5+bj0lAzA
qdy8LGihAgqrIaA1jtPXM33hRtqiH9qexFckJUrWlM3DWh/mVsNS442x9uv8lhnmqfpe3b6+lDq/
sqp5R7hz+pRKziEZcRVPeVqg14I7Z1UYsnkS3xzrsLLPsO8b9w5ZDyr+cyOYLWcNwpkUEedc+okD
eW3ryAtlm0Cj3I6+gm5aP2OK6i0LObBGjETG1x2mrWNgLL0OkCZiNV/Z8UIetKU/rFme3jLIxmRI
ez9kKgcolgZeEJ93JbYr+V9BQdPgsUxXYjmVdLbvfdUSomFPS7xMjIvi5kk3RWk/6CQZhTbUQ9U7
ZDNlK1gXYUPt1srUTaMXmsg+iRklyqFAf/03k20pFoRu4xoqlemBZFPdHreMl1UIP0jEtnyVxlWI
kkiOdihdFS/esc7HOmXxXs0wqFKqk7IU1DQbgqJKtlfc+eg9Z6MtIKqoluQi7p2A26sGCVqehpAt
5J1CNoVIUA5a+ulE3UFp+cl8i01KpfY01HBMNpRF4qFXVDt4TfVW+wgknEWqC5iHB675hHnmrOgN
wGsjSe7q5ZnRxy9IkBRbUgQGzSk2/K59/bb9i+AoIoEGimaik0f/cGIEN6H+eTeXDiK6TUhJ+CAH
k389TDYiPKs2pkXUKi4fksNKkFbACboQV24Jam47mseZYKnzntHuMjHihWfeDE5iJiNEu4sbetsc
OVnw1+wEjYmjtQllVjuwl9PkeOSK7vt3L+2ze1aqoBh7fNWRoAGUHjtNVA+aL80SffHIw9kujBsN
dQcz6+3pL+eqfy5JFUkxzw5b7hqABzI5KoNkP5G8yJnSnrj5O55nydb05g5untpROh0D3oxWAtzn
sNJXQaS1FgAZj77+sbzQv9ixUvh2baTFBLYmW2Vxa9LlZq0+mg6vG5P37q2DjO7PY0LZguyVc/YL
3AXfoTcJyNqHi+8bn7+CisMvr2GshymOyu7sjIONAaR3r6n99RiLHmUV6N8ZuSYW7dGSPW0pD2ag
GmcA8GtH4ihcQbtCtafxu6VYqUPnUXWvyl6+dGpzE1FxoEy34L8Ro9xVaOxTOtofljN7R8GzJ/Cg
Me54kzwf1ldBC2FBKPJQor439RKcTtdJkehY2Yepq0MbMPHIQ7vST1Pl3BueitwISQI802WNthSV
4wtriWFWlx/VEIlVWvtTRfCWgcHtYSTbDaPqAf35040ji/K20dY6C00A1Jmw2KyN9+g1RiioWpDH
r+WynCC15RAKd5NwbNL74wlSyhT6cyqqgENXR3U0se3YuWsia1WIMj1pfkh0zUKIUWzBRMCmnUPG
Np1HwdiraLTzGz9AupAUPwdXivhaOElzqCPJWElKqHQkRZj2c113JYFicyr2qT0/Mow9A9F5LfbU
IkEIyerl5L7605InEcPQE3ldxWG5ueogdsBQKNmbcDCWK8NZKH1Im1JwENs4g78fRbXBI04UVdS9
+5wHh72enXAsy0ACvh71KT82K++bUFqbJ/9wUi3XhryDv2+D3IfLE6JnhAltovSoG6Dg0IcClaw7
uDBGGxseRt+yEH2dotg5wFj1U3WI6FL7gKEwEIu7fyf2y2WZ8Ki4ifLG8K5qNUprrboXFwFMBrPK
IIWZlBPe6yugoFL8Gluh6mKcP9XzrqDWjFFuVsA+fpgXO93zjRjd40VSJGDXgC3nh3vqRgZ8SrUk
GYymLVltJGi2jqnIFCSxjrwkLFy8lC2cl5I8b5bfvwWsRnJrIGwoApNDtGpb1bC3RtLrB98eDyAp
vaIEZKZccvbv4Mppbc2NUm9UvWjoFSy4gMgmBwkbXgRAjkXQMpig2Xw/ehqNFYAanKrptbNmwIUI
UXmdQqzkw5QFkRaqc2PLF1FB+kRaGLhlEsxs2okjNNxAXerGUkfKT6rLkzKA8WMXj0lbM0n2CCuq
jQlIVh8nFfCKd2+nZeW6h5yQ8awao223q8e2J+MMmkWvmvGSWEGEFRbsUvzFGWU6wSE1PxWVHIQ8
wxh9E12bd/b3BNJ2t/u6huhjCR6MVJjo94tntkyAGSb0/67kcDpqnMgCXJKKDTOPb93OeOkp61Nk
I4s4v7mPHLlfBYZY8K2TuMbxjeP4nkINAzAj9VngTfwVIaiLmFuE9cfQ3LSBmwho2xiQWZ27scQL
znr7j9V5wE5s6I1T/ESqicPceUvHiUSypWQi6TmKeMfWlIj0zhGIh9kbiwgv9T8rPJRnnmw2L+yg
/4R4kmFdvXhXjUCk3pSPq4cPidt9nP5v96Prtx1RznJqMHlARCWMhUy9dBQLRflE7UAL5MQB7LvP
RxBF99Q/ak5ACa6Se+tF8Lw019Oc1yp4kUF6MbwWsMNFersMevke2I9RM90V21CB45rnEbQZEHh0
seF4mxUWvUFJL5maLpCH/Zs6rzzsBoM0kGvLQefiNEHb1jMgfK2GU0lSxq6x/S/JponE2/FlJdno
6/1/0qbjKsFo3WgEbXi6zL8D4jMdzPUCa8HkBPdpbdtoSsMKxCpymv1jeLE4GqQd71SNigtGi691
W9q7Xwbl7ehTiSBL1g6SNW+5v+gu1bRoctiBJa6BbUSER021lo64jzbszMWlRZdFr1sqbUtaMHtA
VeWvLMaCctjSrIZw62mZRE9DIthZT4N751cX3SkNo6IaNp9bLh54grZSexNrZqOCmFsujea18XeG
TeXM3NrwbE7UWiaOP+4yLR+ixrFgmbvKGe5U/bqRKkups+ML4A895hmiUAtftS///fRs9w+hhdwa
qUn1RyaHqrwoP8dbINUnxPQth7otu2VTu743Q2yi1rm2oZSMw6VNBMKAjuw+VjqVs9j1IxZDXnTA
dyXg/goDgIV5VuYL3eB4A1YY1H4F3ZlKjxe6KZ0ow+cuMUp9/9ccGsl9W29wn+wIiChyUb/qKypZ
/f4hEeUCcfjtX4XqrAARYerrklOx55V4aSIyq+nlK/fCy9lmnQ3lIA3uUX2VWJbVfU8ANY0VQgMu
YO697CqyjaI4XIaMuYYGMjBKYJ7jZc8SljCdvmD6yKOjCbJmsIBAoymBQ8DCbzVeIxS3pex8u92/
1+IQJd632jTXlIOi+nY/Tid4elWuUrk+j8MbtsFUIqRSUMd3oV/9MWGLVkiWyNejRI33VGJ2zqM1
enAcjvxfr+LbDaQ1zi0KNbeqQase2Q39ybjkiyEGiHoYzw3OvTU1YT9jpz5ijAlGioR8JI3+Uzja
e6kYFpb372srAqMUKN05Dagxq8rNPo59kaYjVgniePaynBaazBFkgwRQnP3dIDWj6vcK7leRqg4O
iTzQm0JNLjatP5KmpN9Mremy5BBESoua+abRwLgxwBvVE5sDnKvFhmhIxeWj6qxzsyzyt9y2ILFm
gqLt4C0lTqPWJvpq5n033Vctjhzp2gyblBIoY/eLYxpeCpOskxwqXQ2BbwIzJWIZEZGgL7H3trlT
PY+tfwjCGuPvetFwa8dOxTkj/koO2PM4MFip8aDR5ZKFP6oews8GUNBTvDCNLPbcshpO/72p6k1f
JLF8DaeAOcD2nrdoZmGkMUm+oSKLwvI+Hs8MjrWxzE+iRuudCIVG3acUGVZPMSPclZuaxm2vSdjZ
mY8RtEwq69Vb1dsjx8DA/WcqlnayPb3/65I/frtCZaOp5rVND2NIz24mgrVcqVxfFddUkjH6MKER
v/YY3Iy4SDyTW9JH6LSQSc6xO4s/jW+uifQYuA4QUE8pKIFsWx5QQ2/Gz7SyPs9Ot9RUI/kj2/Yi
BQ1K2zxkz1YfIT/4d4MjSw9s/xjdygkLS88LWGPps1VxRy5aZf0SW3MsoK1qH2kgt4RKPT66LRwl
SbcrSjMsJoyQsK1bK2QdRB5ffppGhGeQNQM1TfoKVZCfF1ERqdoV+zrNuvCaeUNiRg3OteOHbttO
XON0X1TV7LMEAkM1vBJR+BMF/4yBVcPOZ0NqDgLWIqJwNLZXGRQARCp0Sh33jp6qZI5YCQ7WeRHF
m48f7YJj3x38gGy9wT19mkKWi5dlD3onsCmlv+QvdSG6o/7ebuSa77B/L06ZU4AfBQuVeL29/Gzy
vYuu8ZgWt9FpKohNgvDff6f9+mFyJLX8SnBT6PaFAVAUd4KPDARxkHGldOeiERmQ5/BrLpz1txho
FYNFqhuYew4sX8/XB/u/eOrUvRH8DUkacithfDa5W/4rVuvA4cm4pYqcdBId86Gf2r7HPOqjP367
OCLBizLGmajR2wNedE10wQE8GovcguegICLVfxwP4ElRXt/jmf8q320BFKN2JkhlHYYVmqDWvm5X
+mujmD7LycEr1dwYnBS8gZJx7GWePhbsVDU/HdwGfOOt46z3J3DeRPTXwm5QaSJHMhhY2kYSxosd
eJ5pnF1OKOsZ/jje2EyKi3/2C4SP9+7PaCc6NYW6aWvLhMbEjAoI/maHerkOUfMIEd/EqJClcwoM
AAXE+Vfn2z8PyZCbKrtmKdgO8phnZJhhgxhHKK8b4GfghyrcOydpNL2aBCwayfqtbJkn9aoTzMEt
yyffdjFg84yyKBVgZT3f0/yVXr1CUpXxZx2hpk3yBMHzC4BUabUWUwTZ2Xj/y1YrkGmNJeoKVjLp
4CHaHDz3A5F4iuvylhK2c433o8MNRhdGZoxZzPaIjbwoib2eqAkw8oIAjM8oMdf3cn4XsHv/fFBz
xvLTJIaYhYM7gtrKxzA0i6k/czO33MIG/L0qM5HyMNte5Dn7L7rYp+066+oA4zrOzQ/tMo5D3GFr
DP9TdBXFpu6FOFGntS8waRqQd5EvuIGlm+7zPJO/Tc4XenieeDOX+bXfy+0CVaB840Iz/3N6R12y
IvyaFCghqwXNB4c1NOuMgySyW4OO4f4MBVT9om52Ohtlpkp3q3hdZuwer760xPXIgxTfUaGOLxDP
dP+sslsSWIfyyzJp8ZwTA3TC92FePs8BW4xqY3u3eb6DLAXosc85CIQHZ/uXb0RUsULS5e9Lp9VX
t5tTtgCrALE7ERm9Sq+ggcsQdqH8DCrJOzevIHgMXNbROFTqAfwFjSMqlY5F0jGXX18uEMoDdTxd
1L4X0WGHyiR/xEl861Abw4TBxhfZqV6+sZK892f4dM8eDHwvYkRoozH3iHpPT6dbK1YkHe2HHNuw
G3FNbZqEXa5C5nazbJP3n5FOM4VlLZ0zKgHXIf/VSiF/2BqqF6vN9fro4VwfSxLbySeM+G9Wzd1U
E5ikRJ209A5BrCYZU8aNSKoPCxIXr6EjrCHD190WB/U3n6B1TUmWDPzPdFBER2idDhAFkqJOUPeK
Ije6TzJgFQGY548UBK4RlfSLOiRtjQkysVAaGXvC2M4WGZyFj5bZEGwBNXaTk8l5Foam343KgRzV
+jfj+B335QT/kSrINfjDd4mnN27trIrNCpWz0niBgWI3rBDVsTfF3apqUdyInDV21RnbgdZ1HYhY
TGaypl0KQYilZMvcsUM1jKPbjlvZDED/TFjPuO3uFClTyun2mtyABHnxqDki+3r/x3kgk4zIm1EY
9AfLGjKEGcxRu5zO7o4EuMhdrBwcfifoWUOcDsbA9+pmHGSZYUHkABivLAZCRxC8rF+8rxU5qKiv
f70Jt8RK7Kl4/fVFZfnfZAjih8i7wFDwIPuukJK50d3/MtdubuVFOxPiOiQvTL16L8XcrR3Tv5s/
+V0J3XRJPELcXYG1DZVJzT2S1fkUCZ99lSD9YXzkyPXq+6vHIEQ4VFD9zQcPHuRKFjxoNZsXAlz8
Jk++6V+/eV3omeWPzdwBcc+BiaHdvF4MpqxFp4wMFozJZRWCqh5g9M6UFpUqz2oNyJ/Ky7M9ur73
E/HC4FgA89X+NmOGdVjHJ71uURLI/0DrMUXtoM/imhUlHEs1giZCH9yrGFVzmrd/0tpTdVz0602V
X8RcEvEqQS4bwnnx3ioQqUjjfhr02g1FolcBDYWMODQQZHZUk9XEe8J9uFgidMOga3KluH18WTzL
f4MjIv/166mjrAN4+kDqj84/c8Msj1+ClQeyjDs+Ss1jr2egjbMUOvSQ2y7/tZTpJ9AfTlPDqJKD
CpGhrlPHEt7b1mpoHS+5Ef/7HFCww7GOz9v8jakGUykduQ6QGo4SF5Xrk8DmsVnzRWMCtaWpOcA/
XBXa4xhpG9tVHXV72bmCJFrmjN/C4KbUozfMc3DasVh9Gkx41M0/ag2xU25M1eIkcGqnYtau278S
RAPwUTbmPfbKnShvz5DnZWI6RxUCmmB1Aj747HwN+kHgsT4nGYzci3yAf9zqTVftPYf2JMFVAd5j
klhhzXUzV1i5brPz86H/ctRP1Ne2HD1WvcNl30j2gmRrEAQ64B5hLFjUvnLKTiWLV+ZyXUAD0oK/
RCPzi3mP+XhgYMvTVAXmmNRbzKliiqIAdiAM29/YzqmGK38I2S0eRYERxEwo75mEmi5TGOq1k6Sw
oAg2RKAtWPs0+xLxwQ7fGeTEu1/q9Yvn8/2rSEuhIGpR8es+pFHnAjzDwrosxH0n5ZYdH9kXUfPd
pWU+ymPoq3ur4TptVDIoZmveWcsS3xdyZT9YoYRT9GXLFc5rR604poxJPBx2s26YDIdxSL2DZCYk
zL0uSYD6L+Qk+cBqczPmLxC6Z2Cl8KM1bEFFDCugOX/W9nU8ojh90ZMSTtWUlnes/rGORkoLp+jt
/JrCzXfOMo/AV0F3qZ+dJ73MLe2WgyHBudknjljWZhOTlfoFFUXojZ++F3ka2vj8dtb+DLUHrHNC
RJ97u0uBR/5J7iQuoskD4GqilS6VNR31ZRA5zhUbARn+ZJkN02vp5d9SkhQPSLlUQD3dbqQ+cLzD
2F1Rnx1jLa/eV0yduzxtZwwsaAlAhlyFWGh9OHSERWT5H+Tw0Rxh8DCfI1kRbLzDDgioSTyar3JI
vmbB+RmD2GVM60cH+n3Rr/3fgqTXKN8m//Bf4Mg15PxV5YIJxAu9An9MNN5Fzp9Wi9AnRnTPHXO0
lLunOalUvcsR5hyg+nu+8r5y0ko9gsOz8B0x9gMqb5e2lSGAyR/aR8s/LkEXTLox7BDdf3tEmRMF
E3bkXtkjsTOT2G6OEh01TdoEK1Z5ZNjKN4SsV4WhQxb+yv2aF9UrwZUWo7a4QXmUtOQVYQ9vHF8O
UCiu6ctCaaMAKSyfRc9xLOnLWnR/VK8rjl0jTeHnj8Av0AD7pQa3Rv0s8R94TvL/8d2/iluWC1sw
SZ2qO1aP3mxt/Fys/h60t/2Kn0L/VtJgLOweK5jt+MiDJp5RJ/sAejC/Lbwm2VsAbO7cnXxTGYZ2
XUNpYhpOjviLjqybDuOEK8KGV+9h/fD0btFZdB/+/y6Z6IsZF2gYTNb8pB830qNWCJEx10JJc7Ms
5o+g2gcMKpGVeOCJziQxdjLlhz9YgMs+kANckDxZa8EGazpCqMx/Ivm0feR+t6UibCQiA5QBms5j
ruGGUyM84S1UfiJblUo+PDG8d9FXRYHDWtHyJsrVLhtp1X1A1N9sSjgXwQJe8UayGQ3zPZIZ9En/
3h2AjL37XYrjC11NiNGabMDd9zDwg3fx4k5kBGJhwpjSGW8iyv4VFH+AZZO+rl6zGYoAEUkJK5Qh
ce3hoFSo23/9nxpEC1HVX/mjlsEqa9FGxDbG0tntSf9X0ljm+zChSEcy3scmRg5Mp424CPotz7Ey
9qFuzoA4iIMqlBZBCABlMEXyKNB+rYz2eCQLMYoiERCgGNaTP1o3XfQmkb60tj5ufA7iEr9lbzNI
PlYQy97FBMwY1WJ3FHSzvpJTUaNGQPnz5kn6ZgyTbkgj2SsKnl3KG0R4UH0raOZ/PGqgHN8EUQ6c
2lKk/8Bj+XBwOX91JSHvXjTKXx3dZgBO77+MJ5RX7aY1Poy8ddOoHQ5dwu09bnO6Yz0XGYV7FvBx
31Nitxto4wt5nv0y+D8y9wakK0itjD7nRAs23hVEpHnV7Z+B2tMg3GnBubD9AR8GbydogsR/Xpai
oUkyLPZnn9RQ0DgozQnJrGlkYAwQZR2cP8YVqKXRfd5bQP6I02qMmYOAUQ1cp2CthZdk1GeJChIf
MvNGknCkgMBs9bFS1kI2M0V+w2IthRSSQ0pBvYEz6dlYyPvgLWbQrws1T5oi/gxSnkKNDC+qw4bM
Ycp9xh30LmIdwkeA2YQynVCGXK+Deaw7t9qLMqnXUC2C7MY0gUXoTKIni7uO7zmr31E4AUozW7tq
O1UMm4k25c++iqEGE+/rdfsDvKmT7XpBsp+QCOK88nMDBDwvQAkCNKoIPHUmsl/iYDR+jS3f4WhB
Ks0JSNV8r2uHt3CWQZUcypA+AqIM/r/y5bVaisCALczEFcrpgi++dWzIJs3XFswnGYwFnThcWPnT
K14D0Yqq3FRqh13+acKWSlng6D1NrXElTQmIGatM5AeBFrGE6eODxwIeTVMGRI7tKgxKqia8FbM8
vr/75qKAQVdcCcbRFV7vLXwZQZqDs9h1z6FHFNUjfiEZyC3VaGWPYC+Y/P69Or13q/Vc3ON+d+3g
roZ6k2sON76BSEZP13OmgXw7uFuQNJyXNmM6qX3Z8wPqFVSTScBCrrHnOk3BzHksdISauIhvbRLW
2DoOrCJHRkVJ0tjKmZlKnAJct9bmbOIWegmStqstLb0XTxv5MiNywD6iKE6YjS7xr8u6FEG9N5dJ
SbYpmifsVX0X0QzvZsH75s/GS5l7yVajwOSKYrpp8oN4ZXrOLylcOXU4AM4r+ZVIbD+KxVEQkAVT
KY3e4M5Rsc+YjM/YYlNZQjV7Sd3iwgY6no9DKXJqGVh1bFs3WXWU9P7UnMt3UgLSBut67vmLXZtZ
kIkl+1Mh62T3AqUI5mW/IfQTAZkI0PmQdQE9NhnjYw8iQgv5ATHy9DGL7kTveDeFRCOlSIIQl0aY
VKpqfPXoyP08cmNYZaTo71xk6/qwQUQ1hO7H3C2qtBnrWhBjNeSpdPLPBGlIlisELg1YFRiwLVG5
QZB0hRiHKDx3l0KXCqCiYsvaQbh8eBeB2HjIwHxO9Xv14AE2XmDGzFuG2vJEwAgK/NkHAzMrQfXv
MP9wXTP3PTrYS8WZFRB7Sl6aiu6L0D5oBaEaXLUWrm7Wow7rYsYfkz0Yk4ADRYoJc9ih9+AxP2Us
Clr88g4JdWtDeUdLucMnefbxeCr6DrGUrQyzdTn6rB158T3zTRLRVMUVfl6mnSyBC3A/jio37jup
9EpVhjrkIZhIabxg1cWIMTJqDBvNE32Ru9eOfMn6XnHXF4BRe32xkdGXlKLnV8YVbB+rrj4BJ+CQ
K+MujwQ3P3UJ79q1XTxnkoLxEx7erG0czsi2xgpGLXDltxu9rTCku9A/UXDvBJ9M35WPFo5Wl2CP
jUXrldbUthxYrRM7+WxJolYh9WLx5+2MRciVeCa+evSf69KPezwup4gsTaC8MH4iq2XOLE5qS7ZK
ebZoRCTyd62V8SwYGUOJAn+e9d84jr6EPiwW00KZ6MqMNAdvJOWWii0k1ynZykfFMnpqNLW72y/9
0hIiJqAo8uduxwMRICf2XtWlqeIxCCYgFnYV2t23YFVJUm8AYmOfN8Ynih2mOx/693hOAlnkCrNG
+RZjlMpoFDYIEVQSeCJpT2JstrzMFYeovnCIXS5WIJVvP6eRJmxFqZyQN5zsZRTEcBBKn8cvj6ST
j05u7eAS05CJZnKspgetA8ad4Quo6+TZ8WgcPtwrUXKsr1HNWxvQglP0XxD0vmI1iNhgGi/muwVt
EfEjVT1Qh62LHrC13frE0ZirQVeHBj1K2WgYMejZQ75G8Ooe8YSpgM/mu+7TVp9CSB9ajdbGpCJE
gt9rDUTnKFPmGazvbk5UV9sBsdQf5vIWkFSX8ufQuCTw7vthKBq6pClZZoMZFMoQjcMkpHwry56t
X7mKSeIve6MVxvfyxmirOC/ZP2xGNCmSGUMmfzmL39bs2zUqdinWfRJ4S9KuRhtMsTaHtBDNmnLo
TYdqA431P4ysyRjgKN6Zly99xGRtIXw3wZBZur2rF9+PTnhu/IYWegu5TYQ8a7jZvESI7efX1kFs
zovlnnWiMmn+6Tz2wK5N4jeM2IHTyfGfxz1/oqygVqK/AvP6MuIxdw2z+j41HocDxsyj3XyAf/aH
ZeYeKiwsKb81VDW1LWO/NedealHZ8NvBLLDjxst0HznPtB3MaZ7Gi6vmE9vsIanSMYyRMSH7IW5H
S0ITHZYfiLrUyIPaFeaZa6SOueiGVGy97Fh8WMJaCxs+OKyq7vg3ZaUTUkt9gzQgCZQmO6EpuPTk
tuonwvtKNZlDWpSTlB+y5OVUjjsHHTWeYt8BBKDBXqEQ4tQkVbZQ6+NMYXUOZJl02SXaij04IYLe
46odq7wC3N6JC003ol88Te3ng01PHJ3e7HYbStiSYONPTcCYqRhspT+LZvPXj4esqOjH4KfXfGJ/
mBczq55HJ/9h+hTuJhmM+qoEp2K7pSTHxN8w0qLbjNySQLphxtROU+hohq1TgYcojSm5Az0GLjDE
lv3NaXMt+nhT78sTX/epEzJIdSyAjFZq0coACAGW5Z6TMvpzEvJCmxIE3K5uV29EJiEvDt1iGsLi
+XXUTPNoO2wEYHvoWBgdo5UKh61qI1uaLAAvwl8IrfrY3q5oojNHm7B/fqhcs+dhTME81hPUNUTv
U7TbIpPI1ZME0NhTIFderEf+THYBwKt7HGc3AnH+XZop/G5j+9dK3aIWK3VdT/C2i/Ho4wIehOVW
9Nv15gZig952fuF8/vd2Nzxi1adS4RhlyC8O5+dD/MBh7bDFGAIsSCVLz1DotkpwxNlVraLXnFdB
kCmwWc/rkVd/ka9Z5QZm1uJlCCQwjMl+DHp0/6l0PU/uLs54/jFYEdmH0TTDoEsDJ0mRn0OhNh4y
T72ovlw0HNOq1bd8EfDT6WTKLU6r9tP9EF3WS8YYcE3XC8LwxF+z4XWBA0bwa2ujpeJzEF+0Dkko
k+KHDeYzccR/c5/wk1kcO7if/UQopIeCdA3cHI3ZfGQ6ZWp8HCyRUrvqxLlmZDeLy8aPYpT6goAJ
Sli09MV3tArlaO0rcrq9Bd4AO/LpzmtBROKXsnpwmJ8Ijs0QIPpOjD0lFxj9AT8qxg1HFdZfNJS8
jcv7XE+C/R+RZqro73a1pXudhNvicGFTWWVhMU4Mk9mgjY3/XredSsRy2RDiTTDYw47VJhDudSSx
v840Z9ZD5JNs11KZRIMoMXeuEK8tzOCdKmPsye12qmXIB+E9LxOTpyeASBGL5vKlw1DBbm0zuiHT
X8bmslXtBuWhR3k8XsmhV2sP5Ile9mqR7mK3l0mblTWTsbHtPLLRG2Wnc/8qM50v64xwwe/7lQ6O
7rG7+NqUxt5tqth3NuAOxzbI5wDAZ43I4zfqYKaBGy0EunymJihk15ihwVYQqTScyVehD+PcUfVI
m0xpKhe2cdyvJxhwL3s3by+e4JVdMnbJUY266yilGUD/41fl8MnTkHtEputNqITrrH1UDUVdr3mI
AqgGrOHGIWCA3QHGFwTK6GIwVLqfKJp805B8Elm/dVlgtVV5sUQKvWKequjvY54AH/wqMTW+Flf5
iE8zsan9YPzmNov2nTjkEEZEuQE2e4Gj+qXrMog6g23DGPLGTHlu5B8jKelCir9C5LKdQspFoeTy
PuJHoqFJ/3YxnOmnHNGN2FnbQl1PzXnjjcjKF6DROVJ1qXnBt1We/JXK2LzpfJy7KYRXWJLlzaV9
Uue+NOpZk6cKnzAPAcLsiI88BpGYzmb2TjD3orKF7dM7xH10/hqthyamB8t386MiTGtohFWmpw1g
bTxNMZWCqTOa3hG9al5ALrhZxG4zieWxIx7yRLrdrTPFLpr9f8DRiVpaj6jr1d21J58RSgenILQD
truFbgkufetYQBWFVsV+OMR/HJe1sLqh6J+3QQDozdR3+IOBfmv2dULQAwu+Bs1hPWltGxEXCOyk
oOxur4lL7cr7zyjrtkbr7aJ4r6EGj0mxa0KCmK+pRm40txDk2aOzU/4Qb7mO3UzUNDft7YOeVf6k
CfuaydIms8QeRGEWZVQkHca1xUL2y3Ft7lolVPxe+rtCZ9YWnq7f5GyPXKE6p8uK990tQJA2P7Yh
i9YcagalafnmaH1a40dLwJTnnF/yt+NvWYch/IyAgoJ+NjQiaIJv5Lb3At2QyXg+5GG/3aRs9hFa
YAoTt/HBWggkndoubHry8FZk07Isuh2ORw/q0F4UuDZcGGq8MzM4X8+lkGzR9YyeUTskak5pKojz
umUKlAQLpX1hbiEfQDobG10D1SOb9pizsm9cQrUmK/rPz0HO1iRqNnQsKSnt01P/CQ7xXw4glAuo
FNZtjIqnQCxv39b0ueAeePkVZx3bpX+VRW8OlzM8vPMIS2KoO6Braj19tfqBOSJxD1zHtADC1d0A
APtSPK67r/06HwHYhW/pjMJn2bmJhSHUe9YSgdMA/wM9waqs+zOAMCygMxuj4Lh6XI83jjT66C47
e19j86DR01KSvAWnshVG4tH7242jvmOWybF/4Wwx/B9ezruFAuyCwk4fq+ef0NBMrTirRoenEmF0
aWXOXLboZhZRultxB4fzTSqkLTD1aBnXetCLjdOhOtu1tFHL1mPDOt4/LrHtnkNbwJoQeXMS7DX0
ghVsjxpB0LuRJLXsHMxaY34xAgNB0pzdlmoP+DZWJnX/aa1nVXMKbdtcnTrogOyQ4VwO5hUOvJbU
vfSp7JESj7CQ+mBhxhXCsUhn0ku981na0SwOT+otNujjTVDBcEQwVLg3MnnnrHvf4Y8pDW3j1Hor
KS0zw5pissmwzYSB3AbcbuBW9IeKymXzhVmMWe6FDlK4p+O7QlRbaRF1vTx4zS7P8jX5BIxWpWEH
5csd/0f85R+F28768VKJgNeC8E3X+V6Ii68Qtd5C/bwbqxhZLOuHjkF/jbcZNcPaAUmLKReKnwP8
Kl/pamlZ2pD5d2+NN7jgZzoVrBGJiMPkfhjIQHRvlZifb9vfxHyFDbxow7O2bz7oBlsxmw5bcZ/K
oZ9RzskoaRxOJlg9+gjHkN8R4Tsa6t/vWgk3cHh/3z4czOXd+KWt+DuivP0N+xbDOvsMP+7Ue0Xb
B5av/fe/Dz/lO9rfsSpg5YxUauZ3myviiQGU0whs71dJiSzEJsWVkp6gAvFCBhWoaVGsG96ptAes
yEVBP2HJIZcA4Den47Z7bUbe2l62zgVXP8OyIQm/8rouAMy6OnuJP+16EGtEfcqNNosUtA4fq6JC
b9IxfDGjaHEgR+FvyNBbRdvpcIlHL47afkhp7SZ9uSItDI9BbxlFT0hMP4w5YQg2+HrNdz4u9eI3
5lTgZtbQi7rtRS/MXNFtBOyXUd0IGOZn9pfZjhrj9TZxdz1cBLTu3uRiuDxV50fwdew/Vyw8a78d
T0IuuEcH0thqEgX2nwsc05gM3XX1Tw4tK4J7ui/ePranv0G7JUVCM7wBnhLEQwoRfCs0TaEoUO3H
VsMTNAnNO/SGB6Q8PmHvlgxlTrb2FcCjqyk3yyo8os2pdrodilnJ9W1ELsrfwtfRBxlLoC3pJuCy
aAh6QnSmrUAXN7rB3khK98JQ27c/zOXGYiJ8lG5u5Y1fjmpUgUdGJrhKlyVAOGDQ6hdZzCHuj/+L
MmM5jlexlI3lMW0pTU/VNZMPcnCAia8BK6u35893teyiaiHiCwcsJDY2NR/F4OUQ4akYV2OgKGEJ
PQFJmmgsC0jSp2rmngDULnAyBqpkbK0h8Qm+1yjR5ysDp188IamqueLoHHp1pSZ+mfoVVtkQ6xTF
5wDCkc0NV82aI8ak0H0x+8htqgqsD1PQayGvvui4FoZMVIta/aZvyDFfNRrAEE2TsCBwaSeb/GVr
aaO84hi4+XM6tGuzesnU3VRxn7+ML68CYYcZU6UKY0qriN1o3qiCveQpVvlIeTHE4sWVVqRTsLZY
HvxSFhdobHf3N5Cy8uLjJ3zX1GJF+6Cv3cd26l3UdeLhS8DYICgoLTl044uwujbRfhDaGT+PiJmZ
cwO20uGwAJII1qSU5avwFz2suo1wKZ+VysIXV4XP698EDWEHI1YUGjN9xFSA5zWf6slai7SuGtC8
5CWBGRtEXCLiZ23YAU5D4qifyC7mNzqXnpHIqXMwUWxZ7/ZdKNTVlaux2EO9yVMnUSsjnVbDC8A0
jc6FPW9/0O8xuVfVXe77TdsG84Lx7D4p+FA1wSbg/aCSHi8+lVuR4jE/+gS3+FFeSnkIlmHe8m1Y
WtyOO8YVa5P8MWlqCp6owq0y9JDaX5H/bU3Vl5K6qI9dlwpKcT0QN9+BhJpqCiKbg0sbGZiYUJEq
LZAPEwg84wmOr21PLfROcxqxnKSbYB2nj7aW+Hbr0Ofu/PajRlVS6rCwPMEsD6WT7K7Dm9b9+0jS
WXJ2ZXQUSHhotBkT3FWVLovwP73c22gastCSpUsdUlexVI2olqZ7Lc9Mm+9n8SJ1WtUEnVW06LSM
vf6AiXZHfj4woV8JI5DZ+1YzA+BnWSvW+kOyQ+84khsMSsT1KhBgNp5dI+KEWKdxLHJU4CDbNwN0
GYQWHibjLKxakZkRP04WPrrz7t+P4L8qlqsP/abgJE5wfcDpCO9nJGXKGOINsrIc3rP/F8psPGf5
SOOZHjT0j1NIJoW9DmqxL3q41jfaS/1NYfxoT6iWezEJBr7TN7xE/cu3F4PfH2CK0fPFb666gmpQ
PSRUxjcpzak5dAX/v9CHTmSq14Fa9fMJYe9I97mNtCBJtoAHUGaAp92Z5ktNpv7unUCpVQzla+jm
s5/pCsEvsUGs3IcGC8qhW/kwjWNnA25qCus6CrIJJbjalfpJXSjsw2JG3FOUa+QDQKOZXo5Kaim0
xbNOjpdGdEW16pyX0Q+XsBVnvjf3vVXPofAPpTggOEcO4IsFxlEi7NFGycIe5duXkOOatQbWhXJj
6si2w2nvs2q4YjP3oUa0KMeOTu1CVKgpIGS0e2NV/3Y0uNn0yapsu5st11d17wBNfv4KHyzjbgzJ
5W52pyENB/jgA25EdBUHTUr9F0wgrq0B1x0kvzgSusnni2FI76u63GjN1gNRf/+kfVIL/Q+HmgPJ
vQlwnhZEkdj47CF3Zqt63sIhMXyvyIq7PcsvEPddpsfnCEWudo4LaH95wR0JlYaHfiHiXh4Uuonv
zEFP5b4Ap65zoTfjFpf5b8P0zUzPddZlpLY07VrnRMq0lfaHoEaA0b/BSJTUqtdTa2HBCmCVl/8G
L0CvqipLb1MMwF0Htl40N53UJYhuVlAxmekQpjq/W81ChgVw5Up328UmmxAweCO/Z6th3xngYBE0
fdVqMKOtPWImDCfeAhVQaKbMXXYBglI6VUGUgx3Ypl+dkst387OwJPKE/yDLhilhCguXJZqgSY3S
usPgN7+EqefGd9vkCnKyrSOe977yLrGcGwA7eRsjMXe3aKa04k0M48ZkMPaWNbccsWC+4YHDaz8J
IqS2cqgAN8BuGtBm+FBA+xfgkLF5F2kSxkxDoSwzkZB+OdXUildUy30JH1dVX4ZeVnOuPQbHiE4b
tvOn3qydMWEC+UtkOeVwC45H4yGLa7ucPfykqUaMPzw47MLZqiWNnMEk0hPGaMqvLMqVBFQbKp7h
sUpO+k5wyTGwKvTXYRsIztim2sHL/QOpydtvg0LCfS5IcJhcnh02E+bioltDkOrQbot6OhAsezjG
q70N5+BK9SFmIA6ENcSavUV2UYVIlrMzulppV7A8j4iGFXvmLoynGdEQpMTfM7f48EAr+P8BFBuG
NqyN3ALvelNSdO5AUtHAsyjokTtnX3T2eKLtXj0agEycuVy/woNQWRsKpeRAK9S594pCDQef8ySn
0jy1ZT1GstiJG2tDhVM8mpqLMVAqMkYP/2Hk4/DZViGGPJjXpXdvMtlzkgUIpa7OMFsOocJQzIUL
48nFQEZ5vJK6ymOIdO8xkuwIm/ytPNXM6PPvJF6L7y5sgZJs1qpwXiospdkyXg1MeNCMh20hfnXy
X+FtJZfLoowHxUoCkgfK9CoAJcaNoXlzw5g9zDDdS8hUE0uQA0KYwnX13ajZFdSZ+cTQDnd9OF9E
ic4iOYkhxBAeTGtXDQZSIbtA4NX7NY5TvFnX6pJ9kvMOhsvzD/nppG1AARWsWRFzDsjF4w8PynX+
nXHfphRv/2ualS6+k4dXYFqjmIoUuIFT2tYzvNOEDLmzMq9rz8q5MqyxnFbpKjGWcSIoZXb7RD+1
PcztLr/FzYVHdCwHu84ZMUcViVj/abegiw/oRpWPVe/p2LpEdltPznWaOZjH+ybTl48xf6iu1lRK
b6PaT+7tY566FaDRWmQwhZzVvrkXN23fGhOX+Kcz1J6DazEjOtK62zzGn4CVafIGXGBPRByb+3d3
4R23oumSZYwNZPBhqDkTRsQxTv7lHup94U/ttj8NhH2g5u3zZD/8z+p/debkWt+CapFVae1UAw5U
tz8aTH9OnYAJzWqFu1VvHB49gX9lKPXlJXY+6uOmCT/pCO1eaciYF82r/AJQCCxBYTdE5CM0slJm
VOsdZaARmknDz9SJ1xTicIF0dRnkNritsM9NmMze6kJ5LfmcVLofvsBb44TVrg0+WE1TcMEMwLze
4K1mIVmEMcAJ0nt+Nzt68OCHbx3D1cS5s+y6Pz09L7RJtscl4BRk7X66BI/po3H10MjDq7KcnXi6
vT9Vm5335xlTxYZqzO7hN+s8wYfBl9S3y+QBQQtu5SDDQFNdlcAdrZGne3v5c0r4LSDniP9hhdyf
Ry9meng2cwNB4qUebDruhpYC+NGkUdOAKQZEAjnGNeWZixWMqyBpQogvfvbC8j6x4L/1WDpUmO+o
AOT9VZYxS1SUob6WJXZv4gfTnlfYkq7cRExKWTcgZMvvt/TO6KYrayruPCnEXVCPOJR1MzGOHDM1
50WqGg6TcNozJSNIpg12fFQGPDe+84bNRMMisic65t7mh17sM8aI2Xr3gGehmnYvLfL2KF6pbsDc
yut5cqrK3sPVVZhEkRZw3Aoa6LNBZBxuQM7u866fQqnnEzldLv14lzCN93iRvAWov8vLlGy9yZmP
XsPr7aSR27nGGnSI+jPDnNI90+U4bHauM3YCJ4H9IL+08DiMuC0aBh+5mZseU9NE1/mfmIZ0nxOT
s69ypPtTrIkmiOdPUIb+GEKpSuwEBBAWsQyiNFbrWDgWiTL5LIs71fSaxG7l+R/apk8Cwg8M+CkL
C95Md255hp2zcvML40p6CF9jcXGBuhZjpiB3fdT03QOQHFAG8Jtcmo1jAj3Iq1O4VcxYd6IuvpVi
UCF2g2yCKSY+kRDnuj3h8UqfM/8sVX2rsQn1hqfWLCaVdJL1+mb4ISt9G1nFvoWC5YDPi0N/h6aA
GcUMxOljCqHOwhWFFrX/Cl6wVhJ5iQIDfIBW6jw59xCTR71vT6/yY2tdg9ioDycQ/kXlFvF62zfG
CeBgVKAuu0FBNAqYNrZ0KEDyiWjXgUPrtuaS9P4j5KeIivhL6dGK2Kcq9Z7Cg43NW8olKFnQc+eX
UngfIAdYfkOG+IJDDAXaRlXoAgLqs9SX4GqbhMmvvoWR7TX/fTeotZOv1zfrfGu47VPI6GgGIwfn
Gh5GUquqldD8c7J9RFex5Lo81WVDBLtlGipm8Fjt+c/795CNmOcGhfO0sMyKEfg/ZkvxhzEjSmRg
SgnzZ5eRYtNzdv05+YNJ4fMMQo73MaaXs/jQEq+oxuCzx6SWNoPUlIfa+ytWez1mT3o7ZOoLVPyJ
McRNn/xXXHmYz6riKOEjxbQMZpzHqndLIkXDNOMwlEo65K5jaNkTTzVsuc8FFMWOhCulIeDux7mX
zLGFohpQrjberzqIBVz0KdBjgkwt6/4p2UYT7aYB+ySo74bE/sNddbhyq5DnUafrGaAA8FhToeKA
k4T8vMx6zo8S3CM93tinhKUrBx/LGXBbukrduGsD7dWyn/YiHrr+sUtUZuutJlowS9bNsfrXmRtM
s5XwCNG8jW2LcZ9uZ7CRpM9iUgr8gOraGdue31LYrcMKcTVjgVzQmtfDJPlDHGo0DDKjDylG8q0V
yTZtibf892cGYHh+FUexL4s1Bu823l8D+S21rET/nV0XoDSBlFyTiDhu4t6QO4/oDvt32clk9SDp
xpO+XxAVDtaLMw2MP3Vkrw5uYJgQrtEOPvKzF4EofBQo4T38zXEQGZ35Ul8HZOUexTRNi3DXC/SW
S0On0Ppnbv15ylAr2j/qNevzY082ONKE1no1Upj9eoJDNMV4nD1gwqa0YWn+aWMmg1/4/OH9A7SV
xw9SbrswnueT/lxWW7QybqT+zFv5v6ZVrNRqkg3hWVCrbZxVqlzKq8UQbwqqNpB3fOYp+ln3c9Jn
4UXPCXUfrMayfhkxmGo7l6+yQHrkLZ43aklKekSqWEFDiYKWoFkb/SALXh/qmL9DWdq5ZkL0mkac
4qp0MFxRx+yNTceRBXhE/coxzN77jQ2C5QwUVN6ypxvaOAOI8G/OdQBljNccucsHxOqgU+VdSdW6
CPNyrHGaHGQG/g1YwhsfcvCgZIIzdnycPWeigosK2E3RvEZ/DoT3KHkvOLz6ca3YBPbqB6uqGrby
y8J07L32Bhiid0GGRPcjR1XrbfpW6MkYKkkEyYyQCaXzxpmssclQHStFDYuTTZZi4TXMjvD65T6s
1bGReXQAShokXX2YnDS14GaGjI+mxlYXony1gHjBI+3E7n6mGLFBxCSxYY3O5K07Dqs3c8dyZ2zr
lTv6kphtKQl5CsvnKCvQaAz8fPEDYtkWx3aQhHj16eZr5LVBoSkhc+3ybjHrSQba/1Vy8ZX9o7vZ
Oo5jkHGLJL+u4DHuQE3IQ/5Jlv1TFU8KA3YcByr1rJHzmG6IbcNxTPP+t1/PXOzgAwGqYjn3ql0U
+izjWfHVGjYs8UayvgL1W+PuKCO3gG6WgyE68yf9MSfAEOOGlY0o9bGwfViMrj523gXEvsFIO8x3
BD1l7AWFk5zJlzjyA3G0EGxI1SbPk8zQeVyxTOmpLXGr+YE82k5wm/Sm8nd57/HRdzlgkILqIMFk
FOr9tlW4yiREErSaPWEWuhn3sdWxzXxPX5lTI1ISvac7D/ry38ie/zMf8GD1+xpROlLSdEpYjTjm
dZT+uk7TNyCTRH/lAodXI9bHAdSBThy/GqI24x0MpwlI02YPZ1lVIiubK3oaPoliPmJZkM5rT6we
tHgXGbm/L3P9Etw1bXkWlKqyilePvAsJMj21ATVPBKngYM1YpdCf2rEcmP3I/iAkpSJQvNsuXGxU
FXGZ4uRLbnyRSQ+SBBfqEy4UrOc+qY89qtbwEbZG+eP19Lf/aIQo5WrAJ9U0BgDqhuDQqSmwN3kC
sAq/O64JHRoWpWvnGUP8f+CT+173T+iTOWTtNRpYGjumP0g2CKil155J85p2ezu5NFB0SabEY55O
NR9gTCOBHqh2MXkjUod6Hxjb99MmRB5e/bW2nj/FdUe6isZEUFqRTt8WdhVVmKI/ut/VT4SgqvlP
Yikajzh9oTundsT3cqyd6CRiZU5uk8YGZyXR9d1dEHEjvse5dflerxorBaV8AGtWt/mZnF14rqk8
tcagze9GxMlfdfHjspC6omsHKYIFWVT+SJMEOd8KHWp9h2H0xhv7J5sVTS5+l1tbhypl9iq/+WB4
kWHOzLlH3sSthJmuGkuC3WrIyywcHOaQUWNTp9tOK/CHjFHGv2iJR3y/JiBJr4dLsNOz0fyBVt0e
Q7M4snGKi+gyWfAE/M96c4RGjHbEj6tSCqh685CVsm8VynbsSToBvS4hP03PKQxY6bMo5CGasdBM
xI0rTUyo5Tpyxx2reUPCI4bf+mARJfcNT5BCam86DQ5wiQUv4wWasirCJwxRbct20hab5NnrnQxj
B2+OJ9rJL1HhbJZ3Soh6oB8YROcnHUua+yZFY5NVGt7Cx2Y+sbm1T0vw7/reHcuV/jhqyoBVgD02
Oeg+ZJRuunRsOs4Z1gWyt7exMa1NMMASl/kdcq2RPjeSXdUKEp2gD6pMb5yHI2C/Lw+/O+2EPrb8
rBsSHFJBST+RyLUxUi46Zo2fOr/g8SwZOd/8Qe2cPJqzsHz/kl2snWlQ2IgybtsEjX7fJUcq2NPx
JIvVVTnKifdQ5ugThJGr1jpjBXgBKlJdfulOTarW0yTwC6OJg9/gkl8kzO3/tyTRYKREuf96c/k9
urLIwzoawLumwrb7rj/9krVbjh+lj7aLkVURGYpCfQkS7bfH8Ut0198HVezP7sHAb9JUKOK486kg
yW0tEDisy7jesePCauGcdBG1SgwAYkTvzWtvUXv+CubJwVz+rp95rjW5v/ClsW9KKLOyxKPaYOO8
NCxJZigaAJLsewZYPhCwWUdoz0nRufxHGKMmPC2RCwKVUcTQu5f9LrnB247Re4yDt17BkbCoItW1
DGap4Q0iWB78TWNhzmehxWpvGXEQUtJkV32rUjbBZFjssMFzfsaafGrqDQ/f1yqO3gC8DYJ3svbl
HouCpA0LcDvOsADISkm9L2PratrsLKvVUBwLc9XLvbVy5ONXKhMKtnWvaF4VXkl2EoecR86U5zae
Xwe2PE1HMbjoyKZUH/BVgJo29jquzlCKQAh2K3pDXuLdQHp/pENQWuZBdXQVnSRLuBs8YC43DvWX
kSAobdhmyJZb2DvvB38PjU4cUyq+hmNDDc7V9d2N0dKhvyQvOTOs5xEB6qjEilWXxmZiQIOYaxdH
AYpVmmybZIpNshjAgqqLH8+1Fjj6AyCNaR59h1hOoSIyN46HgY05JRv7cLL3KHc75xWIuU5rsqO+
2ZUKbXFuGuY97DtZFSbGRYSUpwvbLb7mX2+Xu7Sbvt0hIaV0qgeE1tZwqjmnBZig0J/fz2ZPoTR3
11mYmiLy/wUSx6WPavgCzRGrNzHVrok8CmTDgLbTlJ4R6UW91UYjfG7qPZkawHZD24jcLO2ST/V9
LMvvGKTl9VBd3l+w5hHKiBwnz+WpT79+odBzdwRtDQwuzU3Uuo1rF4qXy70Gb2YhHzVoES+DBDLe
7zhauiQUPVuQIXFQfkuwhprYkfEqfQO2m7GXhAHoZ+WjcoOwKJrVxlG5grC1R190DVxl/j7luCZU
JAVnrCMbGv8MbROx6Or3sZ046rXUXisPLDD37QIu7gBa/QA8MCImavPxbgCKmz2MOFW4LusesAox
mRSGHZRs3VaCqtUE9S83NdLN5f7ZQQlL3cuNOpYHo6pMe/OmA1laR10ZIIf2Fr548Bpih6QSQKK2
AegvNitHhCQL7gmMvTk8QCKlHTObmYSuAjLOW4YSgRrwH1qgfh0wE3tP/Af5bl9VtQqEGRbcqxH+
B1upDkzgyu49Z0qw6JGnT1GuYKH8PRdPs5BNl5+HoApRixF7yT3ck1TrmOkwRbsjnKuPCEHOC52C
Z6r1FI+krcOA3QnztG+7wNhL38S/Ni6uki9+s7z2j5uVO/W423jW4XtG4M8DE3nTMLhyHNRboBOn
og/776TI5WlVy8qal94IRlVYXQFhTGEEXs06qwzshbFg+JTQsLQOgmfCZba8nCpUmJkTp+NIfb89
Z+jlO3CX1RxvDmU+zFRPWioegs3C1SU1XP7md/u8efQgLFuO2BS89fw6NLIlqjgoM4unQ3hkwr/F
iRemtlYIQY5iWTRJUuJpcE6kEL72HOmXUdiXycF3OBrOwh3BgW0wzh0EKEacT8UJWEC7f4UNVQOo
vNXLCZ6MQdL6EHuHJLgTuAnL2LHtfl3cx6ng2ve9XKTiqmOTkGtnI2EBumxO0uCcPwEzWo45NYlM
DFu0SYaiRZ7APJtL53VJUytZ+KdUu93iREuPWeKgCzXcNG5TXPjcKmTZbz0IQDKi/8+i788EUypL
7/4RJ4lG9/xMODUC8g55RIZYUxjABw4QtmIXlSyZGF/XysMm1V9ZAWPvHz4iHvwiRm4VCwiGV9S3
mHdKSTVHqZCtadAOogVIcQM39StLbtKDAjfQiuo1OBDL/xal6JRkfV9PGpEsXrYzne7aQ+NLf56n
+gDProCTmBDmwwt7zaXBV7SDCK+5/sChlYCaIOA8kWIUN36AA46rl1ZC/DPZfty4qj9cbItez51U
SE9poAfbEkQaKWlNifZbUMvHf+LdWgkI6yrzU4RZe0lgL7VE5T8jhyHpLEeOU0F8mqwk4SyojPt/
Wf+vVHjPwr9yR7RSIEiSFicGo4InccUiLfRn+HYjYNfZJe7F2qbnvh+kbvRRtUhF6FcUD77CwVDk
JAoopzZeja4TSMO6qGHiM7H4do7aj9reiC710n0LC9I2KGM/7LLPJc2T8jW466QyGUYEH6OozRmb
20T52Ss5jBZvv8OA9wp/69JXabTX7kpY4l5vYNz69rww35dY86qam67bFXsmk+kzNOZCBULIvBUX
a6jKQGI5RfpAu43xbENzlKccNcMaRvvZUfArWFUNP6/P/fxjcTNwG/3pkJ4R4YjMoraK7zSM31ob
sPVl090a4vpndrC/yEMGKeO0gUOelGgl+yFBaQpbhGaNUtqow/CRaETrveUGLJiWsSupHnLK73tL
YBw3pdNBLTlqKCZw2DCwwj9PPOeYmQUtroZydbIc/rYxscvyOL8FHTDc+h0kv6fsyAFChY++KEY+
YmaI8tPAH7Ad69Hfd6Bd1EciKj2wOAXlUy7UX0++sjlX7GKWYLJopJCbzzMPUysURyBtnjOTmbD0
t2Q3OAnCrhr4Yz7DWaJuD4TdPxy4u5gWN+BCBp5RUx47MOxUirawLNlA5mWPD51sdnodA69xwZaJ
Iw6fNrRNTCykbvrDsB8VPeBNWpH/U6IKqfU9nFBd9Hs1Dx+iVubAywNLMpI1RFJ7bvdwH7VZKHRR
JeAl8oskCGXEvn8jfxAtWD7m5HNxHuav5Ya9ZB+QNnxt5F2JKIoKaJkEdbBoANZdeWELmYJFtj7c
xmJOaox/zdDxE2YfUxRZrXrp5SzFNp+2nJZx0kMm6VJB0SO8jwuO6U+rl8VAmMgjsk0eNMAh0Whb
OIRrMr9RvMeUa5yZ+DvyuQw5lPxG7zcXovARoksQA9b0p/U3d8tiDAwDhohR9zo7LAa4BFLMo98z
FHz1Tre9oX832l+BtJRvs7b/40pTYjZ9o5VOnkiniPXSF4tJluEdUFzbQXq/qcyeK0kukTNhDdys
PWEt3UBQ78Ue9jPC9c0MMHPb3tEzBq3Cycnf6NsShuY/uedZYCizq7M0QsuRRvkERbljC2vRmDa1
vkU0XBnHw+cFAKgsAijxfCoBhiGz7EbMgKBXV5eapd8j5xnvROQLYH8D8epR+n7+iSA5Q9osV1+H
jWVQR4yOe8A6H1/EtXGpNC6c3Y/uqHDdmzUxfVfobmZ24E1j+kO6uzLezyfex38Sz1SkywiBP4Eh
VQVrvEYuy+wvaRrkVyMrMvrJ7JDXCbBlPOvqUpd/fgBDyJgr/guZQjf7kzJ5NpX917Cto941AoSP
HBiEYJMPywVEjcrfqyHOMNBOZ74ggZ9wof0/fSauDPzuWqdIhLQKcAuXObeKuKDFFEv4q3iHsg7T
/f4XhRv0vP6Utn6+eT/vUN2uGT3mFyi7Jca3hTX+DxVQN51IRwhl9ZsTV+VKtQDXXyu86KEwVMgA
IAHJMhqsfwyL2ZkpZ8nH/gT6o58A/+V3zQq34EAXXTr3rnS+4oPi9VQetL3rBI0Z2HYW+AfDlq6t
AbkuNKvLKYC+q9iRXPbm1TnqejaRu1VqcQTaHqBVrZXZerA6a7Lo0EiGQcY6Yk7u22uJK2laMXqF
KJhQt/Ev+6tXBOlhLWKZX8nandUVDc5IGrdHIupvhD/CLYKw/lRJEcNRcup8MigRYmSBcyvHZ4Fo
7iaEMkLxLPvBffXsBrS5/+Lty0mzKfRi1RyQxDw+PtP0I+uvcjAqAojxAfW6Vjnlplh8shk6Hde1
nwgtmLtHRMyW2+0nZMiEG18Tq2rw8JehenpCpKDo6HbwDeye6Dax/FiPsCPFmyEHOk8+0Pt3hbnU
3KSx2JuZwOhO5b5/LgvbA5nzSH/cG155Nzb09SLwomVT8eixG3Urc8aWPDpmiZeFuuxnKACsdKiz
25ZJnKol0qmKLnbDxkSj5oSfIyv5il21eeAkATJQWKw8oRh0Nhc+vb7hKMfEDIrbK2GdaLHlqpOp
xnzQ+J8sgoRJtZSIDnlZAJFA/shuskaFkrcGF2iRKay7Vg5dgo0WhkSWZAuwqnotGEt3rYkBM4sq
23ye8T6tE5vhY5N9WRbs7MjY/zlgEKzxfV03FlniPecNLvUiqKGrbvRKXGr7k/uEd6tm7jOt1vKq
2gHgjh942sjtlcGDCOC+y/W/J0wcvA1YiWJpBB+lGfARJioqZUM331B0ze8jhNAAb4b+YhGJY5RA
DFY5TPNMZhKolgkBwWYBYbA0Ax5AlgsrGPh1GPOkup54KFb9LkKWPqHlisRSmjVTNDVGZAC15RQr
rHBeMVkgIJ08H4AtP3bY/Rynpt47Ht1sEkvKso3rZN7KIuSwLrkWhTIOOHBfUuYkSnjauZ2GHpJD
PW9OYT1a3KBm2B8tXaLPDvfnGSeb4aoehuAQ3fLDRBMwb1nX+JNAtFtSOH0Mo/p3wbu0h+idS58h
Z2aWBNcnplUcAb3N47K0lGG9xTII4pBH2w3bVUmDBQVXJMghqgNqFGlBLzl9VWBKLzJX/2/IF0T8
nHi5kxdxKzNGosaHFr7Jw96W7eACZFCzfzol6i4T5hM+2s5PorcfxtdLhlzab2MBqrwgzgTE1EY3
2YI+TtBBDy6hJt1cWanUdDR7M2ICtLSx3tu3qpmb/uhnP+5ylaqAZZ7elM7TQKnYckVCX54/y0nP
HlrOHSpoN1t4CjsGaXghrq5cPflwgcxUkUghEjIx6YKJ7p3rOgbjEKxKVF7XghHeB9cWRc6JykiS
dKnmGir7AhWtOBttmLY/ihIvg+5BExiVJL2/Ap5+rW0jIV5pJPHBhHa1FChaMdreHaj+ihIn3smk
hu6L+C/8xAy5IWSJaCmzTVaOwMdcx7GonOReruv2sklP7q9pJ7tF8HNXYuteRuugPu5F4pnzhnnl
Rx2q6W1hP4NTYPUg0UOh9Rs9uBKOrxh1VRoaQArk4W9JvLntMpaWMtchr49G7L2ZN0XkZOtBqDeY
0XVKd46N1lRAmGIsYPrIncYVECslCmZ1URklnUIU8u6Eo8Gab/XoXk/gPk41rgAtG2f9cSwazV77
fsOTWk7Yy+9f4VUwT7yPkscfaEcgmXZN2/Q9d7HmFWdHrXkHdzkdVSo7UBeKi4dS4+eE4kZ7tGo6
phSeu0euVIEiCZ9/gQ3sNaoZZlzmF5Ai7fUN9d/ASAXGV4fsX4qZ17M3B8ba3NKwNI8zfFXdcGZx
7Hho+/Zx7OvD5M6e3sTlhU5Eyo1Au79haCII7erexVGkNHa8mS9CTU5T7iVEbvjhmpmm2R1Dj+Zz
xuK81anlzvA0FDvtv+jHG8SmFd0vqjc9qKKNgCeWzrAVMBeM3AK8R/9UjBBAvymETtSlG/ZeEEO9
Z0+F0ALQyGHt3YLpe9HJVTnulloEu/NEzXcfaB/myLzxWZcbtXv3UNbi3+hFk8sksx2XPeO3XTly
oKZy6r3vursP8YF3epmrcnmeb2z9MLG66Ed6nU0radpu6wuCUvK3IO+BzYddFqZQv6FIQN/rpG7I
pV1T6sSeZuN+t3QoaE7hyL4cgy0uC/piD6N3YYTn5cawxzcfGf/X+JI4LvuhptO+y3EkZmmd6fGq
0r5/U7qVlF3F0WnT7QtiwDFcxAr8YsZZ1XXcAKcRQLRc+l/zkZDvqRIbVv87xbGsSlUkB9RQrMSO
ld8lEWYpQ3lg+znIm4Ep+d+mdl5LM8enZ6hApPH1AcgciSsyx1BpCZlQ3tP/LmgKYez2zx8AgPob
ydKmUKYyuXpiMpwr8ApOpJDjQMLA/07efCu1VeAHr51+7TTIO2lTr5cPl7tP1xusjO1c0c4LVFF8
ja870vRI1TjjXjLENMfnNTVJJXxM6x+Wr7/cIqBspi9REFuZtoS+6IkSSgTbTg7fgRDQywaNsIdt
BDoLfmJOMEmi22Ihr0bASTBSgRHT7KEBBg+nBdfLOBVZA1/5jfpc7uXXMwxgRLajD1QvJZ1GsmPH
FH40Zs/FFaFeOB0dphOblNTT3LqHQDSAbXvCouo7txQRC8FjvTh/RGw25Buama8JUovyaywvOU34
qRHUe7K0S2Epc7lgh8I3Qu/umwKHzR9bbDDfHOKbLPavfH4V9VsDmnvxHijSeL95VK3Ri2hn6eEY
VsM42QVmVnFB+DMjs+zjY1saaTxEni8qrFD+33UVxx5LMWnLgu9W0cLDH0BPcaLrBAG1zLMJQmhw
U09S4YiWy4+0z8+/Bz8I3tcbE+c47Sw9tUv0IbqNZ8v8nl+dHpmG5ICIOK7fVj+Ew0QI3XajT50r
bJbkjjpJ4MXbIDIQ50m1IZvPY8kNL15YpZ+3sBJN+DyhjKEv9rMjviLUbEjrxC7LTSAEdDJhsj44
kSafeFzxAB6V10WMR2xiPiI+eVty3sXjxAxrDUO5vI1h1s5QU3T3dTToQPmGKwa0SylzT6eWbevj
DEzs8GOJWx5VsWWjcckSDyfuoD3R9Rg9npcfH7N2QFEVKnXYajzw09Z5jKkJsDQOj6iFlJMIJRgM
LAxCNHJ2cE0DRH5gPjkVChdvQIA898tXRBkN8FDBdaFZ6nrYbJ3yipPIKTuHgLV1GjAGyz65mItc
DK5oX6MGO+7dGyn916wttiT1mEz0SMTsyJRXIQoV1H5lJKT9aRmLnhgH5D7mo7R1oLVifF6pI0N9
rBRE2PADqH1ZeZ63Dhwwe69HEc5QSWUI6cKJhPZ0KSIChmWGoUKR/oBsWZYMH+CeH85DHe/zdnDd
iy+kwIjbMHG267a9YYUrSsKgSfQy4ysvIDGABKBkC0gPwDAogKXPk60Z5EgtKlSFbX9L1iXIkX9g
m/hT5b5E4y8og2WV3v8JNmeMDUZrv0DNrpXXqsa/61XKdzOt9OvQX3ZlvNCyiJ5UPi4Ho+y2D5UE
pK6ggfgNcGJ9NFjVFzF2EnWVySsq+yxhc63j8rKP1a3FUrDYETaaKdc6rQkG+1tMUGHSf04NN9rD
+Ad8Mf5/j9VND+28AgZLKpjHnqUwiXDkqsoZ2PJ0vaL7FtaZX3sOz1gg08wpOQsSTCtTA3egqvNj
BUlVOQiIslL82ls06OjJcZrTQI16IO696gHqQAA6DaatIhZrJP89lC1NHS098/LniOV7TZ2KR9NW
endQdv78i6z3CK0Cs67jqOHKiHSFEEbYgox/UDmGQFFVDn+PNV7rL+yC7U3CGaSMgjwcwsLpU8Zx
J0YGO02Kjb/ZNP+rqbpJQtzGXTVAu7LmwA+ct5o+SOp2l/deuk9oUQ1EdO/LkfOdVWewHdV57IsE
35ozpEuNKAA1sFDapXRMYCYk5KYbXtlPsysXzq+gLfBeHE5mVQQQFvOLCleyGQyIBD5HvZHclqA6
TFY6Ea73JSFQEq84Mz2dNhSJ8sipylgIU0hPbCeR+957i22C8qIljrcfQR9Ol8GF6II6d74tk6sw
F4rHlRODvXDNXPDLho8FqnwFl/UkTqNuXz9HQKUGpNpYK4JNvPU3Xvo4WzNo3zxIne29xXK4V0vu
GORP/TW8l8cou8OF+6n43hLcmvpCxlW6I3Klr+YB5uh/frjCxABx4GKOQguCMPuo36F02GnOLKMw
LnwbI5JDDi4CUNqdmVwTaUlOtmHqcWhJQGdgTHe9MzbcfX+ANH6gZARJ9VOAAYiqqp8VTuOl2HwR
xw9pcUF+3lI9e12YSqya9jGspm3f90fpzJiMfnDRP7kl2TZcsbBwt3aYIaf9yD4IV4abjcJyAGWa
F5zYji7Cs7+NwlcbyhJHRUMcT1/cAfR7XC7kpwtg3yUi58HbJwfFNnkYkD297rQpzTOYj99JIMe1
YO6vmpplvHTafzIwG/2WoUYc0gICfbG8LtmmYh968Li7G7MqNnNeb4x9G6MHeBq/QZ1P53d2wmMC
kXZgZdISRTMXpG7iLOVknQoET7sGF9qm8xW6bvxRNFGL6T7Uq41h4GMSQSuk2Kv6ZSKdUuaA6/ov
0x3PKGTiHPtwKxlEUCJ2qkO8kZNZbQGAQnE+EUMXYBDNCgJfQpFKIQ7CZIqo7RUv1ysY8nm6rcIB
sGygJwt747Mw/aakkNrmb1g3SrrJgvRNb1qLt5kMyh+WwLmT/q/OUphnUtxK2FVlACe+NzjelV82
IkhuOkxwuU7NHofcpYrx+IUvEY8oOGJN9yiVs04Zhtw+1OZbUfN5CDDgzGykGl5AVmu3IQItWQRs
EeaAXKCbsnMxPux2Df7FDSsPt7oa/+Ewv+FaL72gT72TNU3yx5eUf2ctuj3jCb4EJTTxs9EJweIa
/Np7QoE9C2jzANJqZbmKcbxLWvdGedsrNxfsV3SSvk31UqXI/1IJ0daYKyCQnhJamzNIwmDajwGT
EbZyHVtH+gDMmNNBscL9rwj+ojtSGECzWxKyVtsL6CQK/efd48M/m63cJ716cvXoAzevho40lHlM
jiYi36KLJWBkilv1+RpUY8Ni0jdTCDzf+bDBAVfJVblfpejcyKtkn92yytcrlFzMCR7O106yYaq+
2Yf6adGebnI77PckMPmXzGiHUA8Vb5TkXeCMo4YBGcZzs4wXHiqNIA1Irb7Eai1+MzaLHREkSKGj
txfLjNPBg1eM8xMDrBlOJAMcgmiQaVGRwk+c2SHcKTCcX0yJLhNhbwulTvqWCmd4HWW0DXj20ten
FGgoEI4S9tDZFfLgUz+q4f61TMRJyAXKrmeyfxxETBpPWeCgfbKhzjEgew1P0pGOqlGSneGxnj/b
kah13oiaHGEa0oknGEa1aPmnKuEAkSiywgGw6gUoKcUJz4+P8QRs1proCg8DG2736RSFFZx2vgJ3
DAkZccyylhwAK/CgEmP9a/N3iv5pRl+WvN7K1rJGYduvSzZVSKt1uDyKIlrj+lJFr7vpVTBUYCHz
xLO5sgoTszkECGTzJ64danEO8NhsjbU/ZPlXn2nveuODc8AUKxqCxRko8H2gJAPDIDVlK1jIVp2X
qDrj4OCsChsGkglT7j1UHDrRpS4zgojkS6bSEkYcTdau8oUi2CH0g82vRPTvdXSomWnSzXMC2LYA
uzjass1eHfvpgmELrm3wGOPSBWr16mdtOFYZkpFuSJ8amYrHEZBnZKtG8a74obg5NR/Tx3ohkSmV
0ImJxHmRZ4fy/Wr0p8fvsPMRw/UGjmDuV4Hr6KjTz2BHR1BI38Nl6e8OPuo7xQhxgLcJj9lGBn1L
Nh4pvxzlQgoCjvB2f1soyVlOcpdEKdrdFzYjSqTfYrDOEgkJKMr5zNAroDG6YsRN3a8SjwR+Jfqg
JBteBkYmf6LxcHI4e2NJO+IWKAPA7W9v1m68v8hUfF2rywOd/pRGpikAqel1lvJyn6EDrqckrETj
HRY+ssyImG0UrJuS81vWnS8sPsROiY52wQy1iWfvgC0J/FpDgprRmSSJKwNYZwCZu1uYV6TqHdDr
473Ux6fX6hEXJ4mD3x3q/LJiiBBcvorsVKs3GaOdLHDItLaG6kaJnFfDDcBvmx2bLKSE2c7AHzgQ
hR8LfDtbTQNl6xR+qX77IB0HDnI2fRAj/GFKOR1VrOl4xMYyC6qlt3+1xswW4JH67f66AY15rmZX
9Sq3T17gEt4qa/7XgmYqk+ltXpYVCFvhoqFneqs6NtpEW2MP1zzLa82XgWADima2nA7WnxdfQBsx
/2oKV79B9ALrjdTvfHFPHWpu6VxmhBuhLIDvym/NyXyA8w/S+6zva2WzlEcOkwU0m9agmTJWBJfJ
ftmEQ76Zs5me4MJNf5T6J+yBuMjhmcHt/rleUs4+qwgapMHsEc8evMMpEzwuClYiFBmRk47Avswa
te5nlpx0jyJH2gBXfhJpMGi3HoBdJLE+Wt3YAqdS5aWmpiNWHZSIGMWu2cSSRwZJ81WuHT+/96ge
oVB7Pr5asNLtiS2DjnsaWeytHPz8xAoT3t6wn+JOdkUpkXw+LlOv3b+tihF5cRlTd8A+VR4Oofxh
fXU1mPrd/ql7u6C3xhAvjBocqwHxpFWHsFDulYRpZwEFt5rFY1ZGWLEC6EYOc+hHqmdKLzPj7EfX
6enHskSbGNtGgK1kHkGk0iSqiqjogoTepp4nd7GyfvsyZJQ7/2w0QYCze2uNAYrncdD23166QAi9
+bHKV5JM5TBsXB/gnIvwyY2D2aF8Z1WWIXs26MTDnFNqW625tnbpW72cuQzi6BOXRAaySFXO6q4w
G6hUfcguh/c8zGweakdkheiS5v8NQyLVAx7Dn5+CriYB2cZ0axXEP2OxaX81QWoiztzI7ignmmyz
IkBJyIjmaWf+RWhu5RK6dV5DxmmvD2hxlL2qri4wKhWa9GoL1l2iyHoTqANkMJbYmEOifyoxKydU
TRyPWriPJCrscz73moPedGb9ONy1B2jpy43q9xtvigUzYi6nYPM9y3oAvkuqwyadrn2DJpwL0FNo
9o9sXNBy0h2ESkCc1pRKgyWgmwO/bQ0jkoWiI0JeyCwl89RL5UP4LD+eXMu37XML+n99HuAL0Gnc
1iz8JRLCO5yntaXN4rlLJ/WwrC1oJdICapX6/LYDmWy8Ii7oB9on+K3u80hug5LWda77GOnE+SIW
4wHdYH6AyVYqO1IqE9t034BrcVX4a+3/Vu89Gt2STxHb1P0y7JAo1LVMYiEbpiEq1YMkZ7JrF0lK
M+cpA0Bt4Y6EZrscxaqZHUOEa71vldhLruh6xgz0btKAbm5Fn31dTG6tjSn/sZ0eeaHGrU7hAu/A
F6vylJUs7Z5ZF6hEGwVPhvMruuJqxiQMLbnRKbG2iaYZxGjzKQaI8tAlwnhI1fCsS0IJBcAd0SbZ
+qyKsm/bues8HzGylOGChL6c5BElekqfjULuH48WkopHFpeimfIL70hteIv+apKrFYWE01gu3mXC
rLPHeY14JBQ/UBnNelLBo90NChM9JxP3Seex58lNuPWQCITRah3GPeENihEhXFzFv0nI0srvuGF6
9qcIfgjnUM8YEpkY5OHNofKNLyKUQyGbpEVQ2DAFc1HU/M+w4BXcFpt31yJIX9telkOBxE/Acplu
J7ntpbEwJxgmH+9A14wdgXKd6LidGfXRMw95hKKDxRjc+AA425o++8wVtHWiW9vNJLPgv61gz7fe
WG9EYTm/hKj/61i28LezTEOSYCFDSsCqrVL3BexA7RwuQW4j97+RDHl9OEtvZAekVG6ak/lV+Pex
M2uNvGZ9e9ym+lNo4a568isfRaP/gczRi48M+T1rl0YvYbXk5zGUSWD3/CXGFe8er/kQDtNj13xQ
AhJW1hG/ThFYhhduohk2PmRjYzoj83zRkeIfDon1kE4VE5IqaLSfQ0fRdox4PwRsM1VgAVA5dG1R
dHFTPRuJBEcOyfw9ekJYWZaC7qyZcTzizKVkDK3qE7tQfE8uSN2Wvc1SLrx5COmE3NFAc2XJzoWQ
kAPuMvXFc4Kh109Za5ZmOGrQq03vtsTxEIi1B6lar5pvNVXkQDq7uYPQWaphOcxSjkbcHw34pdrA
mlFNPiQLvkwXAlGPEIbiUGBL4jYgBrvPK9HsQku899VoMcOmn8wHjy5ko93gKgus36tVAnMRIZSR
V6vGTymr31KvsM11wqrs4TuAOBhg7U7/xOnBk4oCnAnU1jkehNBYq0GhCG9fxG/zPUrJkrZgAies
iQiDWyvZIEd3zCFnzMhLBOr7EjIETN/a7ljVd4jYjSfw315oL28hy++pUHtR0uybSFcWwLHl/gfn
hxJ5qq3waEsbdlC8SQu29ZxjHqz+tj4SpdVx39pxW4n5vK6VPKM3K868749l7fjIS2AIVqH1yfQy
/4qWjvoSTGobZ9SFY4jEkmyXlVLfUO2ijNRtcrGY3zgOl5OE7jEIm/hPuZnkeV0dCw3ul77do80T
4EYkjUXPBQs6G7mdoPKoQJxr0QEW8CGItkdZuqAp3JLbhzTmjIlBt5Cjh5Pg1MmlMHKA0GdosWbA
iI3q/Bazr6d+LRK8SYSDJVLa1IQ97Sf6hIqauHGopxcoC963uze7XCWbSRACJjIvqgTmYmSyxmnJ
hnz6YdjYl+u4P5rMjlyoJEiZFcs0PuS1A8NAEEbcWTmFk/+qrPHe2ITJ4X4hfdmHYmUPVFo5JSCJ
Mk7ThXiIVEcY5Wvafju17hNJcjWR+KneDG2KGdTvyNaCh4sNCj0QD/+d+SVNH91jRGrQFDCZx7Kb
403ErJ402YK4lA+8rE3hNqe19x4xYRuzpGtB/C9oyIchAxk81r+Z4zLpZED325OrcZVF2YYXc4d6
5w4ofhqVsPR2CRbo11Pu8iPaCmBYC5nZ72zF1l10RP9dybVGwHbBsV2J+YChdI/YeO5QxDAfmMlA
Z0pGifUGf7avkUSOFCbcB3AcaJGwBZM9T7nz++KlQT0csLFP38VGCnJTirpLUBMFPJLrI7W8gEBq
qdVbRKszOCaoe1KnrCiuEbSPHQjok/yvwEKNqlRt9qDFGGUtZA9tKD2g1PNQEjYO9Tt9WmTYAIxZ
RN5gsWmwQ2eETd8krEc61uzBRh0fJktxKTatBV8MyC3TG9E1+9EP6/3GsTV3k9vjz5BuJnR0PLNU
67ON4FzyY0HwHhSbhSFRQHmCW4ZpMEeu9HcMcND81UWX4Uh2F0G2woAEqQZ9fHgkykqGnwqd3Z3c
IOvmb1Yy1ZjvFC9InlhdPhgx/aEyYa4VszXA3WYUZscTXq4SuprZi8Z/t5t0fMIIKcRD07s29o/X
5V4eVihxO176fDlH3H7FGABV189KTJ9uf8NiJ5gge0ZsEKD3CtANE+tew8gx07DIA27SIU32fkqz
m5OqQFNuZHG2xCBjR4VqBnqBWgspLae1GXEHm0cCzGv1wUzphq8A0lZrZDEKov0vzfRVjcsm6z6f
Tlos1stRIZe9adg095TUPN/wiabwSE4IyksFnftrBKVFz7FGTm2k34s17YmkEi2GnMPTRYt0oavn
dk9s63XtNp9L6X77ggs7hqmoKmsdoZ5w/8yP4Byx0sl5fBr9bwexsDoHtwDtBD8rubmC9BE6T6un
oCC3jJrgydoLEvG2NCOYc8a5e2AVsr0zAk9oXziXvDmGQSWD2GbLuyOge06N9oTvkxzFXXCVG8zp
amoBskUASanpKd50XnQB3AWAgejdLi9iLxPfOYRD6qf5vVbtWlKiqJAvSSpHt03Is89KI/85/wXT
r+064NlDOOiplkEY2LpFyoQPaeJabf8+tiEWX/e06HsQZD6l9ALZEfLGPoWMyFDe/3xBT7kX/Inu
xwuZkeQmvlbTdtxGs5Exc6im7rvni8t6tS7qcjSWskylRNpUvjANKd7WQkEpDv3gFMbguu/PUvkw
zzTiFqMYN2xYHPyvvFRJdegigpodPAU9tYljQF7WWnHL+8saOo0BzJgzsR+JNAMLf5cDF/ohMN64
+7LJQn5xdiC7PUWmpAo00rYcJREpgUMZRhQrFiO1/s4VrO0c+TEXl7yEnKWMq+uBQqc8QW5kE8gX
N7FQb6WlfNiOM6/oJAqhKguMLbjJwnFhgkEwZx8ySKeU2Fb5Suhu2VxRDiTgKENezLmcBTjq3Ws6
encaMFHPFt18Z3MVlPIS8sW4ilvagliYu/Dzbg+089ia5imM1SaOBLqT15pKZVL+dEw8W+5vtzqd
K5mPV1b0+yHmcs7gLUrqP7NTNlBQHKfgJOS5XrBQPEzZEOkoVUqKwQA4iQT92fGbfusHbJBN5t8y
Sp4DZCBTqEDh2OD1xdWzciJz1UYhCIN1vjOmgfHYCqUx8jUEN4Z6XX2MTevxagrptQnI8F69EFjb
EhRi0BdAfSAsSz95GEKPJjI73oCZi17Sl5Oi2eZRNsdOSaEjC3glgTCEK7Sd9cXmbS8XaItkgHKd
t1w3WqJxukAEuZdwlLpWXKx5tEp3o6PlUdH68j8oMZwsQB2JC6l6nOf0291YmjG+ZyQ2p2xs4YmG
Wetyq4T+jFmvx9oCdub60Vh8XUCk5s87n3Lmq31I/Tgg+I93rVVHdo3FOU4pbT7e/Sy8zxDKPhoY
jNzwxctnEB8tqCMeN+lEUAgyEyfo3oaSGehOBcPkrlV7bE9p8p3gRXb0NDHw8cClrcXgaiKsbPTe
wVC2YU2FPG00v7NdCZkFtyiBVF2L9mL/bSnR8BU/dxT9FxvvSCVnKdtFzgwuxI32N/EiNoD4xPRP
NPKj7ppOf6u6TtmTTAAN+Et9VC/a84oWYloKoDfmZmdX7SWU2Hi3gke2w58QiMY7D4cjOpoyinOZ
e97qCSAozvso+ZOYP3ozvFNSrri5UKPkvKuv0axUB6AQifqLVXkdGJjCmTiQ+gn/5RPJBgTMOL0e
EObfsOArIQcz8lnubso7vROV7n0i55qmupK4F/fwDmmJ56LNxs7+eQZOT4NzNSS3oILAqiLTRXf9
7MbQ438s49yA9BeP6GcKS42yw1R5VBQAPOpFCtDWpwZlyRzf4NJBIXsu2MVl9k6D5wATZnce6YjZ
EjX7AsBOG9bjs+3uh/raCFqgPS6KNScqAA1IqKxOrhaG4WZPIFYRZJ1A4MtyCmsjm6VqXV+7xgms
OrYxecF2YsPC9f4ZIoHNJ7hdNfJfo1/CpmFnvWd82kDHi0GkL5cW8YyERUoAeqZk8WnIYK9L1+51
m+5HsOQXtQaybofaWy1LCGs0AaF91J4J5q0wXTCUY2fh92tDr6O96yiLte+ziFgElG8FwcMCZxaK
ioLvMuvRMJjuj3uvM7jk8O9AX17LRWgOt2KSpmO11DIvXwvdahcppRBn4QjvAKn2TVuDy5O5IPJ1
Ukv7R3f8yqP39Gtjf3BD3e+YghkNSJnmxnJtxgVAnJRtBUtt3OAsLmr72dENZQeLDXT2UbDqXyW0
DPKwA/o5eCfSlQs43NEItt2AAYcsb0ZHseeWjSJNIPpXoz0xp5lQ+L0nfKrBu82KILup8SeCVc4p
NoStuh5kZaXqVrkmlXykhibZxJC+zMsl6fs4xHUaLdxn6oZFWOOr7oF+ioOckrZhiXL9d6IQik61
uspui+HQbJpVGSyjM8ZqtESug8VN1eXtpo+W2DQDsEci/kaESlyPoflUnVVMg+CwTVFGOks0mZPa
2eBeC3YSr3t1a8o104MN8Jlm5PtIegEnNlMW8F+vughyJi8aqClxoVhfqSAkEk0irOJZGp1tu0rP
FPBkIzmJ62Om05V4u+kGgtltO0WWoT4vGSyOoKWOmbYtKHXcSpBr8kZx1nRLQfi5Htk2L/+I8F7g
azwmn5G5SDFdIPsPmQzmtDVZK858aHHr8AVD3t9cxQjCP6ZjyNFueiKCqQxqOfhkR2gxHXd0yd2m
N1BMz1PZHEfCCwt9jInwOoEXHfCbQoZznBQ7PYgBskl9rbAWTHWQGxdMR4KXNG48BpOhOgUN2akK
5JI+Lv6nA15mgpoLgezy6H3saSFlIO8AIAOQMCJizgrLfQqlaZFrYIZTmw83lIeBGdegNnwIR8Ea
QHC3bRVmz8EZ872G5tBOdZq7ml1iAti9BQbYwbLFc+UDg8HluXkn9b9f2m8FKE9SGImvH4DsIomr
KhvTuTfBDl7DZVwPXcXp8Ny7ArjetjLLmXLX/FPwgG0cismZOU6sFNnpA5V1BuRE24NhdoIFt4ZK
cz9Tw2qlKKw4ffK74PRZtsbl74O4kp43Buu/AlB+ULhAeq9tu4Q3heHcNXytQQ3L0LvAK5931Ahe
66Zj4H7r/I4YThN9ZY6AfAWLvtH+CnkSGyHIIhfwPEWkLhxDpTk252WV5HsN0Ghx7UHVgK44ZIna
vXkKvDATahVlX99vJVS5AbEuMc+OuscLnGlcViZwbNM3Gt+L4Ss9bqIS4zLTQwQGAIh2Kd1jDwp7
m6qWNtES2XEtf94F9dplC2YNUXwbUm1nWA14nE+1+5ghjIyPVfSuCNb2SPAGYpGCLryDMDELll/D
dCyZFq0AqyPySOjX9MupxS0Mad74bubNu5gY5b5ZZoPYtILjoPiVda1ypp/PRWiKeQwxWBvc25Zj
U7h4fsnvyEk0ZObtG6dFe4tkGaihOfFqAZ0o8C7DV0AGONTFnUTo7MDUv7QPqbyEEtdk+zHUFper
HCZdNCINVSmWbAK2tiYkzmvJQKKCZ4ttpkADIWTAN/wMKBHIiO5rK3FGnfnZXsL9hxCnv6j80Qyh
IacNxwvnB2hp9CLUOKKLuiQhVEaflU3N3dMq0JvDy6tbtu4NWCn4H/8sFQZEUQVnojD3jPYkejm2
NwyzoQtuabRk4IxcfXqsTQA1Wx8hePApycwyqLSI/ffGNZ3EW0Vz0tvCFs+JeDznzFTd1pNxIltX
m2WBX2eETIXRcqHmraq6wkXxZv6wf0F+V/y8eI7NL/rg+5WY/LPpZkeJnWfoAFByCiuXpN/sedeP
fI6FFaOLktrKOcOaOF5OhPG2UKqMir5ZvBBhtZMYAL1/qP5yfvwbzfSKLidzsguLghiRAOjEv5RP
xFbyub4ZUUfZr0wUnS5RIMVsVdl6hnPeGMPypEi/k20kKHXwF1aFiHwvENICkS2YwYYYw9UxJ9hU
tZ9lvPuNILsI1UoqywPNNYXSvyzmaVCvlnW9ZK56Td74kLvAcwjcaarx6f/9jVKI1ExBrjaKxFrl
5w4GArK6w4frn81smiJ68HU85pgqn2+7gCywD3zifwHi9XXdQ9l0UlCLm1n8yRQaDa1E78kxC5vU
T7r3F7hrc60Hn1z6iouOYTAY4cDMeatmrXzjjNPCjAKFD0N5r929gQe+lYKXjBQ8zf1RaR8G+KCp
mNCqzNu9MjlGUvoAgenjRKXCBYZc4fx072xhJLx4Bqpow0MSOFJ1pRPZtdsgbprEEB704TZyYpbC
Bel1Z8a/49ExNxCpcCzEY/bxMef3guIQZ4T0ruzoIF/O7+lPpRPzoWOkn/wJb2/8JI7rYo5gK0VM
HyiDCTDOKeCQHamdTET4q8lFdJEMg4+haKd6lq0fifX/QxMM5R3QwFM1+ac7nEH8AodSC4MgsX1B
B1V8waAYUD9MzzRJaIko/WxNAUuu+vqfdNpIJc7MJo6dGKHzoOwr4XTQXuKYeQHDe5zHUHi64hnU
34dU8Xndg6tchMiMjCYaPwVnbSZ6QfwEPwvK9SM8zJrMaOgUrUgFY7vlc7p+ZmNHWWY6GRotckUC
Detw1kT3YSnRVdV5hIGufhVMIArlPpcI26B/ontVbvz+G68ct/ypeDoq6K/+iOnlHzUduImZqBnf
sSFPr71BAE7jUISUI2qOlxtauKTqDy/168wYy/Jjk394mPdBUTgx8m0sdoKPkNXo7n0VyyuG5hem
IRe5xFijEz07i2jvkJL2TdkUgIWHLTzCuyEnjzdi6wTm4sJ9PuL6xVszh047RS4VDloYYjq+b8+S
yTFlZBtP21VI2nUkwmSDXXKO9bbAPq9RF1GoaTUrYneZSzmxRE+chw9Rax5QwGADWQ11dLjMGQWg
En2RHHn439EZETjp2icqvVtW7RSTvkq7tigg7DF+1GGTPraNu6fauwnSLBloBlmSAMiw4xfeaHL8
JzHnGG35bVqoFANxcB2eiFfH5fLFGZmdSgh7kMFyPrRz/tb0zBAXoNTLFzH02jOaT5Ev8ja74p0n
MRQxMJVH7+d4IAUHgZy2PU7vr67TSbjK7YS7a/Z6u9ZCHv0p9rNo/mu/0Ehb5LG05t13PqUvEXVE
3oYrm+QW4RMveu7OTk54nvh+8u3R27mTcU6qniJsorOpRszSIyebaEej7Zggm32aO0TK1IuMY3vs
bNM5WK2MvB59hP1TwtOk41yRnkq/1nf2/hVtmCKMY5G7zrdrnRtKAK8m3G8HJyZVHcrftJUK0Ydu
9S8m9awmxm5C636GV+4mKTEORoZqaEt4BduxJuTjmPUecHG16s4XZj/S8pRC81xb03ffVy/9amrN
bvUJucJEDgSMXuaFElHaHHTSy8/GkEu/Z4fsxIjm+GE+aIs8MIFQQEfdeP3kI/XjsUR59qeCPvCP
hpDmSa3lOUBj24730azBPsBBWWXGNnRmWe3PVvvRTYl/Ks3OKlfg7wLC150oQqkvCbQD+oM0G21Q
rStDROShNO1JjKJ6yla+Rz8YWfMq36gRfo0KefXJT0mQUn5K0bSM0MYVpzufl3dsM6iAhDvhNvsn
cfW0EJRVvhOhj7eOZNuWlIz7yWRtSRC6NksJinjNT9QhHV5vnGJP6J4OlMWFT/R9DR+IC6fCl6pY
IiwzvyqBzLdVetbw8KqQ5bXgL/gWZio7CWFOuywzANuSDx+k6tmZvUB/J2mDB6bq+3D824S5vrLM
M9nPu5JJ9o4hWmnBIqWsONjr+TpaMTTu+Z9eHc1wNjMZQ0x3rSu7nVQnYJpmo9t1NM/1P2Pj08Zk
2+xQvLKmMoSBsNJHTZxy6J0HPQPKbtmAfMqi3ItUEGDUIBnoovsGXFm/bQM9NbgpAy6s/XuC1XoI
BAzY2krq3W5wJbwr3Rqe8T5FXHa9ZKfoStYIkM/gXIB7YH0YG74011sJsii1NQPW0C8cWyYtFw9v
j/XdrvokcVrvic3R4P5YCWI9WGD95q7DN4kXnkCAE5NfMlenFr8LcAnrRQXdc41sjHz4qkE6aC9K
1MxLfIzhlivOA+OpxKokbyhGobMCe57DzP0Rp5kIGHGsWHsqh3ZV93fqLNpgfGNosKe8dgu4UZk6
V8FFlIqva8Twtuh5FAI9BOsKBzhgoxraWJ3mrw18iLhWifhRWCbXf6h6PsG2YvAU9fkSUO0rCxxd
BeZ/BdrTcQTE+p+lE9kzUSekTeY/BhV+a7wlLzZDRPbLKERqnsBn82VJWWgSH9/AeMgwZ9FOUfYR
SOgM3XgLY7LgxGRrFu8musDaEj8A1/OS5EkQEabBs0ed8bA+3c8nPrCaEjQNQCZWOM+j2C7Ijcc4
Y1bVIhTNfzjIHpEzuaiyZ6AMEMjptE1a3/6OoK8oAzn5vtObSia7m705Mksix1bV6C9ezndQXCZ/
iG9vatJeDSGPNrsWf2wFMWq/WA1+puihl0usVCkw7qu76Wn9eaES9wlfLPIhudxL4ZclVDOoZIFV
liR1emZRTdH5c98gb6CZ5f26Xo2CVAw3jwaYhXTgR1hEsEaabmSH7wIbFWCOrN2rCIrNgulwSh4G
yrKcWF3DZ48BSCkHrT9hLvPjgsDJMUNu2Ddl3ZoV43qlGIqyspyaDe+ZyTgRIRSfFoKtqGVSyb2k
HSqGj2XHP5KOKJ904n9BXngNCXLpunhFwZ62d2sR4Oadq2d4B3GplC/EXYQfeIYhQxs3zspsq4R7
js0cGih+BJyXkGD+eFK7BFK0y6Ue8nW0sErEmxq2+W/bA0R4xhQqPtIFLWIhXsKJTklAHJsVOYuo
6jCaASIc8ekzzmMAwbLZiFG9+fZWArDIZmsCiBgU1cFxycEYyxCsVFXYVQOV0j0mEBGtqCJ+DJNG
0wegwjE6tMwRbLJXEHnw5QwvC2W2RbC8cSzmuvOVDhkuTjB6NqyvYOWK2Ufx9GUAi4qleM+iu5Kf
o4IHqRUuL4StjOHnHzBkuYxhaHINNiD6JwLA4wRsX9D4FDAeIlF50A3sv9uAu1CTLsTZ3pheRGCI
GDtDJLKoMs1a4r5PSfO3DODF+nYqj5+kdWiK2c5givTQJYHUct9KwxCfcEymZxJHQkdsIuuXz78o
GvQRSvM+VKr6goFhuP6yGie1caJt+TRJiuptX35B1fk9S8oqwS/JkDFNMAT0y28B8x9r8t4heIjA
tke3DeFMo07mI6Wj8nCTR64DyWluzFCjNZZ2fOaMgIS90h7vYTuMFhKZ3l1nugxl0I90ifgOH5hN
nB0B84lRMJ9NZRIGpb75dfgiKzAIIM95SsptL3Mt2RtkAYUPQR1FHWMWC8wMOomopB3l+Tsup3Ba
BUPsBQ7sagD4aK8lAIUFZQDDP1dcBNMrycx+mrCn7OnXPYwQ6N1bVyD/DQjJl2uqpFrSvPteL0bx
RJiSsVEjRscmtDjfKim2WEpwyui8vD7Bz1tjV2n8fmnGqCU2tcv0i3evZcnyiU5I/rZtoiMYb4Mp
fQhNiaDGhrOmHRkDcN3ZM/9HwSS0NGHHUAr/6DHVzdA+r9F+egBsY3OdCciQo8QKVLTovrc93+Qo
Cyf+9L1ZBZO+89o+f+PmxFRVOUs0TUZz1giKEVgARUR3u5DDPi0lNaXuhtgJoUcmAQb1CX9OAmp8
8mANqVHfoygqnzEt1/k6S+JHA+yTQuHcpaWitpuhvREiDjerzXVx80PKuErc6MZAOwVNt2hYN6aL
aFIFzI/WVWq+T/ifvtldm5pYIc6/j5UZXYBJsTJroIRaPYeY2Ae4feH4HwyWak4yid1PQZotH0kH
wtK72YBJ/8Mov9B4JvcDvOoVdQVKjrP3zylYO6/TZJEskZiH2PtXIjAhAFTkW1W1AjwRcPGx80Sk
7hkukqDOCSGwUbhJ5QJIQmZVEzXuHkN9vKSwq6nj1KSGP7LmSn8HMAdddsevPJOnQ5wmqy9G7bsB
DeBVqJ8HLv1GmZ1SH0vwoohrBe/kJLwBLaTy7a1wfUE00VAwn16dW0MReRXroqJesSVr1QVc7KZC
0/JRiwhzEP+xGsAvOnREqEWxpXaw+dLE2vHUcnQ4G5xHX7JJDaCapSYbk/jwy7HC0YUo4mQCeGH7
U76/rnVhYE1E67LldkxL4STG89u2A0iKDZILsLxUSg2ktMma16A2c49Tcaqr+rr6CLZnzuOBG+CR
nF/1WwtTWb6xr0vMTCglfBa6TQkPMNt6wHWEbk5YAJ7DYvVniE/+D9/BDcwdJJ8sf4ZoucwE81hC
dYwzvAOYwaydY6ShwK7OhA/FXtmIdlItV3iunvodf1rTCaoIjFdAL22HQRcjgM9jxDRKA/3elLA4
jZ+v3ANJfihS38pyUPYe06rtlu2igV9rr80TD3FKN93l3XjwJfvl8V1fHMZU8MPfmRiDG310XlKs
ygzAqr9lv80QFeqtSPMW000dVyJZN1GsrMsZj8AG5oEgWpsb46a7GduYHobFhCunGnR20foKeOyN
a+Eg1GHmBON6mhHCLasRFR6V9HG/Riw8zX+CJmT3fhne6hVu/Zp0/4B7/IEygMuXzYXy0U/Ac9rd
wJ+/WPY5rRTgKxDvL74YKej7mM1fUzN/e4/+YS9cdzGwpOj9NjgnDt4AGOIx9dcUm1GeHzgaVuf3
HX6rF5L82kSfHZ9BrEJl690BEdJD7YLYZ7y3ZEEfyxaEBE9uzGaNF1Zxjm3I2qqwh+btqK+9H2DV
TL3qTvxdZa68f0EBhUALwyr8CImL7Zz1m0oPRJQXcbLLhL4J25APQIaiD8MvS8GZj+FamSZtQIb0
4akkki6azrnI3Tf50tuXfZVWlKFKVGaHB/tx58nSR9BzsgT8stqDeXGC1oKo3UnTa6nrvRLzs5OZ
a6/zumX4XmYfsIDJRaapHkukscQsOSFVWJuSbgbuQjrUTXQ0G9KzKTcIlx1znN+TUIZ6ZVj39hO5
3WY/QO7g3CzrKKRP9LIPVQzgUoBbgXKfhCHfHus2kvTSCFeqsNJzleGbc5GN2Idco7LWjLwUy0Zf
DNt3Hx7g5PWJrXYzhga1booAqwd8khBphpph/lbIvUd/ZPDSu6TwD+LeKmxBMAo1RKsQbAa2KM8Y
vc/Q8AgaZqxTkO4wRJoC0+yjoNF/e6DxSFunAtzvENep+pVjLvD4UPW3NEHwKBNHBops2tWLQ7e7
+n+uqLSNmYWqmxNQJCb2YXhcxUuW7RWjrwmejQXZ4kOlsBCL6ZfUWoGfU5/fkUCNHNO4l2AOBulv
Sf80SkQCaWPCJjGxAEdnw4YxdIxdKAOaLkCbfHKYS0PljZDjsjDDNevnY+kRU6hRjQlcB3EBEelz
UztUuUwTO05CuaeFdCm4iBoR4hWCZ5CBKuUAF1DrYet/lltiYH+fHV0lPhnkKpOJLNdLolAqi2tu
jVcJMGECYj3ysJiGeZyI5TQEFMepK8Lmr3/fRQp5qCoj6fcIzte5a/BzvyBnNGoj3P88bbIY5Nyt
kzYzGvg0QHrSEI1wtu8n3XfcuK1Q4X/9R+JaoZBhrSToW5OONGzGlXA4laD9ZXTH94rpgHGm/K/S
RqaIT7i01eifdtNr8WrAZI7Tf7di4OX16xG/y4gnoJrFo3BCzlpYCUr7lAS2cCnAenN3AuXyAIc8
+x586a67nr4RwnvbsnhRdhpbHFxkzgaJ3mTsjkLXwwOS2hqhIOwDP+AJ2M9Do1BSfCGFpZcR0P8W
VKVAaACGHZd/qCSsq3RvnkQMQl8pjHnnWcyfZ/x0yjxKvWfgBGxnco/e8U0G+F/NTLXXCtfGdQSJ
Hi8We30OMtWd/kd9G1H6xqB9TFal7/cFEzkQeg2wQE2skGRjUy9WthPCSZkzSGD1LcfoG0KJM6Im
IHeeidsKfBvb/mPfp+Ko2jmYmzCHeNw9zhJI5EsGsLEziYLs6P3WlOxmuvHle4RzFDTE2ZNLAqzw
dszHAVb+EJA/hcsaidu+gQlofhxWvIyCVhmCkS4vhSZCAjV15Pc3c8QdaIvqfuwAUk6qEmlX1i0y
QIsrn3ipbN+DqhQ514ogyB91veuS6/rBBWhPP4OWp2hBwRf7DoucVZvYM2CrD0Ydj/ud/9LviGHl
wnyAIWqRkiYRrpjKrUSmGErcYlFLrE3/TWIPgBWJ6paSR1DIkzUiRTgIagwwNqmdMBn4MfcY0Y2O
Ze57AdrYhkCXnT2LUl8FD+i6fCDtuCkpL9K9/MbJCVX12qLxejQm6uy2lh6/98Y68mIUy65qCe8c
nAegdTrL9LCIfFbC1kg9MZS5VnRXwpGyrYGdBgb/OKbZfghHsaRP28gJsmIoFGVmx8ob1Cqpfwim
zF9IlU1VqlI62uGYeqEUEjHhSu5C9pncqo9wRLJAx3fTfVSqMefaJ4cLJ0KFOaKnqyVXYrMYX0hb
e6H4o6VaRnW8ATCZGtr4Pg1Femf2ArIBetDTfC2HTGtnshfSVaDQhMeo3ByqQS6wA3NMnNiJ/vvd
zvCgJ4/sutNgUbMH0NvSgdw/f4KJwYZ4QwbRLd55jjBtVK6Io28B2CHRlkrSSrz+Yufq3AmQstCF
pMFqEzEbmeeip2hm4TbkyMlRRqU0dLB0M3Xb8y1pp9FkqFekOSkGJI9D3ZFh2ADfQE+rKCnWpn3Y
H4D3VctorwNjMU84dLaVGriEnuZ3QkhWAmCpXkdGIgq2IvMkcVgqZgI94fXyivlofH5Rv+AHjMPB
wfoW8AImHJojWq9pa4Fjx0zZQOcjOXSofLaFvbcueiNX1U96bJcAyiLKMEbLmqWk9xXayu+ynLsR
/y9JHeGlDHO7O+JnnvQrQ23ydPvc+haTzXyyVwaKr3Kw69+PeAKRNvnS7uhxALCP1Qtm+nZEDUUg
k2fjSOCtYX2/yYWs6rWtWkR/7dbyRi9kjF8cqbCpLgwtNG/JlZpX0haGZzS6tOHcThJ2K94Cslub
PlyhChWvvcei4ytzmT1/iqfdjm+Gn4EvbPCcKp8db58JL9iiAOCdb/05cxIKenXltk9VUHt2CX6Q
QoDhmLbEdXCZc6EjDJeB/AYiSi8tFHCVrwkBFKsctm2rGcxy2sAR3Ktqgz04vQXDNkXvjjyJoMZ2
zqzlfWQ4CsRWnJ2Y8ekIQQTPpHzm/f7pRIqH8gQBo8Ca6PYuCiMlwAZYpq+jn1HNS83lfeC1ylYj
OS2kRODcngIfNlvS620vSByeydoyp+nuZdgTfs6GYeCZ4w0e8aGmwvxvfA0yPtj+MuxEz7SW0CuU
YkgSH1zq5BQHNBRlhoX5fYX3DZ6lN/Mw9WAfTfXW+AlT1PXdtHOQX4XXDeXcXeRXaS3uM+A/2lQ7
+3qVy9k0mFX48NN0pGcHTb8rtE+3yjJYN7jaVrckFaFoYGMbUkbj2jG0HzO2thkhOki4W0/5bpSL
I22ZarykPGS9mwN0CpvK7Ra0UjUPKLd3/g7iFThDYfrGK3pgFgHW+MAPQ7HDrTjzmumObuC+rA5g
7S1q3LWHc1Mp5gp5KJUqsyPN0mNulwMsJ2gYYIw2tJ6Kgzu41FRJiO7odcdhn66EoggQvntkSsMD
m10lBGNRPGxT7ujs4DrI/Ctp1sDhgMAOj3iat2KPFUZBgPC/vUg7PXfvZkK5TWgTr4S0/zevXrbQ
CnxwlhftQAGdo1EehzU2vAovWiRGOGgz1v1Gyx0QBY3uCSWPcad8ARlArLT2FUQeastGfnOuVovy
O9/nGvpbr68NtS/d5hgJQKnoxx2WM836p8E16PLQNXRJYswidsoNzpbc8dmoEL+ZzL64V2kvuHRw
W3B7xgYxtC9/SxwNivxzUjFXwG6TiW6KLPDimOoJUbcBkmsxlqa6V7m0OJ/D3jwEYfNIWKDnZw42
GPV5UEEWkFiwCXWQAIEWwNwcGQ1/oMeopZMABpIuBllgyknfKA0XjoRnBADJyBP6gBBJQorzAssy
F2vECAOxn8cU9Erkvut8qdTzDIuHQxLWw+OzcCv+M4YCaf6bkiTm0BMUNblI1SBk5+dDp+pjBZAv
OqRD8eaznT/KfpRVbkHszp7wPmcY1NZ/dTcyZ3wNaCmDnIeCgJuq73SYOpfR0oej99lG2joB5EzX
BqmPNcc25QSdlJgjWMyi+emLi0C+EDwRUCA/zhscijyxFwjZnEWuaUYj/hvD7B6szZ32UyJnCsXd
oCnxMw5TgjEzjp+2viLOnoSk8HfxHXUgwhjDR3MDNbV4YVnE8Z4wSTZEjCNBQuG+7b3rdyV/6svi
SOI8MPHRFTjPrrcu0NQc5rnA9IzHh0+997wAXGXTDZnwdAFv51zMN9NHeqLqr8Sl2T9WzaiE732B
+fWe7A1BV0kOT5f9V9UMZorsDNp6feSRFg6WlR6LQZRHMBkTG0enXtDnrtLVLll3MInkXi0CWMHs
niOod06uHHCuhcCMWHT2I/uKUGUbaKjXqrRem3H0uinBuD9peHclilN1NwscmLYgRl0AGJifbHeR
AYg8RSb6d8Ios/7X33cMZ0ZOgTtpHwVQLGnvZg8rik1LW8q4ydKREOsfbuuoKeKxAJegngG4FgvI
DBelg+FDJLM/Rs5ix/LZpJAU77gtJHGeU2OwaHCkCSDvxixfsHkLIYZckxaWtxqviw6SWQm5Q/2y
ln3KWWg7y2V1TRQFXNSdSdMYEeC2Mp/oBBWie9QzQ7ZLmPPsAbigzSsEzZ3CxwKULDP5WRZ1u23s
fYa1WOfU6ryR1yYbnJF8fyWLi43QhT/tHVZ1T665oyIHFiQK09uTNiRh4eUkhT+jGr6GRt3JtK8o
7AefeKZDjDjGAp22v1X5uwbG4y6tsW0Tvw2yvlOvjHqJBCkI5ntJ6svZUyUS+30+qNprqT7VonvC
yDXQo9dBDMYG3wMt0ZcNiS+Z2XHuqf77loTP73jIy7Jr3rKsPktrdwcsoo9Wgmz9C/tAwfH0Am4C
6cOug2nox4AzaKmKao11Q4Wd+b3OBrSKSUk38rXAUjRMz3KmWiHIPA1zkFRNyaNyVV+WbiqQKpYL
nDxPw5iMYTWyTvs/kVdiTX7Y50p9aVu/JO6rprXt8O9Y5GH4NXlpXbxnlfsNmuSGUMxlkJKRxtQ9
FINrun6sPZ7bRmeQdZ6szuqulUWFl7zSELYPq4yYeJDjDtCb056M5ZiW+gX/b9HoFvmLRTrTYUai
Nc5haPm8iWZUeGu/CaGqYQH0ZCx9VGT2Kh4QWkr3+R2YeJB/qKdks3UHL+f/58JKY5IczP2RoMR9
cAH17c/SronNF52Sxa6N8qofBrnfC5o4zzQkGgYiUd/bShd2d/dVdbda+rx1bVTSz/jwYVuXgqX3
fzSv5qQ8yPiXoyjSpdaSWA6T461jE9WS5OtkIjsKywLrGRj4qerJG4AGTix1GOOQ8TJ6paci0rH9
l2DcpIge7Q1kMD3krQyt1BMKzUwUHRj9fuDJ0tSlCG/ynz93R2VwY142bvWteyOsb4hK6Tc9goMl
7Uq8ECYb0eekUlrHuMc6w4pihYhzl6RoeIAh/NrXLr5PHaTScnsiBmKGEuqlNvOUGRM1P9xIUCzv
ZaEtZM+qmLLby5tTHqzEFsGe9JvOttAbgCl6TrPkT9BSVg0TppJ8qYzSd9tJlkiBfhwFkIyeMpN5
Xcl5qKlU0M+cKydGuxMOLF0essBa8g0WIM2DhLeRDbA4Mc34RUkAuWjxoBayKc6UElZZCk1fYSXZ
iLUNNhZTtkNDAEWEDlUUA0D89RHm8v3Ys72QfsZ3YCDQCNoi+n06FlFpDKbhBnGAFtsOGo807sxx
jdl/Ud7sZ9ysvwsgPWVSaT7C+BPtqdrXVhkfAuLt7qmx/nqr3Q6fLRK7RqozOoWMnHi915XbSy2Q
xrXw6vNc5FZ8JSG2ZCsZK++oASUmtdbF1Y55pbXP98cIYKFprz+3NnV85QLc4qBOsB5oOJIK0NZ7
ET3MvXq3o3ulOBBmuoZQlJj+5ZRbwcPnJK1R2CItEREVifox2bBvihPFH7JbkTbNMdGpnfucEmGh
p+Jkhvhyivo1m/yXkPks3OUasyfKVlyWgBV/TAW68/oaJ2QxPqPGVDIK5WRUplps5KfawQ5PCOrj
cJule84z/f02ueL6M6yWyDXxPfF45eB7swI/SH9dUnRMcZNFzcMNagTLAjKprj+B9+feCKdU4pAE
IQN9+BfabZ9pZjUrwy5sxl1JbjU0fG6HVF6+PBjRq1G8Kn2rNsr8j850fqWG8KQU+CzXgiSl1diR
BW6Vhzm/LxUBvVivUKaDlD2N4bvSATQZNxW2LHjHULYGayV0ypIRp7f2chNbx6FVdP59yfynPbmA
d8aDFt8Luy2tdt98WtkvS7kmrrw41qA6c/TtaiIxtZ2QdAC2I7LlQWLLXN4BZMeXXPEzQ9GFRQE2
1Bb/3BkiNy1QZvO30Ffc45dRGnuX8qzcktNYsM3OCHy5yAiElRwbMNCUUoGasViVfubdoXT10/PE
uAH0hcrMRd+CMLmP4Hfz9eJpZjWS+SpO4yyFW4KjZYFa22aCaUFexXnsIFHJnARowJ3tho8075nw
2TBVzPDMZuEDpFCMFEx/R9me+jZiZLBn65nGnZPrK32+PQ8WpMrqXeSeEE1FqD+I/ORjQdkAx0Oj
jlr2owcuKkZUev97JQctCipwTRqVJohIUCkAYu2Mt7v8OYkP+5W5D9Egy5PuP8kYoc29ZxlX3/qw
WMZXZWxLOfl3QMRPmFBrlEcX6yn/+xwo+oE7SW76KNOgTqujJcdxMAnDFzJj6VwTw9KwFMAswHQb
v4PxpWarNowf41CSByWqDkH1XTLZ47z1mX/+gpHyBBbYE2Z6UhP7s0r9NONRZ+DDrXRQlodqx6Dg
hj81WDz4KryeREq81z+6J68YL6jcesWaE11JTgvzqcUv/iytimv1jHyXlHx7RB5kHOmUsQt6Qhnp
e5vP5USMzwi4xVKvfUeCv/yvp9EfIR7WA9doJvHWljvXdgPO5ChyBdjmVlXreFdqbnge3O4JdXxg
9hAUP3JivnrZK1oJbTY1rZ/TETZxRI6AZiYeZVGL5C0Q3uvm+CoalROO7yDbKMFCR+jgw6dr7eU+
mnKrvkruoMs0FBpw+K86APvAz3skiuOjI8OXuZTmPlZxD6d0Sot0keJA1JKVt7a2q3ootXU8vl5g
kwnAY2kPsi4X4VbPdhyYzvAkEj6GYfppQAs9wv58rHnBJqTyl54LqqqaFKyiEu0Kwet+HjHQKr4J
2M7zg3//H98XRGatP3MiS2tfug8b1Pa5qmlqqPRaRXUQXpY//3lwE+iZlPPZYDOHulKQPl8etZsm
A910CJBQ9sqaihKNAojXttHG/qnBy3/jxejxKwAV4scvzXV94tmqil/zqh+yScRH4mxBQo1aAkIr
bJq3uwTfOCnJhLDJqsEwaCuEI68tnlfEYrPPL9A65Gxqnq6bZKMFzko8QYmJGNqHeNd8CgfoH0B3
yz8KdFI0JMsozRUqFn5l3gakD3ASv7gffNIomhfqTEPVgL5OMz6uYMQsfZuLHV3Jx4dt57h++sZu
XaywemSjUGmXN7t3SR1IWEA7n8i9bvpUliOhSCKqdb1rLK/j3lBQAwCYSN8QzOW2h+zawKu6giTy
7rezY2DM9+MgNWZC+CNqMX1vZrPQ9r1f7KM4/7d/MZC8Rpt4AzW5MIOeIzQWmoKY7JiIGgmsvLFQ
L/yTi1snMnDni0ZquaaQsl+Kx1tQgrqTPXwKTQmCNitAhfwr4+yPPdkpp0Y+1lGbyQKWjBYG7xgA
6tURFZ8xcYpagxsqmJwrIjqbWZeNxsLufqzLgwxi7Dmdwnqu1i1PQiEenCapO2unMMXwV5HBruTd
FyVAmsZv0o0t5jGSjhPnCEhUr0h/IFciC5lXk3qMXWD12fsV29pK7osY4vqXMI2keVLJxIExYKSn
TFg3DFkCkpCGNumv+Z5Ikl4h2uwibYPhjOD6UhkdWDvL9YGw/fmEDasK3wNakG0fSXLKi3gSC9e/
nAqt/Almbz1Wc4gMqq70Ttw1x+KliXtBkgJk22xmoUzdxAEHGziMuRmfWgZcKSVGfEtp4CTzBcwd
DZYKeRbjsmXbGKtVYFIfrh337ZYGb0gqJ+iHvIOfRpFehme2mwF4q+IFL9lFGlzaZhk/EBDeOJxG
ZczyIKAZUVPYJz6j9UTwnR11uRPW8vTP3qAYmRsf1e3h5Xf4Mq/sBy0XAVbSpo/iHfpOEwfewBq7
8z/NPsY7a/nSwVy9zoX61cXwMrZxNhFZ9QEcLKjXT1R2dgS5L9TjVw9ChRv6L9Zw8++Fxv0KEvlr
jGt/v7JCTGEXkZo67fBzA8o4184+zTNOJItRJYPyAjMLShC5HWeCZrDvJj8mPMZ/vzaR8sbMc/7B
I4ZRN2JiqV8lH9WxT7PQ3rsPVItc9ZXfM5wsz+EGQ9JWiNTRCWY/MT/fd0WhYGp4PkUAVC2zlC0h
S3XkSTcDRMO0JTbwPMWJa45oTdeuYsS178dflqsANMlVc6d/Wk3i0WaV/rhojY5Ihf/pGAHEvKb6
Og7UzQSizNxp4K5cf/7cC3CZeTqrvBFOI0ygV5EkOboI3/kwqhaVe4XvZX5581YjsulVg2/a0Klw
0JlXtCUQC6eEfj42yyX+erV5Asr3g5m50jj9uu/wEfS/nxnCXNYDAfPZJ2g00NTiNrln4c+ZJ7Qp
udieq6G6c0pyqLwDJXOK1oM6u+5+5F/Qul6HREBZyI3jvGQ/8Dq92MeRE/TPzYpG/yq9+vxh/PB7
NbRqjI7XBGh4vjqGO9IzzKgGIrnuu26Wwsvrxqoh9ermSpT7qSqjHOrjsrRBwvDxWhiylGwW+xNj
xPnB+J3VVV7axECVhfiqoLf5roWOgBwxuJo4z4awMq2tEZnWIId3LT43Gn2DZRrD5nx/3hcl97bD
7fiTRNczexZt6fpp9kMfWmlQXGAM3mGzZvOqHMxf/zQyNlnHPegXHtHEzqht3XGIkrsPQgIdiWLg
qyYqbsCSao48yH40W/JyPkE60Y7I6ELQ/ILFwKS9TKUqeiNeqwAfsLowAMBxlWJBDrR926MER5HM
AFEUHBGRM4JQa+541W0DRQmNuqURASIsRkn8OKCmNlG4Ymlwl6iI5u0PZpRftft2YVE/iiI7QogL
ZCa+ymcvnSh5EHJyx9uqIWAZ5FjJsYnKMSjDJhbvHzJv0/tvaiCK8A8VOnP5QdbIsffmdLnUbs4L
mJbt7Ud9EcUrOZ/TQRVjvIJnjDJtayZHmXgMVhIpFmDzHYTQBz+qAdNoX1T0O0RPPDBw97O7Vc45
RANQKLM8Rkv2a1XGwNnveS/ZURxH91OKjDYcCUOeG7aF+1EDEl/9klWVFy6pqJLkXwHaNtX61LwL
UKffsHVogBbzXS8fznbVGZKymaHlyxNtXhhdbrzul8M0R7dahL62ymJZuXDTu7xn1aIkyaClBFaJ
A/PmiD0BDPuvFdX2M5be9qffgjLBWpN0KleFROxNBa9u2NvTrgL7jjZc7dgravBaA2Okg2z9MahT
/1w/5I5dHyPM5tEwHA2nKdMZN/fbrU7d/b7h8CR/ObbZ0K2mEtb+w04JBc69eB6Myoc+s0b7THK/
guTK5BSeqtuLmRwNAQVI/xralcZBCkw3IWLnGxm0q0HONYnPA54fBQYZtsmGe9eHz2rg3RZC5mzK
gIWadVlwyvYxbv4kDCYd/M3cTiFkoijnNjet9WDUxADdQNQY7fIWmTO8KEKPgKnxUfyu7FWpM0CJ
eBiLgcqmpnBExk5X5FQ1xs/yhHvqB6QORD9W97UAvmxp8Ws93SV1PXo7CF0yNoIq3Knm+ErW2s4E
01ynCIwbbKqe2kfdGoyRZqBxVqIwer/VlWdYaT8BkoSFkKtimOeA9HMzy7ZXreOnWrjZPbHGBXNN
rNMH0zdsSPN2+KcDrybv0ZHJ1REuTqP9r81Pb4xoBzefDl87fm1YHVmZh4rxusYnVPjMwcQiD/ye
uRkv/GXOpbXQ4gl1gI46T/fxHylHAguUOoDkYR7I+Ka4mGpzJKLqG+NdHP1CY/Ylxo4FpMYgAL3C
Lj5OAyTvxFTldqI43k238WMcJpAlXLrzvD+73f9oq1vNk22CZVh5FPScJVHSP9kFqaXGrqcU+XGJ
8rOCaOQ5tDShHISzUN2IuoKdjUpRwpJEd/53LoIJ9FntxOYgxh1+ZjtUiiQqOKKQ3wOvB8iYCAtw
rqmc8G5WTuDH8KgzPxM6HuwJYjhwD4hvPaIsoE8GmokMqr47et8m8pqss7LF5jVMNOpV3GCwG25V
UzjjCa7JErpm7gpwzVU0D4sRyjg4GNH2KW0aBJBGvgvx3SP7kKU5o6Dn9lFS6OKzxG43c6z8d2Ux
L+R+tvi5WuWE7uuBqnvazKHI1m6jmZlWq/3iTHMN1AecL/fzuVPwz2zi+VYbDYGNWwPFRttjPoZK
qvHAll+I9hq/aRYo5hEz+6SAE7lgXtZgP0JYju1mc64F7a3i/D2LaoB2uLjsfiMA0jcApCJAsq+b
1JGeHi3ZJ67C3TkQqhI3f1GZGjwdx3bdw3VDYiRyArNSZUoyr/oh4nxqGH7fLMYultX2l68dHzhy
S3gYrwh6uPAtA5i7WypeFC2ccc6fQ5kF/9l9voxE5JWeo2goM07HTkqaoP7HUg9dajj3vmgBuR4l
UnG9xIyceKYbdS7stnWGANVBAf/h48NuhODx3E6PmB9ygry8fJUGERierJbHbF7f45NYBKuNwGMu
Jy1AhUgJazcisSuOU7AKl2gYfW37tlWGAqaBTkWl2n8pbkbuxavw5B7YEgzVNOlzO79OOZyRsXqH
FchSbbcf5sgPfyuCtmZ6UykeHZP6u58VVzvQgbTnibQGsVOuf0guLr4qDliambqm/08Fiellt8Np
M+vPuCaJXJtTdAr48aCuLklJ8ag2jXgGMrq3QEN2cx9RchOm3MjEGwBo8EhOFf1U6VJ29YP5LU98
ars/jqejvOLROQq9cduUyfmStbWySzjtXbhUCtdzQZsmXY3ZGKOmHPWjGfxD86MUJsX+7ylsYXfL
Q+Op0mr6mx6BfiWpgfdDhoGMtb5mXSHKxN+PDPNSByIZf78JK7ZFADRG9QHxEXiokJgJXj1+fzMQ
dHWi8QYKkYFDHZrMkgUnv9ymmaMcRZIE8zkmyA5uoCkbP9G3hmFM+AHrkO1rgImJy573Y/2SLfui
+vJcBJUo4zufmDoV44bPM+qsKvNZiS3auzc6dlrhB+aCaK7R6+WgNwGkWG5BAd8bhxWsuC/ELjbC
pjsp584ifFX0GYeVc+4yHS0tjCkIqLs+C6PBqc9KtnoOYkB5x5IFz7Emj9jd0uuMrA+8URJEait8
ww0SC+8S+Gq5t12/iJFi+Pg5wg6jUeRL0EsEHr+rlVqf93Cz4laGRIkNoZavTbQwsdNlHwAgHUbq
IWmwohy7sbfNkBudyDjM7yFrLLy5VLTsIi0J+Mbmnr6BqgJuqGnorsdkRYr/r3nBX41KNf4gVpSm
ShIuIVTk0sxKTQqpHXugPRkCoqZDke8R1BenKMG6+0FjFznBPSmDMxULdJhPRo5+q6Hsl2eDlZi3
MwD03a0EL0jMdpjLqwq++LukWldxq2MYDfC7V4cWPYZJq6hACZRRUIQbH0+GsfHrq3L0ibVaTFN8
RD9TjBqh2bnCO0lGmAIAT+90BFhfHFzEj2ukla1ceRcj5/aTlwi4gW8PPxLawMvGl9CaD69WVnWR
67hSNwBnnGlkUkWSx1YuXnHAgGJA9KQ5fZdR8VOxC5UNUBIu3FuojE6T9gOjsvtASA2G9eHmc2Go
3tA6AiDMVVJFjosmP1GYZ/hy+cHMLMBR4lkEqwI8SD54BXo8m6Ckd7V+uczH49cNGQSk7ONLk1xC
v2qqjrzACU8ayAlu4C2PHcCGeAOOgu0rvi4W4zzhTT1rpXdtobznZvC/wFfG7sY99V6WKun6HJWZ
liNCwayM1BivWHE/7F+kmwmKgh7TnrEkeFQrSAaf375vZZgaTYKhvPB1X3rdTvM4/B76+DZw0xa+
hftUy7r4wWuONSuPiI+08SEsiselrVgryRk7tXrscn6Jg/YnZF2ktFhLZ9mf59Nz9v3wwRZfDYup
ERPOm5ioiOZVB4QwM1RRGwvIXANBjSEYdaS3UI/3myv3OdCYCyDjcfXu4l0lE18p0sr2n3fVFyEi
B7DGNQPOlH9Bmgsw8ixp7lmmI0kLQ5VcseuE+leGnM/OM/2zWzexFPUa/OMS++hr0fBeYId06fob
5+BuxJ6PyLbzcWgb3JcIol2aeupA9Z/hICNs58Uz5FSYjEmBq2Kzmgz3ijc/g3odERkdoPHtQg7x
3lr0nwN8sSj8yeQrR5YYwb8doANzZmJeTjXulBlBVA5v2t2aUtWhjyw5MvdEpTNDrrppW9fybDsy
yZ4tAf0VROOTBzSYUJpJHLBmJkR3Oj+6jpRlbHOHYJ+dCWjWhnR0fpp8ewOKR+y+DJgbW9z8EesF
A0DBsgIsTBCQJuX8ZdWoIIN8GyvoqjRfGaYtlV5G/V4vPDAfCvBe/h95SDcRRu2XbGgKyM2BrH0s
AoVcNhERoAIEnyzR9vk/ttZneRbb8rcpCCEhKmvqRoX58mLOm0Esng4L1hwJD+af4UxQUyVX55Rj
dlFy9CXHmHPVQgkUBnUft62plPNXlyiEp+SA4wfCAi3fNaNu0zCfU+6TDNgABv6xY/Lc+GVb+6DB
q9GhrjG87x/D92SDk7TieIH/HXXuzwB4IAEJ1p1CcgGLIB/0cRgnak/AC16mWnC91Zc3PtRUja2c
OaKWyqUuWWZdxUwRC+4I9guAkK8vU6oLZOaHyH+wJ/8lypFA1G86aym082r/COXbUDESe+Jlg0jX
tdLJ6OIU0omM4tmYhk1IKp0Ux8gGkJgRTGQypyQuV42rUdhD9d4f6nkRFmtKuXv3lppIb99JUjkc
djgbdH5gHOPTF/3RV1FNNm1ZQWbJBaJnGUXry9/9mH61/yV6jL1l9VLZG01ZuJHX35fDasaS0kxR
fYhoV5f+zoOiih9ZFt8OcYp6XFmg3PRQTXPeyE3BJ7ZymluweKWnpeobh9RAdxjhD1bkc5KIPB1n
Uw/pS8zaFQEk5y8ZH5PHIejkNMO4PoG95hmYpqJf16gqWtyGVnoXTP08hdD1vvxOGMHqjCZ1jxMq
jZZ1NMWEHGs85MM8FuFDRULnZGM3f5HGm+fVRWSJu7irpi0igtBiUAeeUwwjglPTmLnz3VernPUA
RgZv2VliZDtn8yVunU91/k4pujGlG8Ahangs8ZtIWooYL3JlYhpkrGA6H2zZI32IcJV07ZzgY01C
CVC4hqmt9zt+OrXQUIdkCYl69JRbNJkBDcsIj0ZVDNR4cVV/Lxw0yghB+H+zEEWFeIY3Xt237GVf
KnLJY5AMUuKzNYqu6hoRm1n5IK4ABH6S8MoMgW+uFe/qRsODkiwcymL0bS3ZuccuR1M9TyGZ2Rge
cYqCpJOQwlb11Hj3yhLfgKrq3tXtc21ruqHS+eJ5/qulHtLUZ1ibMroYNpKe09TUdTxyZc7mtrdU
8/tL3xtLZiYSIvvGFnfc7Aauu3fH9Zvqv+hGUNA+sVeAjjZ+hCLVFaaeViqkQh7ch3CzruAMYAi7
2uGFCV1L+QNQyRLA1BLVBczjTykRo+9ENKJb/wFZidXsG78xf9f8AjG0eNH9016d7EiIMer7IrrL
E11WVnI3Wy6e2TfTs6xdnVDXbGVG6k6wROMcSNDNLLG4uB1MovLXCKuBDG0jfrZiIKhj6qKnE+Nd
X2wB1V/T1Sso3NmCTQRPAKJ8q+BW78Uk+C7ZLdahbZPncfAAcB1Kzn3D3a2mU/Itvra2W18/MIgB
AJOCJ3V4QbnBSrjFWC3sLOfC3aV9QXSRt4xSh++KCmOH6lLJCBbz0CXytyrOmkRohoWNv1mHS+aN
93V0iv7dFfvHdXr9yuIKT9Y6sK5dJ/omAAyzwSkygq6DrWbJRT9dS3LuxSzyYrnGqSHClujRReKM
gY5cdUl/MdYGF5pNHJg79UsQx5kYFY1JPa3PUEfg3emNQFlaCGu3g3ANTiV4O+XlHfpTGS3KicAH
OayMK353y7GJC2JG1sI99MIZVprhemh1UTkbh92hLnKKVwM+im0P9DOSsHYBqpQHFNCA+vcWOetE
r9Papla4EoqZy3iNtNFzzRLEBjtJvj+YPsfH4d7Qe3noH63FrFbJe3DfMcDr5SGZ7b54mwjuEybt
ATvPScnkh4X25nIzqUVxzOxzJSwB8z97IhuXDSaHIYIMioZmmCt3WAtrGArT6C62mVufmkQzNWZp
vV2q2H9pdPOc6U+bcSTj8FpfXzSSXqse+7q6dsR4dPHiDMOjSB3IfQaUhXAVvMye//n3XBxDqGrz
BCaY+Q+TXdLqYGd8ePxgpAc4b2TzNB05qAwTdTiNU5aw+nNhd4u+Gef44nSr16HqPEthcJTRSuTq
ceYNr2ZW/BN/ajGXXxMK6HiWHFAsHFMB3ll6+JYxXOdVoMcaJJH6OvEY1TbI4oBTaLVsBVdEJSvt
jI4MWZ3I0GGmjQxKtSAZV5RGeTRktBe1r8oA7ymuAGZC1p+2bnFJDKlLEpdrsVZMCwCnLtPRXMvE
JC7JeoNGJo3YYB9q0Oaw8aPfslFLf3dazVrBL4NiEAeBaX3RXcrGc05z07FS70aOS++EEF3Xr73M
D+bGDCmhVXlNwSlvg6WodeVYLm85jGwKLlxcyaMSWLCKy/FnWNFw4wRD37me1qL00s5k39OWRBUU
3Z+acB7i7B6ym9nsN1/agdFWLM5p81+Qu9lAYEI4kWFjCK+KFVuw2wVAjZpVCrHYO2HfRUCoaAOP
Zmo6sHvLd+PYyhDFu3VgPzMYRlAgT13z9NsPk8w8N3yUSmBiEKPhcWGTnd6xM++o/1cwJ1yNdbQq
9Ix0f83L7JltOCA8FV0EsANhIRzBrbWXmIEpuF/SViKEOXU9uH5gUjWwFn1gsr5K3T7Ver9bsIs1
Vm4X4YaT0qce/8Yoh4esTtPEHV65YPuultlwi/rFDby0ejDJvxjDqcBQxOURUEPR3hAlWHCZ1U6q
mleBFyPZO97FgWhC0FIbFG96eFd0Gkl4a0fkO/dugGAKo0GRwET8y7JwSVMmr02gxd/YO6E4RKuy
2CXgu7B6T9wEHyyMb8h2KWoLWn4jb80OP3trel8nhNIdElz4pBaOjk6wwyZDmOEvivLxQoPur8BH
Guq00TSyUZ5ofqFqv0Td2KTq4DFjQYlVn6tKCG16DLHBixhTHaUwLe13OJ5RtBKTXii+JUGVVN33
GTumdtmaqh8V3qz2qmyZh9f48WB4ryCAFxcMAytd+xlH/I1BBqA+2b3rCi+zog9ZXsIX5JEjGfKq
ubhXIGtIxKOMYIIUqZIKIdlHsZsSJjCCcwQpgUD/9eyhOJX1i/xflztX6NKqI0++XSgOaB30NCoK
gadQJbrfRPeLHV9197XO4yjgOrbGaJ2DZ7PEmq0pQpO9PMgieJzRoldxl5swqJL+WixtGjypkX73
VwXwh8YWfNSPohgKfUkzs7CNpQ8SKCnsQ0v1Uw8pJiCgYCxfcwnX5VlLk2tsBJiRZycHjgwiHYwl
/i+zVpz4JgDT76o60hWd/0hn3YenX/WpHt0xQnaTgyCLR6KLfdkxlyRsRhbP7+wVQ6pfMohUjgiX
I6bahrE1isxHw2Nny2FVF4hzhrTp5HBvmF9Kl4ld59MO/1ZuttQIfrQp9pnCLZK3iVKEbcdiI/1S
jhJ5OfXUhrSGRqzQKNfWnrUviqr2RA2ESC1E3BzP4eqh4Dpkkaop/0OQH4qfUvUDWdTAAIeVV37T
TFnf4RyUNq30pllpJHY2E59uj/yRyQ5RIjNB4U0IESiP0+MA7VcG7DOlkauGVdXyw0WDfnkvrz1M
d4Q2I5OedFBX1xHEDdz/8OYqZxZuD+xen2qv29ixHvczvlXkcWmu8Z7YjvTtEVHqSN+jxNgxPTfF
v6cqQ/iRxb3biMWDxXslXYkqfmKuMI1TQSabsjaVHxs/IHUzWmSQu8xfezcHhqelW5pwDjbdHbpq
h8/NkjPllswHTNrRl4OWkH5ytJSwpQb/Hdt6cj5iJlvGfR6dG/UcHUBy74bNZ+ponT8GanLUohBb
bqBCVFFh/snbP/XqM4drD+sZrYGFU6utDUdbfjPrarILwpO6WfRR1w1078Kdva6sKFfwkRCjBGXw
gdh1fEjkNbba/rSH+WhXF3or1vWY11/mSL5o2LBFEylw3B1udFeQpcqZ5fnYO4wTaNX/k8NAb4Zl
BRzEw4pokJ8oQFpMqthpfqqkDYmLtUnfSyy6Hd7QV6LRllpk22WWqclLquua7eZGh9TVZkvjMrbr
5OG1j3k9qTjuwuSMCJeu2LnwWbumt4qfCSHO9KhU3ch4M+Z8pthfmSVi23uHC/jYnlI2OUDP0Vzk
Ia6nrJbjZP8tJHAxYkD0+49bvLbVcz0He5zaLopcYfWA14OW6HVsBkCEy5JEBy6Ru9nzNafwYY+2
KsQ1JWEdcetu8Ny/reFyMNb+WoHrdDlnM0ZZNtwh2wAD+ss3H6yUAc8w+kcpgqfpQ4ZsWH/8w6of
NyV2D3TDeF2He4aThN/WyURS1xcCrtKyh+6DLAEEkZtwoK0IdF5gqIGaCMrXZNfsBBRERdrcqhSj
J+f7zrEDMQ4zGRCKJ+QoTQ8oI3U3KR+ll2zhZ6RYK2lioFQeRS6tdtNCAYSn+/Qg+KTkqNz6STrn
grjQzj2XnSfMNCCp1SPg3BLOZ6EaSZWHuvHvXVYXsScjbFPVM+0kOMW7friuti+GLRoljUezSRPL
W2JLcv1iWToOue7ww+3wn67VChzVy6mIC7YWzJVqMurnt2D+Hp3aJVteplm8E2MxxwP4BZwSrsYN
Bxe4mTQXR4U1V2wVAYiDJ+M3c3FnLUgtc7kHTQ8qBncaovHEKgkGwJCSVxL/FO/T4sVdNf4uDM5/
CueCLJLsq8GNmnRCH5uN+LXh8Vn167lvXMnwOES8CakLDBtGa4N5B3C+HJxJci+O+CYNB7VJtEV2
SYf18SrmtWqC5cRDTd+jBRrMKOZt3hNYCUUCaQDJKvicTHOYi3C1GlcjQEaZCoDQi8PVZeKeFME7
LXq9fYX4NjhDVFAtrG/bfzjh4HANmArNrf7iSP72PdyzDA7PIbOCOL0yHNS/+FaVeVvmi2SSetr9
Nkl3HhJ84iJxvxJ9jRKUVX4sPwPmzeZ224vRgraseOxizQjsQj+oKFhh8x6ftRqI0ypS9OoJB1cp
ckmYIpYlrW/tUPlR6Ioe96qc6r4X0D7nJFP6Veb3grerl7RmmjuqUqLrqE6iYjonX0DCYfanQ43M
SpqncEt15Kxh+nwyv7O4pBZ62w/3Zu7odDswfoEZZvXb4T8b3jiUptC3zzPTlCbUj0vlSh35kIOt
URoDe0Vl/BT2z3B1Pr1iqKrGUPaFuxY2EBBIOdn4AheSCp9Su8D6fKpdTvr7WkXhCVi7mGxyA8AJ
G5H3bHmK2MEKV7sEGpZB/PcYT68NBs3VkBdMY7p+FfRRbfrpgYYaJIps1dvyBsPgDtE3h3VUpawL
v+byhgwTokiQ5oEt0detFHYQ4hc50N0NM94O94WwwXWrMhsXPpYAwVvvfw6qoAGuOe/K/k2zmjj4
jOJtei7EgKYh9EHuqt9jcGvl6KxnOoNhHOPxbu9f2MDhH/sBpfjxlKQ20awztBh4BPRZuioFZiSD
hpXRzhFCRcBdQGPukLDLZ6SKlaSDk5rScKbyB21oU/GfyJptY6DJoF1veS/FSVg4Y6d8Dgc/mRY7
FiHpqQVsFwYUigwr/iK+S26b4D45x27O43T/J2dSrLIrq/BeNkb5yt4cbCeLT7RjrqhYD+TAqOcJ
hedF1O1w9i21gXWQ25JUMgqMNfV2mBEsFozXdY8LL33ivPWwnKWOPlwgXeTmfKxxGrm5L0+WTcuc
xQUKFsg3plnkAZE1Cvgmm3Ccu8Ba9WrDPRUq/hHYnxHDTxR8B3AsPhG2Gtbh5Xhsx0hv5vuuPr+M
wby/oO9h/btGpoaeXSEOj+J/j1Bf10cxe1u7LnK8G4x8nCRChnUzx/k/S/oTJUmQkkavUCCERRbT
x8vWwXYGHH8hEmKQWBkEQCpxI2ZYhewF3Y9MtV0m1TSYWncUJ/mwoNAbl2UCwZf9M5XE8+nbmZap
LU0JRcRxC1S5D+u58LJSxjxaaVVTAdB3QnzNNg1MrstroRdCegX34fiNN9bYoX1KKSXABAGhDEBo
3i2XvoyaN791ZT8UR791fWQdoU7HKJpRkV/0e24ajl802ZJFqo/2P/y2VoU9+dU74J5DKaLKPnA4
8Er9lHf7T1/cU4ps5OL3//5cr0RtTsWW83dQDWja4avaHj4rc3tFKgQ4PQosMm0yxZPwmqTnJTm8
x1G9L2+Vn05i29LxGcCl/Xk/TZv8ESgpVzjkArwJiWFTUVSQhPZiNOPTmDJNP6D++Q2bBt2epfOE
rs5Lpqjq+y+saKtgE1Em6dUO0Y7rzRZbDo1yebTXLO33RDKPDI3nQ24o8ioRWQvgrSlo1ewOXy1t
HLa98C+jGL/aey1THEdqs2h4UpTcsZIAip8K56xo6KSekmHiNjqSkpX85s8RYl3IyuWVRBGvzlcg
24q231w/NpZMRkY/xkO9Z7n+uJxemuPFJ8c/YSfvVQ9DEKYD8FtyMr1olFAm6ve3i+2YSKDLtYsa
QUeTcwGyW9rc7b5KE9T5oSJPBGT574vU6Di+tjuTgGZpIW8V9S7eFgZAQXenQdqBoAhCb4o/I88B
7tDssvX368qO9JaJIPgvyi/ZmJLCdnhZWwhBztgcg1n6ClJ8ygs5cAiOzTdJuDVH/7HYZcnzWf+Y
M+Gx39XaRq0kUOAgvIUFfFV2i44i2W+W0owkw+obzdS/his/zjk7O/yBg9PaabHUZM3QKs7Ua9kc
BfvqSMY5e8/gNdYIBGgRQGt7q1Bn9BKgkDEmxAmzDUoTJvkPB6U/PB1s58Z9jJLg2rPiGaR2BUAp
qrVH3bqrJnci+G6mjlsMrWUL2bSJRJcjjQpV5a2mCDw18xlwlEbm7+gC9TneQyhKp92c/lc+eP3A
KsJH4a9uTrNp0CmngbnTbPUP91oJYvn9XP36XV1nBN/mjfxFx1xQW/L9MhvGKdphDoR6AlmHMI1D
5pSAmLM/R/GTBZgWRZPO578xa6yyVhLBy5aiuJ4WIdEqTKQb9nZnJypeT0Beca147Qo7aZnfGQgu
nOP9076ocJEllRJUBXerZvUvlXzrcqjBYLpqAmYgvZLDJCcMJFvGEEG8vYeFEZuUYoKJhWwMrwQJ
YMPWcvtYKyRNDy2oWm28cdFzK8m9ZLs4agGnkZDtFLoRJ2K8PpcKFmNdMJ8g/ZhqwMxPwX/NjbSL
/urDpqzppXgvLgV9vasK1Ht80vpzH29bxSISudY14ufarqibEuCtn3ekXTYzcRLwQwOgy+Vsnpqj
e7sw1erXNQZesWxkNJMYpvEjNLu+KHRQIZgFfMb1+h8yY/U9JqxVPljzepxFc8pPdDK+3PaYu8ZL
eltpn0Za/r8lRlqaLuW79Zmgl0nt2zUaDMEdOslPM3EpYVDj8IpLq98FfL4hrZ9UIUKPqlR4Ipjb
UnvKkj/MAB268MqjghDJAZ416yEll37KuilTES9vd87OwvIMhcaIl1sP9UVtJZ3pA/JHw9II9WaA
wzm7e+ovFLOkTtFLjebz6U4OBhzY45fP2/7D1+kZ9Qnd2xorYuuUYSK0DctsyU6vDOxQ2gL8WdI0
0YM/OJNaFk/Oe0bmrt9xYnSjwPmOEvw0mmfY7POgKJh3I4DopzYW5iFZ/fewTmtUw+et39QCg0hr
UX7nMrzAWp2UnsFH8AhcWx4ocDr0O+c7zRgfTNRXyx+sQC8s46nSvXdVJiLaveOTrsW3KJGuXqOx
cMTZjwizu3ueljl4SM4PNgP9YJk8J6V7CcdvjpJSH6lmppAX4iR7ZkfTXlmdHuWjQOvSayNYapc4
lSBou+xxP2ct5oLdGAABKZH4eKhyZ7sj4l2am4KPR6TCGEyDg8ax60oW+8dR8JUFf+FtLcPbyPTg
dnYsPWoC8ZEos5D6+LafdWwTw2jsjl5eFuPYIoZvshkUE8Av9PxaNWFdYaxN+gqtiYiIpDPJsniI
6NaUXQLUdrOrNbKSX9avvjs1ZKC/AY5jx1ZDwY7oN6RKDQJIzNuxzEFiF9929apC9+dXVlktc0bZ
fP5IZ6UqTeu49ehM0eszLMJirLghiVOhOeJ4zFIy7ONG09oZ4dyZ2A5uaP9v2kCDSfqnV93xis6C
o0gzvvrKzxCzTF/3scacIJvbXDhvYfH5SexHB7U7BSvE6nmpWR8RpKf2SWb4MzATXlV6oa1vSbqI
G6YVJhUKqEOQPC0xzenBPnRJoC/VBTGb89G4V+Drn16POaAiEoo4ZaabPgXTn0QASlYyauG8dFmH
hQ6SqvULyvQs/YSwbyWL9Fpap+CH/K5zUfBu5RKZVFwfc138LuWGXfRR7m2hsSDCFhyGrfpjgMsO
s0dE6hGu+AiAX08PPQDM33ok2HiGbr+XE8AEtlYeKkGC15+uKsHPTTJ6HX7WQvpt76/W2QDHNWij
UoGmmkMuIgFQGwmfr6fdgcc1eNrvm8HtXdeSL4CFQOKeXJZabjf7p/abTo+ZY3JxYhcs1bmuxGku
4wMI0tcDPgCjqZz0tz2uJAD/rb+M9+mVfbaIuW2hhUIEoK7/XQEOldWjUZKIt7cV5HxHWz3otTu5
sCN4+9kAp/AIdW5wP2abXESxYf6AHo/pHS9xWafQg7YKOIJdKHsb7cp4X07M68x9BHmFrPWUEsGS
7q+r9iPv11zlRC1IKvTOQKmpoGroC5wXJ+CY7fahkQ9FciLUMHqEAypiWyGNQd/ZomIs3gtr6m0U
0ly36LdGycNyNNfcHlR8UqpWmIB3SenLK53AyvzVjjDv1XFJex8MDooMiSLIACMjoPjkn6mfIOAT
gEtAejyO2m+Gr6uTPnThp8zrNtZJfBhb8Xwys/HjT1HqUbQYx8N/2+h+fkw0iwXHSceYCIza4aHk
vqbv/5onwl3vs3LXekIHPDVPopsQwxo7l3u9ASVXbdh4lU2jq4qNm6TRsJo+R936rRwo0pwh9yu4
PCs9CZOu0oP3OYi3DmZ9/QsG+sJRFRPv1RGdNlDJ9edDTtqUf2dRjnEmff6V8DIJBnfx63iN7HlE
pCWFbrAUbhTrAo7yoNwbhPVJ8X7CbsW6A9i1f2StmIgTjZi4Sflx2Fymd44QE4cu3ipn1D9chN11
I53JWjmcG+WVVLHMU3DXO+orYoPUfbBQQc+kn/45wZz55DYbejV3V9PbD4BlEdhIpGmLZvORjok9
WgOcS4marL270Hw9naQVwAQF5pPWXkns2kknAe9rnCEjb/c2hkdRuF66BvdJi85xV89p8Mvh3Xkw
17IQaYNfSqkataCQ4538aCkBnOHC1PA9JD5NONQOYsb3aSUkVJubs6VrJIG/dWGQrxDmOPYE0hEA
tNzpshSpuBPJgyNnOEnZuwSlkoXEzd5FNE4jpDGViaHnO2DiPfQq4gLnjECkLwZtF2U/BnLXNiaw
4TAVmgNOxO1IF4e/I6VTEob19rZILWss1uwLce1MQ3lLayZK81yVDt0P/rOOs022HUyrsIDR5XlP
TsaJZ3HjRruMh4/1YRSWRUwfEV+E3QNy24y9rz7PBl+DZ4A5MacIqpvpPiTlSV+9XzT2icHpjgLH
PzCJk0FEWAOvB/kVDggEeMQBJL9X8qYYeaUH33uXenPI9yzkJzyXZ1s19JHaOMB3bNTvImv3C+kV
oRJJ75wROk3Tp+a5Yl2kAeyS07qbOaUrkCElp6O+zB8Y73sz4qwuVvW9JPi82j2Q/FMC/RFqOcDf
yfvH0gYzzFuQI0+LP8NmLd73uQe/y+HNWWE9OkbOzQJUqq//xh1MLwoz6tCuG60X9Ah/pBaG8iKg
XcyRsiwOuAlnLFhSUGeWYu0bw9Axz3G5zeEc7jwYCw95EAr4Oso/ONdeQ6qb/HJR/TlGZWTPJuEW
EUDQbV/7zgpECOa6HL+cbM0lt3xEVeynmCB9AR0nY8/2BrtkDW5+3y2N/0aDEWsN8uivPl+PH86M
+wObguzWlkuZsOdVwzoq8yKE0iikFEGbX4q/+3lQzYMA6bOmgUGVhyng7pkPB+RysYPXXlVX2EsV
NgEJ+1ABCyllGqjP/5dGQ4Tcq3ioP7NZ64osXJK7/8BatYAOTGIAD2kY9ewX64LKXisuMpexbLpB
v/j8Zq8Vw7tvVQLGgcC2tpXSXWNr2gdwRNZi2Kc0et7wuHFHJ1mPAeZtzBakFkJeWsOZGPXcA3dm
1iX5EzTC4ZYgNEqJUKvGjSVA3KUi3g8FnO3f9qpakBjTwVFMwZXjk83i4CBu6oKJFdDGAHivf63/
Z5j5z3TIoVNImsBLnEpnNTfiQIhX2o8tXeGZMc2xId3iMrTit6L0Pj3wibaE7dgaXgesTApTMyz+
whXFf8tKg5kpOhkxhPi6EaCPW0PVpewD0XK6+fnIj9Ko46IKUKHlb3U8P9sW4dVK7H7sGzc+OQw1
doRuH/h8WTUzjq4fKH28lu6etYiZUZA/k78Ovk9yrobUerjwXML+K6lUpGNvSgfDH9NdYeYCRJBv
VeCQq/cDzb53Dn5N81BYmfJCkCSJQa/IYvfgDkCPECqtqv1fdsD4h6Ba7bQMdzDfVDV+hwvWW8/i
dv2A8xTP8yghV5xp0eaGyGavWOSXjwiq31uP+P+2WoA0zJAGXykZCDH4t/SQjJvjldzZGZsTwW27
TiUTM9F5ESfoSKnZYUMjcA2cj9fDhaN9H/2w0l6OOzkl3b1MfjHE3Yy4W14+yS8uSK38ziBM6m/X
cLZgXfTRUFHtPSgD8mu0CDB5f2JJ9UG8t3mPOR/ylz+c9UTzWDoibC8psXZuB3aoQt1gKFz/Z9/T
j7n17w5Hrr4zH+fEGdBJ758arBzYnr/YlrC1D8bfwBIc+9NFsw3a/vpj2qfL3PgsGU5Le1HTXuK1
L3OetDjG/CV0qoVUUa4KPBPL6YYAJsXfvKkAWZhZr2vFALqS/est5u7oOhv6bWJSZk04yFD3WQD3
RqqlSW9dge/EF1myF5e8Roa7uiWn2hOCnKzgWuaEjzIxt9UKIbSx769Z9TNvQfKD6noR+HgH4WX8
+NooRIsQeRDZegaDL5zrQy6LRwW0d46YEYBFHQyMjh/9Zb5nfwdrgRwZDyGVTetz+OS/UHyX5LXN
OfWBfuTtkGlkn1Z+ca4ZUMvV0KN9qwQcVQ/51AobcMMzdAN+NMEgYGzp1eAJtjxHZ1Ee/FUy8yCq
s0jbf+GKw+hb6ntm7B4hRWmV1L+0H2O9kVxcLMK5gPHFT6VR+/42mN3e3G6MXmXpxihiDQMAX/D6
lJWDz441WWYOOdc5vT8hk3otz1H5jDN7oJchMlKhdLWAMBFdDh/0CBF+3/7qYHWoy7xj86Ee5u+N
VytMpPkl2R1SRXJMg37DvM8nn8QuaIfAN+Ldl7vnw0h5c8I2TNnGNoAYjVt51yis+xLTjxyY7B49
Lj5ARqRI8Hhiiwmytv9TQy5cQXscShAdXXCI3xSjoRMU/ARA2SDvYdHlaDOTFGGVzPIw4J/TerEm
JEZ2tAaI4oO2Shyfc4l8RaFXnREyY3k5tGT2vEqeSqtp+GmebMJBpCPwY9qjKSjiIVYA18uF2zox
kyqco7sCBawyjfZAWrerIwMkw6CbtBRO43m0+DIhDzQL68ES3Q5RYtJqUZvIA/FsY1CGBKQltcwd
lh4wI8G/OrtkiTRq3ctRT1k3KuU2+lhcSzll/R0vTSE2uW/nTwo72tOKFGeTDJjgxAsoNurDlUoe
9tP7Gr0rfgpelELFBCooAaWEq55ivrratnSH64CELbG98Bk1770r7kdoigkgVh/CEo0xdHRxkMGS
Iz4WXY5yiiZOFzUrR2b4J8RsjO/jh+h+ZLZxsTh8zt0vwx4PLeZL8T17HsbHqN+DKSSaZF56Kp7K
v+xtIpwOGi/eZvaSdBAV7X00xykLXt7xG9BfIp7lb5VmhK0eHz4jwjINd2GHeKkepEP6DtJFscPo
v82Z/1IYMlI/B5HVgT2mrZap7AD3tv3TSHAWMBf7mzFdKbXX0p/bhFBSLtRED8xkwfBsywU+Su4M
as3EUFSXkm3Ue0lxt+UYYYlxkCgMKM4RFHn6p4wY9nKxYvDHmHGIY9CpyLFm5KwjaCYcIH4WxgmV
2nDvcz5iIyR1IsQZ6vRbM2b3q6J67FbYpa804zuLJVv3dKAgAPV6P6wYtyQA/8qE59p5eraGh2jI
1CY2ipjk6M4hARxg3XbV28D5G1N8/WU8DRDTDBh+AXjxtbWUT+ZvfOONafmF0kAx+v95auIsk9UF
rypD/pvKCQdlCJ7Vd/ijU8JK4dtL8GU1wTYK4+xYfcY7TZBPlXXr8i62xZ4D4mQ1ecJmqea06fPM
RHRdhuZ2Qtc4CU+JGNB06x+VFFZ8Dn8yitX+xZooso8C1wEt50VGq5vNsZirDdkjw6DsZw4SV2Vn
zek+ilYYnSA9us0q0QhkC324+RGIsi41Qv7hBS1i8KGIND+SF+5U9jECeux2loSic0jOUYKsTdVi
1r1mFr/awLFvgSG18FQx6mIwJEb8nf0EcM8pM+PlXXjWoTSY3vjwgKKMwZFQ4yJR/0Tl5s4fkUAr
/TeLQJflJjEZTxJUdtCNbtqxXSHQpcDHorKHQWhjGoMPECMoHiSgJ+3tD73MK4dKgS7M9zNsNFd3
E1l6wrqfV9H/LF5tQuPBtq0WE/nCQqbu+lHHW2PWdr7nxq/OcFMj6djYwcWOyW99bxcxj61zlk0/
o3CeoyhzuGYQCirN25N8bC6+PG3uG8uheND/CDsyrciAt95rOIgXvmkSfRgueLPnUzbW7S8H+YgA
ThtPiMrodnFwgdsohPHx7DCQEhNpbyzpXbXeH5ZYKwIXUwdqqle7IHgU5NVzAHYrekdeTbGYlKNY
BSTrWnZxXlvv+3OOzwNWgK81JmEqemzQ21zbtbw2uqp/JagP7oYdUgs4Y0BSAA15bMvSuu6mTJf1
vy54GtfolDwh/OJhwdlNUDTJKeOkT0KTFFm/aynMXgdafOknmofad5yO09ie1m2OR0SXgZdM+8eR
ogwVFWmPotUsrVYx+Q290fcBYL+OjxdEW+W8kw9grhsewVmqW8qWMlo9vsQoHrkxVUdJQJH20yFx
dX/0Q0DPexVb1qvKO+n0M2puxl522tbijiDr18uOP07kZJ+cUd5K3rT0uG8bTs8VNS6+tt9do0vO
wJ0BcEgH3mhj0vXfAQAxb/04TM4sqA7zJl9PcSzSZDdv00eE82mCZD+3dioq67xeBYwGZagAg8+d
dAeczGDccoMtB9FyjBBDeftHXScSblYYbjXkqxrvQmmaI180uhfWDdhsLPlqKGDBptatqZTX9Oy1
PirRAGDa+ZTK5MMgXHNCXSEpHhW57uGvNtPxniZp/BreEmTxWjgWSxEE15bnRjf8od1DZDh2TogS
SC/7qsXV2Low81dm1E46a0oft6AJm+F4zmtQgupTMHbkIkDhG0CAxKsEnY3oQvXTjmKC4TTKFGGQ
UwaW+qT/D5XYu0PdXL6vlK1tYhAwQ1qVgpz0DMaCjU/HB6a725zPDAg+6P1dIlSnbTi5xVyvIWft
nmUfyteOOUkg7wZRB9zakGsb3XOR7PKxVVYjaaQ0Muomm80+b0lghsn97mzJJtIahD4dotq+7M8P
mzX8l7aKQD1lnFwhKbFNVuCu4TVEzF3WG0b+PgwAs8ebW7Ox144z2r8yRNvgRiz/6qTxL+poXTVJ
+6gpsvhW4dWvVtL5LXxbbHXIUjZh+rOH59LabUN8GeJOfzV5Zuo54bnGDQIcBDmu6kkWLt5djTnd
GEbxxUyeZ6DaRPDjN9jB0yv06j8/paQNJo8GeidDTPQI8Ex+GQL2+/MhEn/rJBqoxqeAdmXqEKsk
BZsFLEzHKSAkRXZozaRhEvmJvb9d0FzK59v74QCUGe3MTclXTeyqxpiwGJXUNAgQIstzhgQorC+g
MQiSWEcjqFcTqDxruuq6PBNxEk/hS+YYncTYFijkruct457rD9v8xteJDH20vYKubbvOUN1pBfZB
MT4s0s9Z5+967xj5tQOLQ9Q4M9HO88Dsw4+hLdQ07BYmIvHOPOKcEJQ2K/M5fs0/9fiepilKfU1q
WeG1IGut3cgmEsfx/tlLufR0r0L1ksUrpZ0sbWWAsp2yq3NanQZeWvQrXPSpWK5h2K8kK3PQT5OC
+itZ96VVzzFgaAPeEkY/ZxOxWdvx0MYAbUYde2uzWMug+MCnTEI5lTka0rToaTfBGPpPAx2PTYPl
BTKcj3z3kNJlRvn9wmGxuROO0nyDsxR5H7/mqhVwqO2B0g/YHwFQlwyfPam9qOKGZHl410MAHDBG
Ca9q4OZfKpd0h+gqcMfFYWsbKZcwz+q/4NX629ITTsSiJTjdMOgDRnJvIZyNI5jQ5IRLZpPOun1Z
AM5kqf05FCNoPrNmD2dodHnzrKHY2rXebgmHN5SrmgL1E7VrU/SQWRbcbT9ChvogIwK96bUT9cO1
ks9Q7xl/2NUHtG5NYitZg6SXko1nNhmigOSmabg2aN2EF/HQUIgmIYAHdYDkCl3RL4oUoHJ/AoYf
wi4FCqj4hkqlaJj4TI+0YmMriuWJ+4QMaPFh8K6Ukp4ZlC4cbWa+29NGxQ/Nn287ImDIm01EVlx0
tuI4mZp1tVIAJ3UZpjoQlJpc3ZEN25HCQEzuQkwKEVUEEB/DH+VOnAcx318iRwmmOzQXjGHI9dIp
LDO3Ys/HV6jpYiJSH4eZSjlmk1nb8nGDx1KU1omQQsh922pAUmGZDBippbSpJq/jqfH09NNTtDVx
Q7nJ9RcLljTrRjbOBGfGyPlmO9sOgIoanbTqIZ9aq2hJnqV0zyDk1WSc2UePHgAAA1gk/hp7JnJJ
I1kbvJQy2z9pzGI4z5B27BUFEDofLsiH44j0xsHZLHPbHDlnp7A2EOXpAemTvMglBiTmDJkDwNo4
QL8XkYeCjWRbXrvX5HylSmJQ2TabsZ+jXqXg5QAIcH3m7awH8fAEe7d/Kq8zyEPAf0Y0lm1zuMv9
eMwzbtbYGrD9d0hdPsC3IODF2ZAf8IbkvjeYmS1xvLGXxr2ekOVLKx7VVS5FwMr39F4M28B6JEOO
G1DlFnW+uKhJ/SUz6CR5VjFVoDctAynNerKvIuOeqcO5t3OyM1WOiM5UYMXz2qK+tBUk8rHJxMMK
Mvfo5mXQ3fTZtblMPLwz/MhnutLj6VAdDQYdHXqSJgSq6/205eKy4OPDHP3802pZXiYZ/fdcYp1Z
bMfdepGGg6zrJ5p1JcQ/LQT3tULtmKY6fDqa3wLQj0ipdtoYne3HLMfLvYv2x6FkqPkEYlCkDU71
Bpm/IAzaOmEYhXqdpgPZ95HPjR/XGV6/OuUyE7pAWktbYTicWwjMUVyKh2aOZU09FI8UbFaaeJ/E
wWUOuvLQ18wzfAiziKlA3OSB9j52l/WUihtLdE859njf85nzur8djhtJGAbKU+c1KzhbpTvdmsXg
t57/d6ExVLT/QrMo3CCjsGwAkvBpqA5KD4YZtdigGuBgmplX3ksHN7djU3Qp6e/7DHqTN+tKZM/l
EkcmqWfQGdnj6OVWlA6/iXi6GMM8FT+ZB0UJraiU42emLMrtkNT2t4S2AY4sgMeTF0nHQsT/z8tV
Vg8/fn7iMFjzBY3j19BrqxZLB5LGExhwoUDm8dmnJ4qKDmJEl6q0767aFWvAdqWrp0rsLrBNqD0Z
DsICWELgpAoQSTST1ILthmfViJjLKkSGsdYI0WHtziDSDdoQ8ywDTnmRpgnLgDr5g+YvZ/8+aw4b
VVSvbq9W+Z54SRSMxbz9Pevulx5O06IraM7iiQsWBDqVuoZhdjqbudusZboDAct/CXRn3Snpaefr
UdnF7eGnAW4XVC7ImPgE0aexmEb2h03nN6YiBO8Tx3u2l8sA+2vJseFMg1ThKMHI0qRYcf+qkheE
dAQQlhclr2EISHgFpJRDTEwFMxDIOWb/vk6FVOUyZKNYNPByvW5PLb4AnF3OhQVq4bztLQh72kxV
8/T8rnXPk/WGbkboJ4kXZmheHA9s0vWnTc0EtZ9F75KP325pAZNfe8EUlQ//AdI34owlZr7Nba4t
pXIpc4n2dLrNlw+vw++Emk4S9Dr+3XZ0GllhAhAsVkM6APLvLj1px7FAwW36iIqlAfHfoO4jEVBl
iRArpzZjysf79Lg4OLDeDt4pnV0vvMQuYMzmDV08pzKyXv6QLduk7a2YMfVsUeiJsrfKBxfnnCwQ
iDatBctIV2bps+OoVbf1YOIv/pRV06uBfg8W4uSj1mzHygr+b7uyOvyvZ8KrLQl5E/iNZH3FvxzJ
by2oza6bwvXKAgIR1HpX6MOBxNg+AY6pcDMowu0fbMLcXQx50TyVw/Dj408ShQhfdh1zqklAXWbP
4pWMJLsLlsPYZoS0tlgh7HtT9wkMvUO8zMGm3v0IcIQ7wzNCjJyP3PRLb6yMzV85nw4+50IaVOJT
SiMQBOesnMVEP7vTxPk0F5/A8GgTg8xeSvI+8CAh3hWqXgLP8rNVmVn2bZY7c8Bc35S8pGq2GVhb
ljF+QRc1a6xHmi/BrQVSRLU/7pj1NfWjXGzTK2oL5YsF9OCpX+jZGKLpN0N3fjuL5Y6dMssFSTeU
F5SzA52mJfE69leTVQS2lH55pKT4e+yCAR4W3FA4caWUT9Dx6xu7A27V7UhzkvJfQhSFTiIhKAJw
dB37J0qe9exXk336nhzIWb7LRIRwFAmgCeELudmTShJr4l9HUnmqgefdwYOGiz+7gk2BcDwhTquU
5xZhBeEz+fMSPzTG18hKwbvXmsry+YiCU2GnyWCaShMb7ndRJCL2eEU9TPCT8etmbWzdWwGEvQxR
3QBmjXD4MMhzIjTwHLIZTVgtQx0zOJWYCjjvnY2UkUeFLwZDVmN/ZyGYMvY8y8EcEjEQ5nAP4a+n
jsnO+SNys9Qp8TTYw3202yyyQtzfT4bbNlLJ7Fh1ArC12gdnpPEP53TOn3mniawunnejJqsGXALl
NEJoQjY/MeSVRTC7WvHxSaC/S7TWHqegnG+Z3u8Ap6MMLypTcd+VW49jdumzwxDdDGjs3mXgeH9D
xC7CCFO0Vblvs9kLZy1g1MRnpxpDRRpS5quCp6AH2z6x4v+Gxx5ePWSk0tuGEDqW/L4BDmZLeVNE
QZMSISZNTqxVjixWMVEM/HVMPON7Ilo0H/7xy/CjwhzrncxNd5e4CSdPiiHm9ntfw7YBwuGMHa2K
EtvasRVmL232kdijHDFLaWXplWT2Ok8xk8IR+E6p2MaR6gfn/UvEHU2gQqMbMEitenbHM3coQYIK
zqWJ24KLN9r/SJ6zFX9RL0K2TfuyM4LtAkN/SpjN69+0WmjqAh0beTdkQuW4Q6ryVHeYQqA7LMGy
ICg9AmNgAA+bQgaPJqXj78E/UgrsBanup/POlEKcc8KO8WbEqlLVoiz4uzAlZfBxFKy/WEI5hsTz
syEUEZS4jPHbmcBnJ68vCM4lygYm9niE+1XPO8Ugv6DxdPzzRniIK/oNmT6YXTgFJo3fOuuHmkQN
pr0uCjNTkP6i+xoH+GqofoaO03X1LGGzE9Lwx3y0pFrv0s3WeRQZ83O7AmpXF7A+CXlVGdknCf8F
18NJmj1SXKrJfUMuk+CVRKAozlYz4O0ZspnD6NJzGe4RqPfz06PRNjqkVnw+RZItivndgpjOCdRo
7AF3GDYSO4cLeEPGyhuHwROpYAQeFuzilwE8Sqz27jvd58cNz4Z5QIcABNSvtg4d1/RG5JgXSFG7
D2oxrPjGlh33g8rNE4w29FUqhc0Tvlxx5fACJHaBy7NtAgcss5KFoiSrhLYlugFwi8miwhnGO7rk
WKLvstifLN0ZQ5kfqVl8hyVsBmL0JgnkBqREqY75L1V9dqKjRDGYX/MxqD3zJKVuf1ronlGw8HLy
3gbhu78w1wM5ObLBb2ijaGJiFDaFtDuCYMZthqSzQwGFhDzBg8/0YNhJdLMScNM0pYCgHu9mnjJM
ek8BmSC5MESlWtI2t4kqVUpxrI+CIaO8YNBRamduTH+0tguYkcoTv19MmaqyVSjeuuDNXVpG8lc4
lyAUKuG08GW1Ka9Yt9LtrzKId+78Z+TKjDdEO9bNZ5tfXh8QGuMX+0qygZyJrZBOblW5JnJ7REkF
WUDZ+VMprwxLy/6Ekb/1dboPJKW3R1eFW179A0oalEwmszw7u5CcYCEtCID8LpoUTCy/0lA60u3D
heFZGy2vXxRbliwjKt8MMI+7SM0l6XVcCKya6kiFSV0fuRhdy/f54ljTp8lbyk1PbTMM5sOUJSJ7
cwazVk4gT12kQzqzC/6c9s5+YFM729vFQQdZOpGlYshNvnCsjMDFmTjpNPSCcTbyiQP72siJfyGG
wT5M76x8VYELVaRAT6I2TY1qFVsUxp5BhYmp/9W83RnudxH9+iqyKUD/y3hBNI5t1hE78W9C75l5
DT2hW9UzLXMiBRhf7SAsZqjb42zsxWluewn44POffTAiAERAu6xV1CElnwdPqEZISDyGnljgnbId
TSAfst/KvVHWIVrz79uusKV3VW7+SexMBvszagOBC74dMUevcE5ha+jJBCiyT6eBVwlQBe+TakfH
CtwyQMRY/3RHoVYsFxiauarcH9B3K6wHNrhWbq29gFgqGx/sPciYCz3XtBpI9RwDJt6oqZbNgU9w
gD5bzVVQINVXAQyGl7NXeZw69KMOZWFiFWFnaeXgwPBfRgk0BPr86oR6irgyhtgzChThrtSEawmS
G/+1Lz4Kj+6jR29FSidfKoQrhZFDXbzFBTo+CZg8AUhDnFWLDATd3e4QRcaPB/Y0l+hhVD+lvils
GYNq3cF6h1r3ekSQROhoqHtSY3HAYow0NSDPOLQ93svQzzw1Gur0PvRafzC6EA4SFNbki2SD3fnx
SxKz+t/5ukIut8JcfGsKVnZ9iP31sCjn3JPRenRnGrbrv9o0kF+FXs+Ecl7ngK8bv9h/p8trnBQt
/N39iLCGoOyd8EocbG+H6mq6vgI1sMsH0l/hYIm1kwYsYrKET0M/V3kf+12bsvfebPKCKXhle+Iz
4AlMm6kmSb8LOdnvwREwwKy5MNS9Uyy/RWaw9h8mVrtHPuW9upPx+S2H9mjW7MgegchJKSTnr+ta
/cPAMhJWbfeuscapyKx9YiE+qHn//f6PDEqGQx7MeXlwlZ3xszfPWsEHK32uUSYkzhK6BlolO6TA
Fl7Cdf7Wwsd72yXTvcEQxKtRyRStPcHRpIRTT9QH4SoUyti98BU5vJ5HcN2BTMpkRxsA1udbgShG
xjGn1BlhOSYHlmNQu1U4SRS9YuBrk2Ad95SgPqFuymcnMqWeIGD+9tHxcvNFJKVyeo/VQ2nbiUQR
cNEQonrcgQ9CDsL6meBMYHzOruQNFVLHWLJ5eVjF+vpsWqYF0vJsmoWhcBmeGrWgrogOp+Q+CEDu
cOv4hAR4LlFUeKDXLVKaFGgZ5JBMJ6XjEV5W/wK4a010bB9JhpZD89/Lc0zHEqUwgfNakTEu7+rj
ryV7vJA/3Yvsn+7SByfGiPhw4v25E90fCHSma3W7SYaiSpRbXf7gtwLjeBnU76nkscsbgEyQUyvS
rXPUL7LqInSIJxcSRXRMcMah0RRZK+KXFO+14F3AWnoa7ix56yyQffbZleR0scEZ8Dy+aSJx6kxA
ophwim4vjcBSAX/3mq+NSgxBlUW/MIOOiZGmxN4mP45x34dnsGE2OW6IVziyy6v6h2fbZYExRnwj
g6CXAeLa7mvlpybIbFig87A5bGLN+RqiuDM5QNWC3gYzh8IYHsD9VKHTp3xi33AFtIKzfSv4w0JA
M43revwwt9ATmG+POwwslw2GNVnXmEfSTZgNpePXso5mXFEUAaf5/86XYwGMzsfOSWRJLDP0TKFk
806het1WBBn+/DVOL0X1Yqy/y9q6cbW1CT7COX+iSO0bKFCHydGurgfEDZ5MitE+JbctvxMzaBr0
Nts3cQzRrPiY0TS4hWg4AEN6wRlzf/1XZi0VQcQlnA3q2JTzEompcgIfy9u/I22FEf+WV0c5+Dur
UBHWsNd91skTs83th5UAn4G9TZp4feo+Z1tZYPrXyYXFqk2S5M7Mai/50ifQbDrTEZUjJYCVpF96
eTc6AV/G7IQyTN4r0pLK0pDEiXw4yu0JF/EjFcVsnjfIR/PJB8+p+/dwKpPmIg/Uaob4uRoiPOvm
A44Zda+2Qg5hGNCQk4qvkVBiUEgr5H6os5+HKERypDELUOVaIyjmYiYat6RsWrnPxZYbfTKHoQ79
n0s2/TiN/+KXwb97sw9vpoArOvH6hmzAwxofeP12EFnAoUE/siRM+yy4iwG7tP7P0lMUm2lnFsdo
snVwtaGepyo+v9fhUukEOaVl08fGZI9+dLs506QE88+jD/pGx2SAd0zUxSg+fYRxy8KyXgTdzZuw
4+f4O76pzr4nTn7YLIcbrFfHD3iM9tQC2NGoDvlFJmcygsIj7BQvUAgIerzJRwRE+4VFxHU08SRz
dl3rYZ71E87gBYM7jGCdgEMN1GHFo8/NpjYxqaSoiok09/ChGFYBcKxmlcFtQ8JgZmqvzxYbNytW
QOXs5W5ZWyREJg1o/cKbIaDCuM7Lw73DPnRB1bCIJTpJ8qz8n2YVQq0Fy9Ytu8D+RY1YSv+3EVGk
MiUrDy2PwvCeHF2RFx1K1GJu7reDEtgGFBoccp4juDXBTldNt+wkLNA7WNU+e/yAk9DXNB5czyt1
lrfZQWfqhlsWClq2B3y6kAFDG9u6i2PUPBj9d7pxyciUluQiJ0PP+BU6LSYYh6USXa73MQMuHp5t
MSVU9uUcLnTQQ8TWV8wTFC3MDkl9AzHAhNavG88l+JAHg91PiaKSwSt/DSkCIwvU8qeiC1ZCyIm2
CFp5r6E0m3C0jymdkuGEbDlasSbeFeF1cuj/jnY8zb+pn5RV3NHP8LGEaYkkQ0StRKB87VjtO9+M
t3opcQv8bPfyurPUdmABjKxorNoXPNV0QtqZjG4uCKu3TahSTtStr7wZUB/TlfvlzZxaAhBI2D5H
Hm1RXio8YvRPhmwXGNJXnYevb7C1OPRb/RokRTQQUINWQE2/7mae0cPUyQHYq8sYAhH9RmevGA4Y
y9NTn4RUfAH6XRWmv3S4LK/8uY2vHSulJjGgMdfx4E47fPo+aOja2VhyWkfIxHsx5wByotJtBbML
sZxDj32aeZrL3NbAu2ewhe7jiSmZ2snp5EhDZi6rdTshqFNmnlg+4oM7qIEVIe7X4SApnj2j17gS
DzSUwxintY2gpzE3MSBmMt3ya5sJx6LAsYuzx7yXlBaq2eC0JcKVJDU4YpHUIPctvlEaQAj2bMxG
0w2VPnNzcvQAo1urCJjSe0XKLn2/GxAD1FADYN/eTP00QoymgVYOz/Qxj348YEJFO8MykyguofX7
Fv59Cr7uGAqsFM9EYGKnErfJ3DanKEIbbZkkbxjsbEiEaBypAOFkcsNL1nKLj9Ua7OAL6xzxNCtV
fjdzc8n1qtF7ETro6Neu/8yAtWHNsvY0iYNyNnVBSRh2RoAeAjhgzJrqwWbGKOjiLWuDz09LSBSg
Z9bN72KYlfw6Ii5jdjjWcvson6/05G7/Tc1aJsLmSqFVSNZ5XVFVB5p9RBpNN61YWsv6K+vS0fzf
yysrK55ShVuEJ3tl52WQECEqtNRH8IqR9UZNHMsDf4KDyH06UKMMOUXn1YttMGlAQsQejO+Vno3X
kazj7ecRNf/iXdqGa4V04NvY8NkXGxEsC4BA868hSNp32yrOJmI0RoyqAuzGHJY6/PtHGn9FH0hZ
JsdqWDUKS1bbsFYOly6rBBNwA3LTCjKmzq3x4m0GlAslGSCkQGEBX97AS2wEV8sS72K0K48u4Yug
agZX4Si96Sd9NYpW4sZlVS2Mlcy9Y3c/Q49W3wqrh3C4fbOOaNoAP2Uecfso3QPphgwns3w+Y7LX
x3MeSgoUA+/amyMwuUQkP1boAoWt4j5RuYwuKqhIjJgV818TL96nxAw7rC38JOM4jTBM/RAeykiE
/yuybNGiB4Si5g8CmvjPnG2eX7IBF6H+fWNitxB+G4FtyVJPfrYReRdR66frFRalzGKlw91QNmoq
2p738x/AqZxWosS9ty6ttT3nbGaSwuuhiiDLJkb8rwH9K+lp8/8LQbSZBnGHKi7bH+n7h2FdH0C9
96tDNvkziZPBfSxTa345Zkj4j0I8bo7F8ZdOv79AUVXINk6m+XVjE/v+XOsJXrKNFjss/D1z9iai
HtX6Ii/QA3yzYiG2fxfJCocUes5pbt0YLmbB1jtAva82jaIAedXO8wdg0wDEcsk7rlPdQpgGBfcV
J268vqYUZZt1FM3BaTIHThFV0iBUPV9xWsvuaOBRd0Vv0lz3Nn58/xECWpgyTUNBygIIjmQEbryV
DKjLun1PRuaICcG8Qo8UBMIn/tNhIN55iilCYcFpx6YSx0EEbTUD9V3O1ZKADgVp4qsdrzMCC/cv
bHUd9wgUjdGKXbslIFzpuafaaGmUeFiaFp7dm0iRo/5arFXaOYn0pzzAEBdW8ROAcAyfsJk/El8a
TKlZiZgD98C4YGYyUdmRyfSZrrPEYvZNzlMCS/gv3rzUpw++HrkLusHRXVo2eTEe8ll3uFT/2vuR
itHqRy1Te/EKrSLxp+MVbwFZ49PcotYMdXLEXlR/vKjXEDHsSFEv6oS1yi0ELvLTba1DXHMosyjH
yO20YUIL4+WkfkEk3DiwWshfw8Je3tEyUb/jXvcyoYIeP1OjQdlR3ET3xmLkRfESF7NzRm/jEYl8
P9tueWdg6MEqXnXcv1JpgkB+Zn1wL9+Nv4mCJV9sl6vDSjE2pnqadMch1oEE6R1NFuT3OnxbfvOW
a5vOT3zkOWNfOv0j+bFbO3PWQ+JYnnp7zQ7LDofCNM2m5M5b1eXT74YXWYIsqy7CiSPR9ZasPYNR
5hKb5vKshEA5ezHtp/AgkSimo/j1mi6NRpqDbSTB5Aja/a3gl5O21zYmvL6z7oKeYZC+hTmkoYcT
AHKk2xr5hWD/OkcfO73mdyN21/8E+pT4WGzchJRPT3R10fwXBMGMN70YPZ49JXIGaRBg7MNHMEoz
4c1jOJGh/OiWw4J8hc5ZNwc+Z9hBMAPzviOHrUBgM20kdz/wE+KGenF9C2wmBCNltluk5A6jo2w+
+yQLhqdzrVcJ7X9wrkOB1VtoVpcro01h4ex1H2MvBwC6sG5Je3h3eDVUI0Qks4jOVipw55WezAn6
RgP+eNFhUaFKHPtGn+sX9Mki9olYvwLQhJJ9ZcbuxseOdR+aOuRu+PxAOQLSiKEAp/x8+iLkZXd6
n1ZliMGXjijZaLDSUzyOm8/yTVEVkfS2iaHpa3t7QLgMkGoORjMzZHgbO2J18bJEXSucxAwuD2Tp
YBSaCAjuE+T+tXc8igvdi1JPqGwOnRrancqyDv076f9eX8EhR6PfK5g02X3ho1bBCVqKM1Ak5wl1
A4Yc6mynDKYfXVbxkSlqAejaugYgDxsH8aZXFg+aGORxoRkyngd7KuuihWMP9vWKnSvUTLuFMkW9
oSJb6/hvtMMT1t8JZJCDheHD/5gU9pGwGzpj433Y1QIDAHIJz6UEJfTotFOZ3GGxtl+pqIDqzOyJ
cK6wWUUus6GH2gw1ne25HOfikLBv9DdJUtz5XiHDhX6+e7d2XK2mBlBuDe1LWrh5EAz67WxPGc2w
UsvlsrkCXGMoE5bwFY6CmhHvaXnXf2hxP7nn/0XG4MiMa5V3WAPtYhmw7CncjBoMS/m6rmkg18sV
sF5tRaUBn0t+rH6wpGySdOhIu35DYUscWlVoGXRDEP8KT+jod0683KOe3cUES02+Dho5Hysd8jv5
NZNuqX9mwzxcS/yXGC06ODhJVcc39fpecLjfR74Jz/ConRWYlR4SzD6yT+qMTHYdl6RWLvKf24Tm
kWU2XkLwBBXDEOVKQOdPi39OiteCy5xEKLiINgM9YJvdomUYXqlnGeUK3oLS9Na+oXPXI1vtNRgl
/YGHhUymzB3fV/W9qrO4S2j4FyxPBwBCmgsyUVPzQY2pklqyTJWOL/EemnnLTiUJ0c1egAPOLyqd
2dSTIL1aV5LDAOsgrTatMvAim17aLu9lelUSB5jASAr3Vn62Bye50QmzO537bvn3bDllklSvV6Sz
uZVHKE6rNojzCNVqtvpfr4LeZ5BL4O2buKYTCXlH7uNLM6V1mQBx9euV9wCN3UsbrtjhsmmnBhcN
NHo4s3ecuTT1HNZMX3ev1zUE32D/dFR6rmh9z+j+jtokJ+lurprVBrEnOxxRFhLRFdnTzdjThexo
MfxPeqIkr5jAlRCsLU4gUBqfc7G4Fv1AQfCsHsO88mgvUlgNdDZBWTgiga2yP8NrQ+HnsTgqtTFu
8/Y7WLeMOwypaSU3viBLzTy5g9HE66D3IHutPskdFaRdfaADQgRVJRxQA6ABM4kiNf7vciB5q0C+
Pg66xz7wpPlMSMnq28dW3SLGJEYc1vHPaAFl8ru3StlzqOqc9x2byTn+fMKNsAJYEDwYzLbUo/eY
6R/QyRaVAkA/71kc4CEzvaEZj3Mulx/O3vCLBmgKkhUBH4lJr6mLCLJHBC2f0Woo1bxqqFwKwq8/
gihwoy/aZXIfEI0if0kvmeNfPOO/50FWGL9NZchNIo334R53evNmplQveVitVCkqF3xfKcCY9xSu
yiS3aXxMQVrKVPBvXJ1T7aOxl4KXpuqzckvl/A2WXK9NjMhUt3iKFEUJQy2ZoJIUGe5+Ix4P/Bhs
F10sg/lQ6kQEsrE9ISz8orMvbhyNIvrVibHe8BO1A0R8pjquOI8wdbxSD+biyeocrRjwxuetjCRx
mR3EJtvB2CvjNw7kYkPOg3dz83zjtYzxinBGePnLYzY++EVsnsUYpZthSXCfRTz2mHeSm+iyzaUl
5Ceea+w2dGcBgAWUn0NZvzoXkoE1paAo4lJ0LN8oBAQ8eNgoilR0TdDm5AnUmDA5MGi3ah8YGI5e
nxB4p+3bDaeOHw9TNOuYSlzO8Y3BzTm54TfJuY4eu8YoCi0Hj9lODLxpmO13qMhXdHBhLNPjMmjz
0thcozGvmCSqHTv6vHyYtyXsiYvTSG8MtVrM88btAn2fDhZ3rPU0WlS/oI1Wu6/z07v5j42NLNbB
Vyw5XSyEMts7WOeJJCt8TgKxVSoQ7LfPXkkHiy0nLgoub0dSFH/WCrN/C2IG1H/IPcZlUqR733P+
JtXlqB57qRZm9qBHhU2FzBuRrtVrKfkoi8aeFwx/TFTxqWdt+PZpCRW4foXGKYftx1XEcdKzDDGe
MDkWhgWuIbyYZvY2vGJd8XwspTHKHdF6n6q5yJ4G8cI44W2vXxBnkl0Y7NrtDv9PVy3H+93eIe1M
6m5U9/aTLNAJoBIxuLEeutlo7EJdmttaCYYFxKlROJYiatdG5uvFALGtBwAGO2v7HmprUxOWMsWZ
17ogX0tW3MyxZmwRJZRAqndp1F/EG41mmpsQj+8phUnzorAAWxzhNNmLGwUN9obPPzqAlPQezMnf
IvheGIN9mPr/4/YTGWBKqrnel8hZ1TG8B9q+8bLtugAWFoIZRLL73cN7Igia88ukhiW+r5D8dvrs
bUKpRln7g1iwll/vuaDskNonWEgld+LWc1+b1s0kA9iGYmP6HnUQ9pEgmss4+m7zpAQIB3zA82NS
srTp1Hm3pWRZbJAdWpb8eZ4m+jvDV3HUq8ob/8S8ySQRzkSJn6kSOmDPBqEE0uibeDwIH8XFiXOQ
fKMg6dvHIP0EJ547LeE5En+1YfDlfRHavNNuHfiG4BS5+oFfnm0zFVWlVqZ5QIl0F9u+WMdiBgGm
uXRrIscUn+N1yczgpyanvasR4d5ji/EYaGp0ZPbOM6oM4QJOxLAMwWzRY07aEam5PR/YQ5Tds1XO
2GRV1NS5oV7WATIHbnz/EEkNz8wDciIyd5iMvlHeyV2eUzTF/mYcVk7pxZX7/Yu4XmZhit84xT1j
/JqpouPx7dSXP/aGlT93gvty8CSJQaQjsAfHzXNga7QYBsJgjOt2bwXpc7dtcn9G78xRa9bdsAN+
qc6EwHDgjmgYKCGqbjbR7/r2nECWWy6s+M3diggOflJ0n9pflu6s/Duq586j/BGAlVdzPH7dp62z
IFsjUbBAHoQ5H4S00c10uwgOnX0rfksxbpcyFFWKkZ7KHMSS3OWBtcpF4jUsTcWRq5Q3JrR/BaKj
EPGc8LRsdPbClizUyTs7Wx4eIxx8YZtb2f/6LvUhl/Yj1/gH8Hj6bQoCnmg6ZJv8tSZ2IjqT8Dve
7Q8QA7e6bE6dxqoZOzDFEYJJZCLRXVnKlGTuhejLezOSuQxwzlM6UjBDhFoSzLaIl/f9mYURSh1H
kpvvxyIlz3ZHFVfiaWqpc3lET0Tm5vl/bCwaIvJTmKZwZSa15Z6+JXsReCELJPxKkwrbZkyLdr8l
83fkrECMO1gwvMDJmM68wWLaOKxfhaYqrxbHmibsBvaHITrVr2K0UEDstmYyvXrq1+5MAdXoAmjn
/EGIta8vcgLKoh7CCjQm2oyM/SvTQ5iPYaUf1U593Jouppbkoxh5ey/bkjUZBlzzE8xfh36LxpPr
SfVxi9OuKoB9ex+i/blHC/qEFqprzDS7s0BU75MgWoEtcwZyfVnbmw+8bg+OoHvdXe5VM8+NiNwG
OtAsgJ4x3lDKbZ2HfA9NfClpJEpE9S1p0UhmtkaVFivZkORg2cT5y/1VC3LU31rPmvkJJayGL8+g
hv0o3xbejlKGuSdeHe8yGNMSnBkgW8gj0pvHHcxW1EasULX737ksnJgGgB4IGnamLzGk4lYMzaiO
ppnBrfP0LxIX2rNgriif5Ms9mb9X6Suv/Z9Ilv6dyjiqfHdXkTvi+i46Q58KKSyfY0YCcx6Uvem1
x7vKqpK35qHkBvIDX+LzDUNiFDok+XVUNi+3h7xRfyTiHnCklUKGAvYepuNnmh1gYhNvNWT9Kf9X
yi9AQgDNsmSkt6F8lcfP0EqfXDtGcYuKEA6CAt8qa4Rer3otYMxofN2G0gzuq+Shl7FWnF/0aMeI
G49uVei8mFjLV3unizPpMpAAtHzNHMFiyZZE1n0+/DYNe0tx+gRKztQdBEzGLOQ8Hi6ajPkbmSpC
lslhPmUlMdRqhd8jDfmhUyduMcSSwg3GqHkd0556J6jyRY+/JlL8g1GJv3A4lg27CPQA9qkEh28n
26s3xKQ7b4ii2+J8Du3f9izVA4StgZuDPBUuOEiv9VinxUJQbwgZlhf4xP/eieV8vHYPPtpi/mnH
BZzKRqn7oNHyg//NoNIvl78VOlTeOQMMSyboh2xPsCgQN2pgfmWnVDtslLRfZjeVQLYqv42R8L/j
R9k8wdxiaWYxnExyNdxvMNs8dmpFrBRNQI3VJFcue+d3zcexRwkuYtll78hRFv1kWpCfaCX7wTM0
YICJlb9as+Z0bVErvVCWUFX4n7Mhx+BKf7jZG5RKUTMmo8xTHK04jOLUxQsXYWdaP3gXMnDGIALu
KTLNQSF4BSqOuZ4fj/0b1muYpw76rCIu+7tv/17wPfyINj6qF+3NC+HmhkgqmrReiQUCKPRUmrlF
AIq0uyKBXdADUiPIH7v/garAOybL3TPBnw0wUdRwfeWng0X660PsD/FPS/S5lzWjYf6voxB/H6Mz
8EWrBBOZKYr2c82VNdw4wHBXgB1U1dOsO32RABYt9OaTgpyTJrMRSP74YnkrYLlxEeK+XaK31IS6
HL0HPArGf9pY+8riYXODdjqiMYqoW4gGk36jdEiOpEgwe/U5/BTaqW+ULf1Cq7AVwzi85kqxzq2c
USuHDDw+XS2pTMS51/ckJRx9hvbGSCFQ7QOXS2iBqqimTF1gfnUopCXTBbrCCFD4zDk+IipuTOO/
onOhOkM3BwxRzGfKAk+g9cYaMQZhaNTsvr9vF6YAub/cBfjrJKtDi5ecN/LNYYq2+N325YvIX1de
b/WN0xGg/cyQtelScsx6R+biIpbwrKXUhBJRFbUBBOU5vbpuf3kmHpB5iwAgvJmZw0FWhUUWWFOf
wWFQCM6YII/PPCe7ECM3bke4orqt7rE5OL/syFKhw6KR1pnX7aUNuJsh3AQuYMAHkSFyh79+y/WF
Z2BndHC6631f+Gjt0FfIQU7ITzZHnUHH5bHsWCuwATcwD4gcGqi/hFeJ5xBrhgptVrZ0tSQ5UvSP
pK1t5iT0NuGYSnyqnOt8hHMSO3ooD1j99fpjt5w3LVPEfF7Dd1kaIOCwpHrlez1VBreMtnBPZZYN
S/3iIww3h3LNxfuHx0Asw8gi+nXeZfLdwBJA9joGkRGchaJ4p7JMJz12dG7um4Y5FZ0i4Q1pQ52H
ulUykdkYuUy9ibwU2829Lgn6Nq2Syg4nKsWGNcHxpceiLX9XZinuHCGp3m/sBDinuS/VrnUpFBuq
wPgxQtBVF5K/9clR5+PsFeMI0MpoA4fH1GI+5ePQ22Bc5BUUOCP1ZaI6GltcnP/UFj1xCUZXb+o1
JYE47a7QIJJQtApuwUUzPZNmc44WGrI9tt0khC1kyZqdPnkq/NebWMLVZvz78HGgQMid75IEOLg1
7gxqtxRkYBpNQExjYX668DzBUBbnzWcpYNQgEj6Cxz1erw/i74iWtXB9KifIfGP0UXQIS2LSahVc
dHRxKpPHgh1d0lkc+uAI1LEIXmZW/DHt659ZOIqodL5dbmpmq791F1iCmvxaUJLXeTYPnR0MOKxS
NeIBmqsP40bVQMeciTbPZqBN54XlZXJrobU68wE4D8aejeg8VSnumR2ydnlLq9KW8wDzY3BTQgdg
prpZVzdWPcE32ciE2l76B7Bznf6YUyj56mdX+b0oUC2qaxMPkxe0B1jny1v3ZLH3MblDLuAlHvor
DfuVYK0oiV2JdAmmzQj4SBRS5nwSaW7sPFUAWpam/UQgvNo21Y4ZOhCiitAKjZE+dNFZ+2vKdJxL
fmfTgLRHXMY5WNeSqi/1C5yGon1I0j6lPLBWs67St1i6UyZJaZ0Rn2kTfcaXrJDdzS60RHowka7A
b8sVLVgqGZ2Vas82wn/fploQJNfZBKbbTqnjY8Ns/+LgcBz4e+MNd0eOpNlWqBfeWWJptsGU/Z36
Yyy1hLfAzedOIhGo3ZwI0TZQPTHMs+cikk33hv6Hnu33uqc5agePeY3v9b/Op/BtxN55zPqUSy00
aKKCVqXzHpqiCZspyQaUe/Vfk4a/VuuAixjnzvOgjC8TzoKbVAS3n79OR0wAM1hRXhVjyXR7uU4C
NRQ/v3UKk2E45RLVAmVLBx3jmVNIvOr+qaaNZLb2wVoWZbwmTJ+LtKxNFK1AWBCm4pNGDSb4rO1a
PZ5AJotOj0080FKVfXTD5/238Qp9gXK4rZWOwEe2TaQOvY0d3xDbK/s37KTWpj2GdkEThg0a0IH/
aFBdqX/gCZ2MfDDGWudwuLmHuEOnZ2Wpq2Bc4KZ/SxSMAXnvQLBVZejBVHE/E6gj+HPQYszQpNcR
0qlweQ+nNiJojZQ7I+IgQ91TbfXDhLcV1rIXm3RUkiqDg2nFYjUUnOi+VYpNl8pEhLq2n7NmsJ2U
emznDla2ProgZB0SAo7q9CQmcPoyovtbMC4pnkuusPo8vT+vcZUN5G4mgp2TBusvfbKOzKS6rx/M
yZ+cVyuf2jYnjDiRqIXhiugB4BMM+j2nznXMviJ1zEV9EHP94MnZT08bF8NYSHMmVym30Wc94K7G
ZtiXajTw+jvfIWRJf05uxAxNcbc2AUMXwN55bu2huZ7z6SkSymk9Sx91UsRwKOx3MuNRTjk++stR
c9JOTjUabn1MX5CRDRLj/Ct/jSdh35FG1tf72cbeUZ0c5oXCVxz63WMfjeFMxGMYe+Fz2UXiIxRa
mQemewyPaS8diOSWK5hYmN9NAGC0kim25agckITcZzWsB1LGqnB1gq7foHtcfbocbVv+INeB/J32
rBklKaz33SGjaQ6CT7iWj7UG5kQIkJ6lreU3HdO+h7qd51N3QluUdPoZaMI9Z5Ns+6WoC8GhbNO8
ts2328sgz+ilz1D3X4D3YjnpwRyA1M2CUP3xBAZzk40r0kSfsjd0Lgn6jIeunVU96aWTBWY8ySiP
SD/VzRGOSXEWrWZVLcMYe4X9Ek6Pp8f+oYwrhIUteySaMmlL1wWhlKx1z4gqkaTBK+3C1MNzEOrc
BKt2W/N2UAQ8Okn2Nzl4DEH6pc6a1uiPTabLIdhLDX9fF6wYKdTFjlv8k81DmR4ifDcBhsZf6Emf
LlVVUc4H69j8W9SocQa4gA+kt2E0lhP2gf80r4tOgtMbBK2L1D10ASnRrjeXyf0dKShDyHuPbxmM
USm8rjhhmBfpbcn9v+4gGJN9DbWc1+Exc3TDQJHdVvooRRKA60axcHfm4OtbPX0kWgJ+o/nDWdcX
3jH3RdS9FCMOt0vxr4nFB+lArXhoWiHFHPxoepU4EOozL5/rlmUyQlpicwQ6cQ+lheNxzFYqCbd7
SV/dWj4AWzUO7RJmsr9hnQg0cYdeLAJ0zZlCOiaEEqNcEkSd4eEUa2m27hhe1Ng9iLqIK8PmQOhb
c/3pJ49OKPcKaGjBN8tzeT4o6eTA3RYNBIsDMPLPJxqjUKO7Msx4HGTVpiEVN+KcJKojqD0BdWXH
xltOfVTULyFfIuVxVAeoXZB6a9Gg7BZ3lPfZ/DekeOWGMkDwZNoMwF9v/Nj6knh7bharD/XljRlP
HsWQ7SJMlzc3ml0Q4/hpqiR0iwm8OEL6+C9LL2HukmfhDbLBoQwXpvI2JLkQFIKpSRIaNz3ojXG3
M1+AB2LsuglzVwmK6pja6OS6Y9mnr4VYn3KxVwHQJwWPdk7h0Un8r1dY80A4lMzeKw9RiWcyHxw3
G8ndlRnLIM9E+UH89/38Aea5mG9AusCzlpBpIhjMnREM+hxQoHicUNxwT/aFbiIiSa0NTzDQkcnA
LfY6iOlyWRILIsvtor/jJI4ORbpHe+EP4QG+4Zy+IRURpWWZ3TekQnFmMw4MlrhXJzfVyP8nmLtL
Zpi37S7NocbUA3Mr6cRRYwXlTjotgJFkmzVoyFPWipmS3C9Z4MTJPDdabbk2sJijMtFEu56/gKq2
3xLmLyGFrdakkt5pQgwklVaAoaK3rPk02kibPySbKaurXb+aooPm4n/CQp52mmDIZiSDXYAlZ60W
ZTjyMrJTudqJT2hTdRzdT2T2+ZV8XT/cnzVNB5o5EMv0pmxas30bw4WLRW6m26j4Tk0RRcuMCRg0
uPyXyQQPgU8JO0AuyZfTWGQoNj0KHsVU3vR3sUusZfOUgS1nhILj7GH4hzKqCkVvfMzBU3MrmjSh
v7Q62snG13fw+XraUny9Lc9T+zDXbQJUpgx648S6vU6uiNoYPt11yiDy9UNv3FrCbc0CGLs2+R0r
pYbBV4IKL/qY4+lgfx9mKFrbVoRUefwchbUV1BvCtd0JJMRoxB2YfAi2efvhQHOzAYCtSDSXM6AF
2w7g+oLn2uLcC1ngD60dSyXIQk5pkeUg6TLWA2EZ6X4L06Kj0WWi+jTHSS71bodELEXaKln+ldWN
JEJ9yX012UpS0l+mWD9n/2swFNkjQl/COsIODF8HdOSiQTPbF6cL4hT1NeRXWMVmUAvdQYmpl7aQ
ezre4Mi+XlzCFTS778amiiR63QiE9V2Pj6zKI/qSaJmHhzacrdImM9ZDb+sqDXDpCyfCaGKEG57f
puDeQBfoORMh66OQLl/O4QF0nYIyFR9PeoFjdWzcNQtOrMMdoltSWtkqr+PBF6HUU/bICCFNpiqh
dHxgi26pq9uRPs7khiflxOiVWbUSZDnwk+Hlf1rcDzBVQNjLUE49r3AqUpCK/hS/fEVJrk4vrVcf
oz0/xpAsFJksVJbiMxg4PuEkODkcftufYiwbxFtcB9dQBdSoUFbkz9IZa/r08PH0hCWlohTWmMFp
xA78SJlkzDWx4pRWi6rzS3hFFs4q/Cbl9HRxuMYmkAu4kY2r/+mvI45r4et7HTwp0cmUf1Y4t1Eh
98w5tGgzVLwqbi02hEh82c+bn8rXAUd2M0ny3oxBXeXHAoWbCMDg93XegM2CbNmSWU1/SDyQ4p5I
e0BpNxqtWuFSEgZ2hDCjFmw9Mw5pgC6/lYHY/eHE+mlM0y4hTdfWZs9PeBxnZ8Ek2vWMQLgp+Bf+
tvRTmhP4M4SuXnFvv9c1/f+okcpZc00IAz6NujC65/iR/3Mz+eRCaS+HMHdHo/FNDKjEYAQiUBgy
qvSdhzaNxGKjkHJlTJWbzt+yNZrCw/e6ejBSGSnCvXl1DcaSQsVflFt5Y3eg8slmjc5ToOd4X1Yi
2+UneF3J/bOaqosny0hqY1Q6kjCg45D8zyMi70XrtF36yn+dBERrpn3U1hX/Ih45FCWEhqgaCQ39
CP7BKDsbj/9yqa255gpFF15wem4MWw0Tn1AkAm9J+hHSHM8tTMU3kgZ1Cgch2Wj66UwR5NBJdsva
9d5ywEX2MDH386dg6KuUEQAxRtW9ArcvVfNI0t3by6jeeYZTYowbi8teLkWQDvE2KuaT0AsN1Eqv
YZk7mdLbosRB+INPdNT6ojdIs7mJ1h7o/S0swU0zrrpPkKiOgJ90EoUoI+35+iIk8o4tB9neiR3E
r4osehHqww0wBSMp8i5MzyjwxZLpCNBQ03vQ1tDjg+cPA0uKMTyV+SWXRmoGfkVyEtuwI6XhARKL
QMaZI8bp8ME5/ZyqhweVPuiNHIRgZGEbcwzkhMfU5+KMe2+Z8ko3/RKfuvdpldlsWm7EorVbBa4/
o8su+lbqABcOyJsxsEg5UiA80cn69zSSLH7urvtrqbu4o5T0C5KuKnmZiaCzIb0BJhJeXx2mLrDA
Y6PVavGyfWI+OD9EwWR/T906cf3iDaCo0t5KePdEq7MuBsE/HfTVUqkTF4a/bIUQgNDygZGDnmz2
dqn5NOQ1+WaOjfgwfAznHhOiTvz8XXHvUojL5Ap/CDnG7FYT/mh+1qxDyuXr/lLjTcbV6zgqmFTx
snttMbEdUBz58ZQ2mvULqLWtXv5s+VGxUJ7iaNpFoxEqMZiLVVnCb0/qAypFPw/ZsKnVsGYlZhHE
NzEn+M/THndNRgpYwrH/aaSTsO5ai9Ph0HamQZMaPbz9x58o8fF7ZcNJJLVWzRxV+/9cdBggRr9B
ZNv92hM8f4ezcMUNRBG6AB/5WILJ9EqADNwR04p0zsH/5GxuaJcC4ZSbp83xD9oAKa+z+xTju8/J
JR5gQ18kFf7dttTCoMgkcigpTKhXiMZYYefDET5CjWCRB44HZ5V+1rF8dLc7+16eMJ0Y8bN6rWBu
YXYOdyORJvx2uvRHuLQru3++w3xqasEL7dRWdWDTc2XS34hx7rl7tm7GzlNmxe9uXtJK86rElLV3
zEkV9LfuFUlP2J3hDyAjr9B8uYy5LMnrF3GS3u6g0g4TY68nZLScNl4wA0Si5IGOOQoEUpDzy3Nb
qubQUyi8aa9fgy/qXcLs4rxVDFWbKmDGCYkyj36QRJ9JuPebJ3NTeno1OhI0MITtXftlJ16aPTsY
+b8tKv6ASE4TuKyGmuR6vu+yeyJ4L25PuOuRzbKhjbv2OsOQrerOpzKHMTIL/EwTHDbMci0/fECv
G2WJna6znW+ACcLEhvc7CaamCrQRxBz/4xRTOK+rrpYSNIuy8YOz9xwfvaEmnJvk/FON/FGTewGc
szhS1AAqF1UID+zwGs2YCMOErKs63JyRmV7IqcPQrrvbB6H4tkv8ax+W4dKXNYbyhq7sStAuD1lw
HwViAJREwI8CSWvJ4qO7NsDLrAEzGdFkXSkvrwmZiit6voD6j8D5m0TPX50SGiAjG2alyhyasz/y
so2s+wGq53wVxPTTfg5+mcc4uHE+GvKMSD1STmEcYzrvXj0LL/htCe37geP35CA1iEaH9qTR53nc
llBOJCBb8LM6HglReS0Cf9b1UHj5ERPTcu7Y0Me9GkrAxPnpdBb7HPpXcMuRFQATLzoD50LHkThb
Ir9rnJcJAcPYjWa6hgFoZ17RQ8n+rVlBXHS7HKmD3rCR/uWDzeR1g/3ur6sgdXQziENwWWlwSaea
DuuSQCC1TMHhzoN1cX2LojYpxZKOWfTQkUXIFHpieIZIgx716OLIcFcmYNFBIOzHiCc0z17zuPnz
9XuO83j61uMBg0bTj0BtOqo0c30tUs+QELdVf9oJV3IFNTdIpBSD3K9qbw25dQTx0z4u9mRQKyLJ
wKA6isUF/r6OWuEPEznG9GLBvuFsVcDYYKmEPo3VIkFsZGZodKP3T79LoLSQviug89JF7xZL0d1R
skQeiq28s8QFLfiEgwFalQKDCNbHTr8MasdaAFHL7f8ZSDwfopYWfpCXRU8X6QSupUv1CECjXYK3
sDAE+dCRQ4q4Z4sAby1pznACGt6MUQI7LwSlWN+P4oNUw0lfUwDIJBNJJTjhNjh5+vS9lvyPo6Ly
5w+qwEV2j5CtLtQuq0dN3TfA7Q6YHzm5aZHGsKV8ZeD5CEaYYWJDxf4Y976dgkgPEn8ywaqMW7ZR
WPiOGxIRMedft9MY/zoLqRXi4wcBFnt4Ic5pL6aCMeMAuSfW4bv+SJ9TO2RedEQ65i95vPunW3rT
/EmbJ8yrC7oBtZg8k1SiVKGSOxsamHvqG3TSVtMkmiyzuRbyktDvoTYZlI8L39WIQ4RD6kLGmqpe
YPrn4GlXrLPoZZzxv0rhTbafTC8b91ZCI8ZpEX4ELYRhMueUasVa2hkYZ9K6Lo+E9gFP2XcCCSUe
2uVBCxtAiKTuVRO2JHg1kVz1e87OCKx2V1gVHbRvT48zGYW1G13WhELsG0ed9yihDDjAPhWESzL2
5P63KaYXWGn1uERXB6ipA+KpvMYMTym6sVPTvU9Ec3lWm+RpUb6E/WGxBpwhdzcR7umWWlv1ltyG
pm8BBF3b2aEj0Ygn99kHct7yztaY82tmdiQU3XL+oCbeEHZrbV1ScywN57k2246aNtkEyB3IbVWR
Giai9T+bkG4IQhgDU3Z55WshU2oe2UMpmbfXz7KrdfeJgTLjDCsR1+TAdvkAqMCcz1Wp3vu79vfM
xgX/qtho8LhSdXYyaORrKRydmQKVOjULEvImwVy4KpuS3S/3nNmuyRWQ3GkwV0dQLXPxXGr3Utpy
Uju1G0qE+pu7Bdn4tI8uGdw5XPZsk/4dN17tauW4oRZorrTY1/yqJx+Ucko5V3fOaPfGdcO1gzCB
fCaqA6gEv/Ce7uvFA+kAkfJf9qcUGkZ7iQJ43grogEMYMLpdJwhKZrxDfur4J+feMtkgJFQZQlIU
fJ0YMi1de6X7KFyRjW0BSu+wUbLY7HiypWWqSfvve2sB/qk3vNbuEuTcSLAVgslcLNncyLuE5ENH
RF/gLSSk6qiWDAY4w/LiZF7rsH8dyUUEAYVkRPB9m0w6aUKyQ44u2PIDM1/th4UueT8EaUHcSPlM
kIPw+Eu+iGrH/bMnIzLTmiFxvh+57t/oDGZFf261fYmf8+S+AvD0IKy6VPESNyuscp6pCdjF2Upo
ORrLuWiDsDG1F6hgKfBaTYb/DI1qHCxx55hG/RfQAw28kw8kNKrvVtbtEsOlJUEq1036biyg0rB3
0XepTKim5S88i8bjxPoeij62L10OZoX0xEgpEI1GraqCsO/CNRVX0/ftsBEDabYP3wu3xeg1rMgC
3UXHXwe6/U3tEQEfmnH/qtoHHI+V0a0EPiNqE96QY9A+9Wc75GJjQgAB7BSC0D+i3L8eN5frBXYP
t/OAK0P4ecgrQbS3T+YMW4EDSHvIkrVDHlUxSLlrd0cPaQNGgsXQbGKD2JHO7mSD3V+6lOYfQAZ9
cL/gwSnCWXeL1DpSeMLzz0X0UppZUSDOVhxWsdBIvl3PKJU2Aj24IHr4vs+nfdRufFThP/3cpqkH
ZMw8Jug9i9Wnvn5/QlxFkiW1r/iEDAbK1mVJ+jMW2yIwu5sVHMr/WTGiufSC7cBq69xYC9432rDB
H2GyTRsJbCD9dksWiCXcrmaOGU/zVtcICEIr5s+ITIQemIcMT4CbmflUvXGUTX9lEEW8Wh1oZNJ/
Gw/ucKUCUK8fgLGkWheAhmR6WToHsflVQsRB1NLrjduIOsgcLUHQm4SCWDnDlQsassN0KPXtrfpV
azDLgspd+J+LtrGyv8pvlEYrEW411JCGm3DSfN/4KtZDqRJ2WCXLj1xZhVEEIUlvnbMsyXH7cwDZ
JvA5feSkmiIOX5zS7TsJtd56SrETECEgKlVRsm6/KsOOoEPR8aehhgvY7lBOsgzQJXrhuw7Z4iqF
k2XKSWsNqLu+MBGOWEa1C+al9GJoz5fp1sPwfJIBJ0DNpuEnHXc4CvnnbEyb22qjTO2gtihWVlyB
+7ZSbIpu542QZ52pXlON1QxRlgaz1VJHydxO9FFRczosWKbz/QzdBu8QgOcbCmG8AQJqn5YSIHG2
6jkm94QqHIqaYjgAXCxPsRSCNIZJglj3SCcjhujooyOgLQeswoMsb5PeJkWP4XmqV+NDPAjcPAgz
n9T/mGPfbyXmHHgwCOpeEMGLrCDqf/ALSGPXHi5AkbGnI4aJa2AIXL6JkhxQrmFy76R9Z0fcAtvm
26ihw8SCVrCBn8GT61PlWJsFZ5mWOFAvZLOtXn9Dm7X+RE+yvU7/lVSHpUrRrTq0OaF9zWKASmuH
BeyJUZXBVRJkCo2q5/O1rSi/RpOnEcqVkHxekyFN/xIh6Sx+wmEo2Gn6vBJn5+Fx783oKPJvcppW
iqRBNaVXnCfj7HsAiniv+CiEns9JxRcaRKjmf6ZmCl33f5T3oSJdy30k1PMx4KeN96KbctTEDNd1
XDcOp5D1BLyIskVlSZV1Ltn9wgd6AtPE8+UswjTx5BYty0vDb3HKwcqAtEsf5HI6ZWTt2LLiz+bQ
6p+7xflRdI0eN72gk5DL/nfbNI1lBPc9DUi3RSU71KrzitbT7GNy1QZtraBdNVznBwPEKPtrhRQi
FjQgsR5apvQWrVzNrSY4RNdEnOMqdH5VqVysNiekxE21rztppap7QDF+rNs/J6e//YkWcPJmZOjR
ePJDqeIYCZgkCfliVeaXDNIsgQBtvS6SoUld41hAnQrZn8dR2ms4cnDnHl3qdInpn/LjROf9bKLu
Ns2b1HZLPbkdft468CSmPXKKHNWsCSvJEnW36pjiIL+q1/jncBs2I4P4uNxmuCCOnAQG8nWevPhI
TyRYa13D0aEzMsBmKUu5or5P6J2gXLPkQhMOwyFHytGUvhmTijarldM/Zxrl2ACieau91U/xZ3lP
aHSwtnhJUrNnyeFsoWlmBfzFboNFfNhg87FHfC8s/Z23hT7fI5b1M460VyflBZkFDFZnyU32T0yr
3U38GX+hW1eWKMe9kJPdJUBFnNwf7jkxDMdX5zpHoV5BMtmnDxd8xp9c/Ti9eNmPPWunzWF8h6ii
eb3fjJKfqtmC4hEAB1vLBXVN6hIT6nH3UiJi3OaQFuPmEcM15brKPKGZqFlLZ/on3ftUFGYo8xR6
LmXqZaW3gyW0Ir8jJZmrKPgWFZUDWqr7yjBmXSfTjI2jG/0NalYQqEkZU4gJSTqVMKgFG84=
`protect end_protected

